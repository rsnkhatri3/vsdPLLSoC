VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_io__com_bus_slice_1um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_1um ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 1.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 1.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 1.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 1.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 66.900 1.000 197.965 ;
        RECT 0.000 61.050 1.000 61.650 ;
        RECT 0.000 55.100 1.000 55.800 ;
        RECT 0.000 49.710 1.000 50.690 ;
  END
END sky130_ef_io__com_bus_slice_1um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_5um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_5um ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 5.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 51.090 5.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 5.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 46.330 5.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 5.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 5.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 5.000 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 45.700 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 54.370 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 45.700 5.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 34.800 5.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 34.700 5.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 5.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 5.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 13.000 5.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 12.900 5.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 5.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 5.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 29.950 5.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 29.850 5.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 5.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 5.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 62.150 5.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 62.050 5.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 5.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 5.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 0.100 5.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 0.000 5.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 5.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 5.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 68.000 5.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 17.850 5.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 17.750 5.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 5.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 5.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 6.950 5.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 6.850 5.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 5.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 5.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 5.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 23.900 5.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 23.800 5.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 173.750 5.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 5.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 5.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 39.650 5.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 39.550 5.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 5.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 5.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.000 56.300 5.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.000 56.200 5.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 66.900 5.000 197.965 ;
        RECT 0.000 61.050 5.000 61.650 ;
        RECT 0.000 55.100 5.000 55.800 ;
        RECT 0.000 49.710 5.000 50.690 ;
  END
END sky130_ef_io__com_bus_slice_5um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_10um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_10um ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 10.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 51.090 10.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 10.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 46.330 10.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 10.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 10.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 10.000 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 45.700 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 54.370 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 45.700 10.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 34.800 10.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 34.700 10.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 10.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 10.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 13.000 10.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 12.900 10.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 10.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 10.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 29.950 10.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 29.850 10.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 10.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 10.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 62.150 10.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 62.050 10.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 10.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 10.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 0.100 10.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 0.000 10.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 10.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 10.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 68.000 10.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 17.850 10.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 17.750 10.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 10.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 10.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 6.950 10.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 6.850 10.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 10.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 10.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 10.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 23.900 10.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 23.800 10.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 173.750 10.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 10.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 10.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 39.650 10.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 39.550 10.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 10.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 10.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.000 56.300 10.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.000 56.200 10.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 66.900 10.000 197.965 ;
        RECT 0.000 61.050 10.000 61.650 ;
        RECT 0.000 55.100 10.000 55.800 ;
        RECT 0.000 49.710 10.000 50.690 ;
      LAYER met5 ;
        RECT 2.600 68.000 7.400 92.950 ;
  END
END sky130_ef_io__com_bus_slice_10um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_20um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_20um ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 20.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 51.090 20.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 20.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 46.330 20.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 20.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 20.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 20.000 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 45.700 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 54.370 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 45.700 20.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 34.800 20.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 34.700 20.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 20.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 20.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 13.000 20.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 12.900 20.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 20.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 20.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 29.950 20.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 29.850 20.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 20.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 20.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 62.150 20.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 62.050 20.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 20.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 20.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 0.100 20.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 0.000 20.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 20.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 20.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 68.000 20.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 17.850 20.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 17.750 20.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 20.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 20.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 6.950 20.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 6.850 20.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 20.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 20.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 20.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 23.900 20.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 23.800 20.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 173.750 20.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 20.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 20.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 39.650 20.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 39.550 20.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 20.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 20.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.000 56.300 20.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.000 56.200 20.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 66.900 20.000 197.965 ;
        RECT 0.000 61.050 20.000 61.650 ;
        RECT 0.000 55.100 20.000 55.800 ;
        RECT 0.000 49.710 20.000 50.690 ;
      LAYER met5 ;
        RECT 2.600 68.000 17.400 92.950 ;
  END
END sky130_ef_io__com_bus_slice_20um

#--------EOF---------

MACRO sky130_ef_io__corner_pad
  CLASS ENDCAP TOPRIGHT ;
  FOREIGN sky130_ef_io__corner_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 204.000 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 57.125 22.910 60.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.125 0.000 56.105 26.910 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 52.365 20.935 55.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.365 0.000 51.345 20.875 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 51.735 23.155 60.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.630 56.020 0.640 56.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 40.835 1.335 44.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.735 19.575 52.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 40.735 1.335 44.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 55.645 21.550 56.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 60.405 23.175 60.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 36.840 0.000 40.085 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 47.735 0.000 56.735 27.155 ;
    END
    PORT
      LAYER met5 ;
        RECT 51.285 0.630 51.295 0.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.405 0.000 56.735 27.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.645 0.000 52.825 21.555 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.735 0.000 40.185 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.735 0.000 48.065 23.575 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 19.035 1.470 22.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 18.935 1.470 22.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 15.035 0.000 18.285 1.255 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.935 0.000 18.385 1.255 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 35.985 1.385 39.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 35.885 1.385 39.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 31.985 0.000 35.235 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.885 0.000 35.335 1.270 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.185 1.480 72.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.085 1.480 72.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 64.185 0.000 68.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.085 0.000 68.535 1.270 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.135 2.350 11.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.035 2.350 11.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.135 0.000 7.385 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.035 0.000 7.485 1.270 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 74.035 2.645 98.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.885 1.525 28.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.785 1.525 28.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 74.035 2.645 99.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.885 0.000 24.335 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 70.035 0.000 94.985 1.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.035 0.000 95.000 1.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.785 0.000 24.435 1.270 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 12.985 3.785 17.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.885 3.785 17.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 8.985 0.000 13.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.885 0.000 13.535 1.270 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.935 1.600 34.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.835 1.600 34.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 179.785 1.435 204.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 194.865 0.640 194.875 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.935 0.000 30.385 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.835 0.000 30.485 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.785 0.000 200.000 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 190.865 0.630 190.875 0.640 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.685 1.475 50.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.585 1.475 50.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 41.685 0.000 46.135 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.585 0.000 46.235 1.270 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.335 1.625 66.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.235 1.625 66.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 58.335 0.000 62.585 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.235 0.000 62.685 1.270 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 1.835 179.385 200.000 204.000 ;
        RECT 0.000 99.400 200.000 179.385 ;
        RECT 3.045 73.635 200.000 99.400 ;
        RECT 0.000 72.935 200.000 73.635 ;
        RECT 1.880 67.685 200.000 72.935 ;
        RECT 0.000 67.085 200.000 67.685 ;
        RECT 2.025 61.835 200.000 67.085 ;
        RECT 0.000 61.135 200.000 61.835 ;
        RECT 23.575 60.005 200.000 61.135 ;
        RECT 23.310 56.725 200.000 60.005 ;
        RECT 21.950 55.245 200.000 56.725 ;
        RECT 21.335 51.965 200.000 55.245 ;
        RECT 19.975 51.335 200.000 51.965 ;
        RECT 0.000 50.635 200.000 51.335 ;
        RECT 1.875 45.185 200.000 50.635 ;
        RECT 0.000 44.585 200.000 45.185 ;
        RECT 1.735 40.335 200.000 44.585 ;
        RECT 0.000 39.735 200.000 40.335 ;
        RECT 1.785 35.485 200.000 39.735 ;
        RECT 0.000 34.885 200.000 35.485 ;
        RECT 2.000 29.435 200.000 34.885 ;
        RECT 0.000 28.835 200.000 29.435 ;
        RECT 1.925 27.575 200.000 28.835 ;
        RECT 1.925 27.310 56.005 27.575 ;
        RECT 1.925 23.975 52.725 27.310 ;
        RECT 1.925 23.385 47.335 23.975 ;
        RECT 0.000 22.785 47.335 23.385 ;
        RECT 1.870 18.535 47.335 22.785 ;
        RECT 48.465 21.955 52.725 23.975 ;
        RECT 48.465 21.275 51.245 21.955 ;
        RECT 0.000 17.935 47.335 18.535 ;
        RECT 4.185 12.485 47.335 17.935 ;
        RECT 0.000 11.885 47.335 12.485 ;
        RECT 2.750 5.635 47.335 11.885 ;
        RECT 0.000 1.670 47.335 5.635 ;
        RECT 0.000 1.255 1.635 1.670 ;
        RECT 7.885 1.255 8.485 1.670 ;
        RECT 13.935 1.655 19.385 1.670 ;
        RECT 13.935 1.255 14.535 1.655 ;
        RECT 18.785 1.255 19.385 1.655 ;
        RECT 24.835 1.255 25.435 1.670 ;
        RECT 30.885 1.255 31.485 1.670 ;
        RECT 35.735 1.255 36.335 1.670 ;
        RECT 40.585 1.255 41.185 1.670 ;
        RECT 46.635 1.255 47.335 1.670 ;
        RECT 57.135 2.255 200.000 27.575 ;
        RECT 57.135 1.670 69.635 2.255 ;
        RECT 57.135 1.255 57.835 1.670 ;
        RECT 63.085 1.255 63.685 1.670 ;
        RECT 68.935 1.255 69.635 1.670 ;
        RECT 95.400 1.670 200.000 2.255 ;
        RECT 95.400 1.255 175.385 1.670 ;
      LAYER met5 ;
        RECT 0.000 100.585 200.000 204.000 ;
        RECT 4.245 72.435 200.000 100.585 ;
        RECT 3.080 68.185 200.000 72.435 ;
        RECT 3.225 62.335 200.000 68.185 ;
        RECT 24.755 50.135 200.000 62.335 ;
        RECT 3.075 44.085 200.000 50.135 ;
        RECT 2.935 40.835 200.000 44.085 ;
        RECT 2.985 35.985 200.000 40.835 ;
        RECT 3.200 28.755 200.000 35.985 ;
        RECT 3.200 28.335 46.135 28.755 ;
        RECT 3.125 22.285 46.135 28.335 ;
        RECT 3.070 19.035 46.135 22.285 ;
        RECT 5.385 11.385 46.135 19.035 ;
        RECT 3.950 4.535 46.135 11.385 ;
        RECT 0.000 2.870 46.135 4.535 ;
        RECT 58.335 3.455 200.000 28.755 ;
        RECT 58.335 2.870 68.435 3.455 ;
        RECT 0.000 0.000 0.535 2.870 ;
        RECT 15.035 2.855 18.285 2.870 ;
        RECT 96.585 0.000 200.000 3.455 ;
  END
END sky130_ef_io__corner_pad

#--------EOF---------

MACRO sky130_ef_io__gpiov2_pad
  CLASS PAD INOUT ;
  FOREIGN sky130_ef_io__gpiov2_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 36.440 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 51.090 80.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 52.145 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.465 46.330 80.000 49.310 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430 -2.035 62.690 -0.730 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865 -2.035 46.195 34.770 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.750 -2.035 31.010 0.230 ;
    END
  END ANALOG_SEL
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490 -2.035 28.750 2.035 ;
    END
  END DM[2]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.835 -2.035 67.095 -0.840 ;
    END
  END DM[1]
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.855 -2.035 50.115 -1.490 ;
    END
  END DM[0]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.460 -2.035 35.720 -0.485 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390 -2.035 38.650 1.055 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.755 -2.035 13.015 3.315 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580 -2.035 78.910 182.740 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.310 -2.035 16.570 0.285 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815 -2.035 32.075 1.305 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600 -2.035 26.860 0.670 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420 -2.035 5.650 2.440 ;
    END
  END IB_MODE_SEL
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240 -2.035 79.570 187.525 ;
    END
  END IN
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400 -2.035 1.020 176.450 ;
    END
  END IN_H
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245 -2.035 45.505 3.055 ;
    END
  END INP_DIS
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375 -2.035 3.605 2.440 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355 -2.035 22.615 4.390 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 102.525 73.800 164.975 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280 -2.035 76.920 0.020 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275 -2.035 68.925 0.235 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.820 -2.035 63.890 7.670 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.610 -2.035 77.870 -0.850 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.705 -2.035 78.905 -0.820 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715 -2.035 79.915 175.835 ;
    END
  END TIE_LO_ESD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 6.950 80.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 6.850 80.000 11.500 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 0.100 80.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 0.000 80.000 5.450 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.970 13.000 80.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 12.900 80.000 16.350 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 68.000 80.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 17.850 80.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 17.750 80.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 68.000 80.000 92.965 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 62.150 80.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 62.050 80.000 66.500 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 2.610 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 2.610 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 45.700 80.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 34.805 80.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 49.610 80.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 54.370 80.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 45.700 80.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 34.700 80.000 38.150 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 39.650 80.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 39.550 80.000 44.200 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 0.810 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 173.750 80.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 23.900 80.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 23.800 80.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 173.750 80.000 197.965 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 56.300 80.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 56.200 80.000 60.650 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 29.950 80.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 29.850 80.000 33.300 ;
    END
  END VSWITCH
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130 -2.035 6.390 -0.485 ;
    END
  END VTRIP_SEL
  OBS
      LAYER li1 ;
        RECT 0.000 0.000 80.000 197.670 ;
      LAYER met1 ;
        RECT 0.000 0.000 80.000 197.965 ;
      LAYER met2 ;
        RECT 0.210 176.115 79.915 197.965 ;
        RECT 0.210 4.670 79.435 176.115 ;
        RECT 0.210 3.595 22.075 4.670 ;
        RECT 0.210 2.720 12.475 3.595 ;
        RECT 0.210 0.000 3.095 2.720 ;
        RECT 3.885 0.000 5.140 2.720 ;
        RECT 5.930 0.000 12.475 2.720 ;
        RECT 13.295 0.565 22.075 3.595 ;
        RECT 13.295 0.000 16.030 0.565 ;
        RECT 16.850 0.000 22.075 0.565 ;
        RECT 22.895 3.335 79.435 4.670 ;
        RECT 22.895 2.315 44.965 3.335 ;
        RECT 22.895 0.950 28.210 2.315 ;
        RECT 22.895 0.000 26.320 0.950 ;
        RECT 27.140 0.000 28.210 0.950 ;
        RECT 29.030 1.585 44.965 2.315 ;
        RECT 29.030 0.510 31.535 1.585 ;
        RECT 29.030 0.000 30.470 0.510 ;
        RECT 31.290 0.000 31.535 0.510 ;
        RECT 32.355 1.335 44.965 1.585 ;
        RECT 32.355 0.000 38.110 1.335 ;
        RECT 38.930 0.000 44.965 1.335 ;
        RECT 45.785 0.515 79.435 3.335 ;
        RECT 45.785 0.000 67.995 0.515 ;
        RECT 69.205 0.300 79.435 0.515 ;
        RECT 69.205 0.000 76.000 0.300 ;
        RECT 77.200 0.000 79.435 0.300 ;
      LAYER met3 ;
        RECT 0.400 187.925 79.570 197.965 ;
        RECT 0.400 183.140 78.840 187.925 ;
        RECT 0.400 176.850 78.180 183.140 ;
        RECT 1.420 35.170 78.180 176.850 ;
        RECT 1.420 0.000 45.465 35.170 ;
        RECT 46.595 8.070 78.180 35.170 ;
        RECT 46.595 0.000 62.420 8.070 ;
        RECT 64.290 0.000 78.180 8.070 ;
      LAYER met4 ;
        RECT 1.670 173.350 78.330 197.965 ;
        RECT 0.965 93.365 78.970 173.350 ;
        RECT 1.670 67.600 78.330 93.365 ;
        RECT 0.965 66.900 78.970 67.600 ;
        RECT 1.670 61.650 78.330 66.900 ;
        RECT 0.965 61.050 78.970 61.650 ;
        RECT 1.670 55.800 78.330 61.050 ;
        RECT 0.965 55.100 78.970 55.800 ;
        RECT 3.010 54.470 46.690 55.100 ;
        RECT 36.840 50.690 38.360 54.470 ;
        RECT 1.670 49.710 78.330 50.690 ;
        RECT 52.545 46.430 54.065 49.710 ;
        RECT 3.010 45.300 46.690 45.930 ;
        RECT 0.965 44.600 78.970 45.300 ;
        RECT 1.670 39.150 78.330 44.600 ;
        RECT 0.965 38.550 78.970 39.150 ;
        RECT 1.670 34.300 78.330 38.550 ;
        RECT 0.965 33.700 78.970 34.300 ;
        RECT 1.670 29.450 78.330 33.700 ;
        RECT 0.965 28.850 78.970 29.450 ;
        RECT 1.670 23.400 78.330 28.850 ;
        RECT 0.965 22.800 78.970 23.400 ;
        RECT 1.670 17.350 78.330 22.800 ;
        RECT 0.965 16.750 78.970 17.350 ;
        RECT 1.365 12.500 78.570 16.750 ;
        RECT 0.965 11.900 78.970 12.500 ;
        RECT 1.670 6.450 78.330 11.900 ;
        RECT 0.965 5.850 78.970 6.450 ;
        RECT 1.670 0.000 78.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.575 80.000 197.965 ;
        RECT 0.000 100.925 9.600 166.575 ;
        RECT 75.400 100.925 80.000 166.575 ;
        RECT 0.000 94.550 80.000 100.925 ;
        RECT 2.870 16.250 77.130 94.550 ;
        RECT 2.565 13.000 77.370 16.250 ;
        RECT 2.870 0.100 77.130 13.000 ;
  END
END sky130_ef_io__gpiov2_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 9.695 74.290 197.965 ;
        RECT 0.240 7.265 37.490 9.695 ;
        RECT 24.795 1.090 37.490 7.265 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 7.265 74.290 9.695 ;
        RECT 49.290 0.690 49.990 7.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 7.265 25.600 20.585 ;
        RECT 24.900 0.000 25.600 7.265 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 7.265 74.700 23.265 ;
        RECT 49.655 0.000 50.355 7.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vdda_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vdda_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 12.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 12.925 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 13.325 74.655 197.965 ;
        RECT 24.795 9.695 49.990 13.325 ;
        RECT 24.795 1.090 37.490 9.695 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 0.690 49.990 9.695 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vdda_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vdda_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vdda_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 12.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 12.925 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 13.325 25.600 20.585 ;
        RECT 24.900 0.000 25.600 13.325 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 13.325 74.700 23.265 ;
        RECT 49.655 0.000 50.355 13.325 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vdda_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vddio_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vddio_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 17.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 17.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 18.165 74.290 197.965 ;
        RECT 24.795 9.695 49.990 18.165 ;
        RECT 24.795 1.090 37.490 9.695 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 0.690 49.990 9.695 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vddio_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vddio_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vddio_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 17.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 17.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 18.165 25.600 20.585 ;
        RECT 24.900 0.000 25.600 18.165 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 18.165 74.700 23.265 ;
        RECT 49.655 0.000 50.355 18.165 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vddio_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssa_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssa_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 34.725 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
  END VSSIO
  OBS
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 35.125 74.290 193.065 ;
        RECT 0.240 30.880 49.990 35.125 ;
        RECT 24.795 10.790 49.990 30.880 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 54.470 73.330 55.100 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 1.670 45.300 73.330 45.930 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssa_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssa_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssa_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.090 75.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 46.330 75.000 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 34.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 34.725 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.490 35.125 74.700 189.480 ;
        RECT 24.900 23.265 50.355 35.125 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 1.545 25.600 20.585 ;
        RECT 37.280 1.545 37.980 20.585 ;
        RECT 49.655 1.545 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssa_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 39.965 74.290 193.065 ;
        RECT 0.240 30.880 49.990 39.965 ;
        RECT 24.795 10.790 49.990 30.880 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 39.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.500 39.965 74.700 189.480 ;
        RECT 24.900 23.265 50.355 39.965 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 17.755 25.600 20.585 ;
        RECT 37.280 17.755 37.980 20.585 ;
        RECT 49.655 17.755 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssio_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssio_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 6.100 101.975 68.800 164.590 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.250 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 23.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 23.815 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
      LAYER met3 ;
        RECT 0.240 24.215 74.290 197.965 ;
        RECT 24.795 10.790 49.990 24.215 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 166.190 75.000 197.965 ;
        RECT 0.000 100.375 4.500 166.190 ;
        RECT 70.400 100.375 75.000 166.190 ;
        RECT 0.000 94.550 75.000 100.375 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssio_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssio_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssio_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.105 65.955 167.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 23.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 23.815 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 1.730 54.435 3.905 ;
        RECT 20.775 0.570 54.435 1.730 ;
        RECT 20.775 0.000 34.160 0.570 ;
        RECT 44.720 0.000 54.435 0.570 ;
      LAYER met3 ;
        RECT 0.490 24.215 74.700 197.965 ;
        RECT 24.900 23.265 50.355 24.215 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 1.695 25.600 20.585 ;
        RECT 37.280 1.695 37.980 20.585 ;
        RECT 49.655 1.695 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 169.135 75.000 197.965 ;
        RECT 0.000 98.505 7.715 169.135 ;
        RECT 67.555 98.505 75.000 169.135 ;
        RECT 0.000 94.550 75.000 98.505 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssio_lvc_pad

#--------EOF---------


END LIBRARY
