VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO simple_por
  CLASS BLOCK ;
  FOREIGN simple_por ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.800 BY 45.820 ;
  PIN porb_h
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.840 41.820 4.120 45.820 ;
    END
  END porb_h
  PIN vdd3v3
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.000 0.280 4.000 ;
    END
  END vdd3v3
  PIN vss
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.800 19.310 21.800 19.910 ;
    END
  END vss
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2.780 17.260 15.740 18.860 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2.780 19.295 15.740 20.895 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 2.780 16.195 15.740 28.575 ;
      LAYER met1 ;
        RECT 2.780 16.025 15.740 28.745 ;
      LAYER met2 ;
        RECT 4.400 41.540 14.320 41.820 ;
        RECT 3.850 16.025 14.320 41.540 ;
      LAYER met3 ;
        RECT 4.140 16.115 14.380 28.655 ;
      LAYER met4 ;
        RECT 4.140 16.025 14.380 28.745 ;
      LAYER met5 ;
        RECT 2.780 22.495 15.740 27.000 ;
  END
END simple_por
END LIBRARY
