`default_nettype none
`timescale 1 ns / 1 ps

(*blackbox*)
module simple_por (vdd3v3,
                   vss,
                   porb_h
                 //output porb_l,
                 //output por_l
);

input vdd3v3;
input vss;
output porb_h;

supply1 VPWR;
supply0 VGND;








endmodule

