magic
tech sky130A
magscale 1 2
timestamp 1606744421
<< dnwell >>
rect 1900 4721 13988 39520
<< nwell >>
rect 1820 39246 14068 39600
rect 1820 16697 2174 39246
rect 13714 20086 14068 39246
rect 4247 19918 14068 20086
rect 4247 16697 4415 19918
rect 1820 16529 4415 16697
rect 1820 4995 2174 16529
rect 13714 4995 14068 19918
rect 1820 4641 14068 4995
rect 203 137 1489 3509
rect 13456 149 14742 3521
<< pwell >>
rect 2274 38993 13617 39153
rect 2274 29063 2444 38993
rect 2274 28893 4298 29063
rect 4128 23588 4298 28893
rect 13515 23588 13617 38993
rect 4128 23554 13617 23588
rect 4128 21889 4298 23554
rect 13515 21889 13617 23554
rect 4128 21855 13617 21889
rect 4128 20207 4298 21855
rect 13515 20207 13617 21855
rect 4128 20173 13617 20207
rect 4554 19798 13628 19832
rect 4554 18169 4656 19798
rect 13458 18169 13628 19798
rect 4554 18135 13628 18169
rect 4554 16470 4656 18135
rect 13458 16470 13628 18135
rect 4554 16436 13628 16470
rect 4554 16417 4656 16436
rect 2274 16315 4656 16417
rect 2274 5183 2444 16315
rect 13458 5183 13628 16436
rect 2274 5081 13628 5183
rect 1669 282 3413 3670
<< pdiff >>
rect 7315 282 7329 3670
<< psubdiff >>
rect 2274 39119 2482 39153
rect 2516 39119 2550 39153
rect 2584 39119 2618 39153
rect 2652 39119 2686 39153
rect 2720 39119 2754 39153
rect 2788 39119 2822 39153
rect 2856 39119 2890 39153
rect 2924 39119 2958 39153
rect 2992 39119 3026 39153
rect 3060 39119 3094 39153
rect 3128 39119 3162 39153
rect 3196 39119 3230 39153
rect 3264 39119 3298 39153
rect 3332 39119 3366 39153
rect 3400 39119 3434 39153
rect 3468 39119 3502 39153
rect 3536 39119 3570 39153
rect 3604 39119 3638 39153
rect 3672 39119 3706 39153
rect 3740 39119 3774 39153
rect 3808 39119 3842 39153
rect 3876 39119 3910 39153
rect 3944 39119 3978 39153
rect 4012 39119 4046 39153
rect 4080 39119 4114 39153
rect 4148 39119 4182 39153
rect 4216 39119 4250 39153
rect 4284 39119 4318 39153
rect 4352 39119 4386 39153
rect 4420 39119 4454 39153
rect 4488 39119 4522 39153
rect 4556 39119 4590 39153
rect 4624 39119 4658 39153
rect 4692 39119 4726 39153
rect 4760 39119 4794 39153
rect 4828 39119 4862 39153
rect 4896 39119 4930 39153
rect 4964 39119 4998 39153
rect 5032 39119 5066 39153
rect 5100 39119 5134 39153
rect 5168 39119 5202 39153
rect 5236 39119 5270 39153
rect 5304 39119 5338 39153
rect 5372 39119 5406 39153
rect 5440 39119 5474 39153
rect 5508 39119 5542 39153
rect 5576 39119 5610 39153
rect 5644 39119 5678 39153
rect 5712 39119 5746 39153
rect 5780 39119 5814 39153
rect 5848 39119 5882 39153
rect 5916 39119 5950 39153
rect 5984 39119 6018 39153
rect 6052 39119 6086 39153
rect 6120 39119 6154 39153
rect 6188 39119 6222 39153
rect 6256 39119 6290 39153
rect 6324 39119 6358 39153
rect 6392 39119 6426 39153
rect 6460 39119 6494 39153
rect 6528 39119 6562 39153
rect 6596 39119 6630 39153
rect 6664 39119 6698 39153
rect 6732 39119 6766 39153
rect 6800 39119 6834 39153
rect 6868 39119 6902 39153
rect 6936 39119 6970 39153
rect 7004 39119 7038 39153
rect 7072 39119 7106 39153
rect 7140 39119 7174 39153
rect 7208 39119 7242 39153
rect 7276 39119 7310 39153
rect 7344 39119 7378 39153
rect 7412 39119 7446 39153
rect 7480 39119 7514 39153
rect 7548 39119 7582 39153
rect 7616 39119 7650 39153
rect 7684 39119 7718 39153
rect 7752 39119 7786 39153
rect 7820 39119 7854 39153
rect 7888 39119 7922 39153
rect 7956 39119 7990 39153
rect 8024 39119 8058 39153
rect 8092 39119 8126 39153
rect 8160 39119 8194 39153
rect 8228 39119 8262 39153
rect 8296 39119 8330 39153
rect 8364 39119 8398 39153
rect 8432 39119 8466 39153
rect 8500 39119 8534 39153
rect 8568 39119 8602 39153
rect 8636 39119 8670 39153
rect 8704 39119 8738 39153
rect 8772 39119 8806 39153
rect 8840 39119 8874 39153
rect 8908 39119 8943 39153
rect 8977 39119 9012 39153
rect 9046 39119 9081 39153
rect 9115 39119 9150 39153
rect 9184 39119 9219 39153
rect 9253 39119 9288 39153
rect 9322 39119 9357 39153
rect 9391 39119 9426 39153
rect 9460 39119 9495 39153
rect 9529 39119 9564 39153
rect 9598 39119 9633 39153
rect 9667 39119 9702 39153
rect 9736 39119 9771 39153
rect 9805 39119 9840 39153
rect 9874 39119 9909 39153
rect 9943 39119 9978 39153
rect 10012 39119 10047 39153
rect 10081 39119 10116 39153
rect 10150 39119 10185 39153
rect 10219 39119 10254 39153
rect 10288 39119 10323 39153
rect 10357 39119 10392 39153
rect 10426 39119 10461 39153
rect 10495 39119 10530 39153
rect 10564 39119 10599 39153
rect 10633 39119 10668 39153
rect 10702 39119 10737 39153
rect 10771 39119 10806 39153
rect 10840 39119 10875 39153
rect 10909 39119 10944 39153
rect 10978 39119 11013 39153
rect 11047 39119 11082 39153
rect 11116 39119 11151 39153
rect 11185 39119 11220 39153
rect 11254 39119 11289 39153
rect 11323 39119 11358 39153
rect 11392 39119 11427 39153
rect 11461 39119 11496 39153
rect 11530 39119 11565 39153
rect 11599 39119 11634 39153
rect 11668 39119 11703 39153
rect 11737 39119 11772 39153
rect 11806 39119 11841 39153
rect 11875 39119 11910 39153
rect 11944 39119 11979 39153
rect 12013 39119 12048 39153
rect 12082 39119 12117 39153
rect 12151 39119 12186 39153
rect 12220 39119 12255 39153
rect 12289 39119 12324 39153
rect 12358 39119 12393 39153
rect 12427 39119 12462 39153
rect 12496 39119 12531 39153
rect 12565 39119 12600 39153
rect 12634 39119 12669 39153
rect 12703 39119 12738 39153
rect 12772 39119 12807 39153
rect 12841 39119 12876 39153
rect 12910 39119 12945 39153
rect 12979 39119 13014 39153
rect 13048 39119 13083 39153
rect 13117 39119 13152 39153
rect 13186 39119 13221 39153
rect 13255 39119 13290 39153
rect 13324 39119 13359 39153
rect 13393 39119 13428 39153
rect 13462 39129 13617 39153
rect 13462 39119 13515 39129
rect 2444 39027 13515 39119
rect 2444 38993 2482 39027
rect 2516 38993 2550 39027
rect 2584 38993 2618 39027
rect 2652 38993 2686 39027
rect 2720 38993 2754 39027
rect 2788 38993 2822 39027
rect 2856 38993 2890 39027
rect 2924 38993 2958 39027
rect 2992 38993 3026 39027
rect 3060 38993 3094 39027
rect 3128 38993 3162 39027
rect 3196 38993 3230 39027
rect 3264 38993 3298 39027
rect 3332 38993 3366 39027
rect 3400 38993 3434 39027
rect 3468 38993 3502 39027
rect 3536 38993 3570 39027
rect 3604 38993 3638 39027
rect 3672 38993 3706 39027
rect 3740 38993 3774 39027
rect 3808 38993 3842 39027
rect 3876 38993 3910 39027
rect 3944 38993 3978 39027
rect 4012 38993 4046 39027
rect 4080 38993 4114 39027
rect 4148 38993 4182 39027
rect 4216 38993 4250 39027
rect 4284 38993 4318 39027
rect 4352 38993 4386 39027
rect 4420 38993 4454 39027
rect 4488 38993 4522 39027
rect 4556 38993 4590 39027
rect 4624 38993 4658 39027
rect 4692 38993 4726 39027
rect 4760 38993 4794 39027
rect 4828 38993 4862 39027
rect 4896 38993 4930 39027
rect 4964 38993 4998 39027
rect 5032 38993 5066 39027
rect 5100 38993 5134 39027
rect 5168 38993 5202 39027
rect 5236 38993 5270 39027
rect 5304 38993 5338 39027
rect 5372 38993 5406 39027
rect 5440 38993 5474 39027
rect 5508 38993 5542 39027
rect 5576 38993 5610 39027
rect 5644 38993 5678 39027
rect 5712 38993 5746 39027
rect 5780 38993 5814 39027
rect 5848 38993 5882 39027
rect 5916 38993 5950 39027
rect 5984 38993 6018 39027
rect 6052 38993 6086 39027
rect 6120 38993 6154 39027
rect 6188 38993 6222 39027
rect 6256 38993 6290 39027
rect 6324 38993 6358 39027
rect 6392 38993 6426 39027
rect 6460 38993 6494 39027
rect 6528 38993 6562 39027
rect 6596 38993 6630 39027
rect 6664 38993 6698 39027
rect 6732 38993 6766 39027
rect 6800 38993 6834 39027
rect 6868 38993 6902 39027
rect 6936 38993 6970 39027
rect 7004 38993 7038 39027
rect 7072 38993 7106 39027
rect 7140 38993 7174 39027
rect 7208 38993 7242 39027
rect 7276 38993 7310 39027
rect 7344 38993 7378 39027
rect 7412 38993 7446 39027
rect 7480 38993 7514 39027
rect 7548 38993 7582 39027
rect 7616 38993 7650 39027
rect 7684 38993 7718 39027
rect 7752 38993 7786 39027
rect 7820 38993 7854 39027
rect 7888 38993 7922 39027
rect 7956 38993 7990 39027
rect 8024 38993 8058 39027
rect 8092 38993 8126 39027
rect 8160 38993 8194 39027
rect 8228 38993 8262 39027
rect 8296 38993 8330 39027
rect 8364 38993 8398 39027
rect 8432 38993 8466 39027
rect 8500 38993 8534 39027
rect 8568 38993 8602 39027
rect 8636 38993 8670 39027
rect 8704 38993 8738 39027
rect 8772 38993 8806 39027
rect 8840 38993 8874 39027
rect 8908 38993 8943 39027
rect 8977 38993 9012 39027
rect 9046 38993 9081 39027
rect 9115 38993 9150 39027
rect 9184 38993 9219 39027
rect 9253 38993 9288 39027
rect 9322 38993 9357 39027
rect 9391 38993 9426 39027
rect 9460 38993 9495 39027
rect 9529 38993 9564 39027
rect 9598 38993 9633 39027
rect 9667 38993 9702 39027
rect 9736 38993 9771 39027
rect 9805 38993 9840 39027
rect 9874 38993 9909 39027
rect 9943 38993 9978 39027
rect 10012 38993 10047 39027
rect 10081 38993 10116 39027
rect 10150 38993 10185 39027
rect 10219 38993 10254 39027
rect 10288 38993 10323 39027
rect 10357 38993 10392 39027
rect 10426 38993 10461 39027
rect 10495 38993 10530 39027
rect 10564 38993 10599 39027
rect 10633 38993 10668 39027
rect 10702 38993 10737 39027
rect 10771 38993 10806 39027
rect 10840 38993 10875 39027
rect 10909 38993 10944 39027
rect 10978 38993 11013 39027
rect 11047 38993 11082 39027
rect 11116 38993 11151 39027
rect 11185 38993 11220 39027
rect 11254 38993 11289 39027
rect 11323 38993 11358 39027
rect 11392 38993 11427 39027
rect 11461 38993 11496 39027
rect 11530 38993 11565 39027
rect 11599 38993 11634 39027
rect 11668 38993 11703 39027
rect 11737 38993 11772 39027
rect 11806 38993 11841 39027
rect 11875 38993 11910 39027
rect 11944 38993 11979 39027
rect 12013 38993 12048 39027
rect 12082 38993 12117 39027
rect 12151 38993 12186 39027
rect 12220 38993 12255 39027
rect 12289 38993 12324 39027
rect 12358 38993 12393 39027
rect 12427 38993 12462 39027
rect 12496 38993 12531 39027
rect 12565 38993 12600 39027
rect 12634 38993 12669 39027
rect 12703 38993 12738 39027
rect 12772 38993 12807 39027
rect 12841 38993 12876 39027
rect 12910 38993 12945 39027
rect 12979 38993 13014 39027
rect 13048 38993 13083 39027
rect 13117 38993 13152 39027
rect 13186 38993 13221 39027
rect 13255 38993 13290 39027
rect 13324 38993 13359 39027
rect 13393 38993 13428 39027
rect 13462 38993 13515 39027
rect 2376 29089 2444 29157
rect 2274 29063 2444 29089
rect 2274 29055 2410 29063
rect 2308 29021 2410 29055
rect 2274 28995 2410 29021
rect 4144 29029 4178 29063
rect 4212 29029 4298 29063
rect 4144 28995 4298 29029
rect 2274 28893 2342 28995
rect 4144 28961 4196 28995
rect 4076 28927 4196 28961
rect 4076 28893 4128 28927
rect 4298 23554 4335 23588
rect 4369 23554 4403 23588
rect 4437 23554 4471 23588
rect 4505 23554 4539 23588
rect 4573 23554 4607 23588
rect 4641 23554 4675 23588
rect 4709 23554 4743 23588
rect 4777 23554 4811 23588
rect 4845 23554 4879 23588
rect 4913 23554 4947 23588
rect 4981 23554 5015 23588
rect 5049 23554 5083 23588
rect 5117 23554 5151 23588
rect 5185 23554 5219 23588
rect 5253 23554 5287 23588
rect 5321 23554 5355 23588
rect 5389 23554 5423 23588
rect 5457 23554 5491 23588
rect 5525 23554 5559 23588
rect 5593 23554 5627 23588
rect 5661 23554 5695 23588
rect 5729 23554 5763 23588
rect 5797 23554 5831 23588
rect 5865 23554 5899 23588
rect 5933 23554 5967 23588
rect 6001 23554 6035 23588
rect 6069 23554 6103 23588
rect 6137 23554 6171 23588
rect 6205 23554 6239 23588
rect 6273 23554 6307 23588
rect 6341 23554 6375 23588
rect 6409 23554 6443 23588
rect 6477 23554 6511 23588
rect 6545 23554 6579 23588
rect 6613 23554 6647 23588
rect 6681 23554 6715 23588
rect 6749 23554 6783 23588
rect 6817 23554 6851 23588
rect 6885 23554 6919 23588
rect 6953 23554 6987 23588
rect 7021 23554 7055 23588
rect 7089 23554 7123 23588
rect 7157 23554 7191 23588
rect 7225 23554 7259 23588
rect 7293 23554 7327 23588
rect 7361 23554 7395 23588
rect 7429 23554 7463 23588
rect 7497 23554 7531 23588
rect 7565 23554 7599 23588
rect 7633 23554 7667 23588
rect 7701 23554 7735 23588
rect 7769 23554 7803 23588
rect 7837 23554 7871 23588
rect 7905 23554 7939 23588
rect 7973 23554 8007 23588
rect 8041 23554 8075 23588
rect 8109 23554 8143 23588
rect 8177 23554 8211 23588
rect 8245 23554 8279 23588
rect 8313 23554 8347 23588
rect 8381 23554 8415 23588
rect 8449 23554 8483 23588
rect 8517 23554 8551 23588
rect 8585 23554 8619 23588
rect 8653 23554 8687 23588
rect 8721 23554 8755 23588
rect 8789 23554 8823 23588
rect 8857 23554 8891 23588
rect 8925 23554 8959 23588
rect 8993 23554 9027 23588
rect 9061 23554 9095 23588
rect 9129 23554 9163 23588
rect 9197 23554 9231 23588
rect 9265 23554 9299 23588
rect 9333 23554 9367 23588
rect 9401 23554 9435 23588
rect 9469 23554 9503 23588
rect 9537 23554 9571 23588
rect 9605 23554 9639 23588
rect 9673 23554 9707 23588
rect 9741 23554 9775 23588
rect 9809 23554 9843 23588
rect 9877 23554 9911 23588
rect 9945 23554 9979 23588
rect 10013 23554 10047 23588
rect 10081 23554 10115 23588
rect 10149 23554 10183 23588
rect 10217 23554 10251 23588
rect 10285 23554 10319 23588
rect 10353 23554 10387 23588
rect 10421 23554 10455 23588
rect 10489 23554 10523 23588
rect 10557 23554 10591 23588
rect 10625 23554 10659 23588
rect 10693 23554 10727 23588
rect 10761 23554 10795 23588
rect 10829 23554 10863 23588
rect 10897 23554 10931 23588
rect 10965 23554 10999 23588
rect 11033 23554 11067 23588
rect 11101 23554 11135 23588
rect 11169 23554 11203 23588
rect 11237 23554 11271 23588
rect 11305 23554 11339 23588
rect 11373 23554 11407 23588
rect 11441 23554 11475 23588
rect 11509 23554 11543 23588
rect 11577 23554 11611 23588
rect 11645 23554 11679 23588
rect 11713 23554 11747 23588
rect 11781 23554 11815 23588
rect 11849 23554 11883 23588
rect 11917 23554 11951 23588
rect 11985 23554 12019 23588
rect 12053 23554 12087 23588
rect 12121 23554 12155 23588
rect 12189 23554 12223 23588
rect 12257 23554 12291 23588
rect 12325 23554 12359 23588
rect 12393 23554 12427 23588
rect 12461 23554 12495 23588
rect 12529 23554 12563 23588
rect 12597 23554 12631 23588
rect 12665 23554 12699 23588
rect 12733 23554 12767 23588
rect 12801 23554 12835 23588
rect 12869 23554 12903 23588
rect 12937 23554 12971 23588
rect 13005 23554 13039 23588
rect 13073 23554 13107 23588
rect 13141 23554 13175 23588
rect 13209 23554 13243 23588
rect 13277 23554 13311 23588
rect 13345 23554 13379 23588
rect 13413 23554 13447 23588
rect 13481 23554 13515 23588
rect 4298 21855 4335 21889
rect 4369 21855 4403 21889
rect 4437 21855 4471 21889
rect 4505 21855 4539 21889
rect 4573 21855 4607 21889
rect 4641 21855 4675 21889
rect 4709 21855 4743 21889
rect 4777 21855 4811 21889
rect 4845 21855 4879 21889
rect 4913 21855 4947 21889
rect 4981 21855 5015 21889
rect 5049 21855 5083 21889
rect 5117 21855 5151 21889
rect 5185 21855 5219 21889
rect 5253 21855 5287 21889
rect 5321 21855 5355 21889
rect 5389 21855 5423 21889
rect 5457 21855 5491 21889
rect 5525 21855 5559 21889
rect 5593 21855 5627 21889
rect 5661 21855 5695 21889
rect 5729 21855 5763 21889
rect 5797 21855 5831 21889
rect 5865 21855 5899 21889
rect 5933 21855 5967 21889
rect 6001 21855 6035 21889
rect 6069 21855 6103 21889
rect 6137 21855 6171 21889
rect 6205 21855 6239 21889
rect 6273 21855 6307 21889
rect 6341 21855 6375 21889
rect 6409 21855 6443 21889
rect 6477 21855 6511 21889
rect 6545 21855 6579 21889
rect 6613 21855 6647 21889
rect 6681 21855 6715 21889
rect 6749 21855 6783 21889
rect 6817 21855 6851 21889
rect 6885 21855 6919 21889
rect 6953 21855 6987 21889
rect 7021 21855 7055 21889
rect 7089 21855 7123 21889
rect 7157 21855 7191 21889
rect 7225 21855 7259 21889
rect 7293 21855 7327 21889
rect 7361 21855 7395 21889
rect 7429 21855 7463 21889
rect 7497 21855 7531 21889
rect 7565 21855 7599 21889
rect 7633 21855 7667 21889
rect 7701 21855 7735 21889
rect 7769 21855 7803 21889
rect 7837 21855 7871 21889
rect 7905 21855 7939 21889
rect 7973 21855 8007 21889
rect 8041 21855 8075 21889
rect 8109 21855 8143 21889
rect 8177 21855 8211 21889
rect 8245 21855 8279 21889
rect 8313 21855 8347 21889
rect 8381 21855 8415 21889
rect 8449 21855 8483 21889
rect 8517 21855 8551 21889
rect 8585 21855 8619 21889
rect 8653 21855 8687 21889
rect 8721 21855 8755 21889
rect 8789 21855 8823 21889
rect 8857 21855 8891 21889
rect 8925 21855 8959 21889
rect 8993 21855 9027 21889
rect 9061 21855 9095 21889
rect 9129 21855 9163 21889
rect 9197 21855 9231 21889
rect 9265 21855 9299 21889
rect 9333 21855 9367 21889
rect 9401 21855 9435 21889
rect 9469 21855 9503 21889
rect 9537 21855 9571 21889
rect 9605 21855 9639 21889
rect 9673 21855 9707 21889
rect 9741 21855 9775 21889
rect 9809 21855 9843 21889
rect 9877 21855 9911 21889
rect 9945 21855 9979 21889
rect 10013 21855 10047 21889
rect 10081 21855 10115 21889
rect 10149 21855 10183 21889
rect 10217 21855 10251 21889
rect 10285 21855 10319 21889
rect 10353 21855 10387 21889
rect 10421 21855 10455 21889
rect 10489 21855 10523 21889
rect 10557 21855 10591 21889
rect 10625 21855 10659 21889
rect 10693 21855 10727 21889
rect 10761 21855 10795 21889
rect 10829 21855 10863 21889
rect 10897 21855 10931 21889
rect 10965 21855 10999 21889
rect 11033 21855 11067 21889
rect 11101 21855 11135 21889
rect 11169 21855 11203 21889
rect 11237 21855 11271 21889
rect 11305 21855 11339 21889
rect 11373 21855 11407 21889
rect 11441 21855 11475 21889
rect 11509 21855 11543 21889
rect 11577 21855 11611 21889
rect 11645 21855 11679 21889
rect 11713 21855 11747 21889
rect 11781 21855 11815 21889
rect 11849 21855 11883 21889
rect 11917 21855 11951 21889
rect 11985 21855 12019 21889
rect 12053 21855 12087 21889
rect 12121 21855 12155 21889
rect 12189 21855 12223 21889
rect 12257 21855 12291 21889
rect 12325 21855 12359 21889
rect 12393 21855 12427 21889
rect 12461 21855 12495 21889
rect 12529 21855 12563 21889
rect 12597 21855 12631 21889
rect 12665 21855 12699 21889
rect 12733 21855 12767 21889
rect 12801 21855 12835 21889
rect 12869 21855 12903 21889
rect 12937 21855 12971 21889
rect 13005 21855 13039 21889
rect 13073 21855 13107 21889
rect 13141 21855 13175 21889
rect 13209 21855 13243 21889
rect 13277 21855 13311 21889
rect 13345 21855 13379 21889
rect 13413 21855 13447 21889
rect 13481 21855 13515 21889
rect 4128 20207 4298 20257
rect 13515 20496 13617 20531
rect 13549 20462 13583 20496
rect 13515 20427 13617 20462
rect 13549 20393 13583 20427
rect 13515 20358 13617 20393
rect 13549 20324 13583 20358
rect 13515 20289 13617 20324
rect 13549 20255 13583 20289
rect 13515 20207 13617 20255
rect 4128 20173 4152 20207
rect 4186 20173 4221 20207
rect 4255 20173 4290 20207
rect 4324 20173 4359 20207
rect 4393 20173 4428 20207
rect 4462 20173 4497 20207
rect 4531 20173 4566 20207
rect 4600 20173 4635 20207
rect 4669 20173 4704 20207
rect 4738 20173 4773 20207
rect 4807 20173 4842 20207
rect 4876 20173 4911 20207
rect 4945 20173 4980 20207
rect 5014 20173 5049 20207
rect 5083 20173 5118 20207
rect 5152 20173 5187 20207
rect 5221 20173 5256 20207
rect 5290 20173 5325 20207
rect 5359 20173 5394 20207
rect 5428 20173 5463 20207
rect 5497 20173 5532 20207
rect 5566 20173 5601 20207
rect 5635 20173 5670 20207
rect 5704 20173 5739 20207
rect 5773 20173 5807 20207
rect 5841 20173 5875 20207
rect 5909 20173 5943 20207
rect 5977 20173 6011 20207
rect 6045 20173 6079 20207
rect 6113 20173 6147 20207
rect 6181 20173 6215 20207
rect 6249 20173 6283 20207
rect 6317 20173 6351 20207
rect 6385 20173 6419 20207
rect 6453 20173 6487 20207
rect 6521 20173 6555 20207
rect 6589 20173 6623 20207
rect 6657 20173 6691 20207
rect 6725 20173 6759 20207
rect 6793 20173 6827 20207
rect 6861 20173 6895 20207
rect 6929 20173 6963 20207
rect 6997 20173 7031 20207
rect 7065 20173 7099 20207
rect 7133 20173 7167 20207
rect 7201 20173 7235 20207
rect 7269 20173 7303 20207
rect 7337 20173 7371 20207
rect 7405 20173 7439 20207
rect 7473 20173 7507 20207
rect 7541 20173 7575 20207
rect 7609 20173 7643 20207
rect 7677 20173 7711 20207
rect 7745 20173 7779 20207
rect 7813 20173 7847 20207
rect 7881 20173 7915 20207
rect 7949 20173 7983 20207
rect 8017 20173 8051 20207
rect 8085 20173 8119 20207
rect 8153 20173 8187 20207
rect 8221 20173 8255 20207
rect 8289 20173 8323 20207
rect 8357 20173 8391 20207
rect 8425 20173 8459 20207
rect 8493 20173 8527 20207
rect 8561 20173 8595 20207
rect 8629 20173 8663 20207
rect 8697 20173 8731 20207
rect 8765 20173 8799 20207
rect 8833 20173 8867 20207
rect 8901 20173 8935 20207
rect 8969 20173 9003 20207
rect 9037 20173 9071 20207
rect 9105 20173 9139 20207
rect 9173 20173 9207 20207
rect 9241 20173 9275 20207
rect 9309 20173 9343 20207
rect 9377 20173 9411 20207
rect 9445 20173 9479 20207
rect 9513 20173 9547 20207
rect 9581 20173 9615 20207
rect 9649 20173 9683 20207
rect 9717 20173 9751 20207
rect 9785 20173 9819 20207
rect 9853 20173 9887 20207
rect 9921 20173 9955 20207
rect 9989 20173 10023 20207
rect 10057 20173 10091 20207
rect 10125 20173 10159 20207
rect 10193 20173 10227 20207
rect 10261 20173 10295 20207
rect 10329 20173 10363 20207
rect 10397 20173 10431 20207
rect 10465 20173 10499 20207
rect 10533 20173 10567 20207
rect 10601 20173 10635 20207
rect 10669 20173 10703 20207
rect 10737 20173 10771 20207
rect 10805 20173 10839 20207
rect 10873 20173 10907 20207
rect 10941 20173 10975 20207
rect 11009 20173 11043 20207
rect 11077 20173 11111 20207
rect 11145 20173 11179 20207
rect 11213 20173 11247 20207
rect 11281 20173 11315 20207
rect 11349 20173 11383 20207
rect 11417 20173 11451 20207
rect 11485 20173 11519 20207
rect 11553 20173 11587 20207
rect 11621 20173 11655 20207
rect 11689 20173 11723 20207
rect 11757 20173 11791 20207
rect 11825 20173 11859 20207
rect 11893 20173 11927 20207
rect 11961 20173 11995 20207
rect 12029 20173 12063 20207
rect 12097 20173 12131 20207
rect 12165 20173 12199 20207
rect 12233 20173 12267 20207
rect 12301 20173 12335 20207
rect 12369 20173 12403 20207
rect 12437 20173 12471 20207
rect 12505 20173 12539 20207
rect 12573 20173 12607 20207
rect 12641 20173 12675 20207
rect 12709 20173 12743 20207
rect 12777 20173 12811 20207
rect 12845 20173 12879 20207
rect 12913 20173 12947 20207
rect 12981 20173 13015 20207
rect 13049 20173 13083 20207
rect 13117 20173 13151 20207
rect 13185 20173 13219 20207
rect 13253 20173 13287 20207
rect 13321 20173 13355 20207
rect 13389 20173 13423 20207
rect 13457 20173 13491 20207
rect 13525 20173 13559 20207
rect 13593 20173 13617 20207
rect 4554 19798 4578 19832
rect 4612 19798 4647 19832
rect 4681 19798 4716 19832
rect 4750 19798 4785 19832
rect 4819 19798 4854 19832
rect 4888 19798 4923 19832
rect 4957 19798 4992 19832
rect 5026 19798 5061 19832
rect 5095 19798 5130 19832
rect 5164 19798 5199 19832
rect 5233 19798 5268 19832
rect 5302 19798 5337 19832
rect 5371 19798 5406 19832
rect 5440 19798 5475 19832
rect 5509 19798 5544 19832
rect 5578 19798 5613 19832
rect 5647 19798 5682 19832
rect 5716 19798 5750 19832
rect 5784 19798 5818 19832
rect 5852 19798 5886 19832
rect 5920 19798 5954 19832
rect 5988 19798 6022 19832
rect 6056 19798 6090 19832
rect 6124 19798 6158 19832
rect 6192 19798 6226 19832
rect 6260 19798 6294 19832
rect 6328 19798 6362 19832
rect 6396 19798 6430 19832
rect 6464 19798 6498 19832
rect 6532 19798 6566 19832
rect 6600 19798 6634 19832
rect 6668 19798 6702 19832
rect 6736 19798 6770 19832
rect 6804 19798 6838 19832
rect 6872 19798 6906 19832
rect 6940 19798 6974 19832
rect 7008 19798 7042 19832
rect 7076 19798 7110 19832
rect 7144 19798 7178 19832
rect 7212 19798 7246 19832
rect 7280 19798 7314 19832
rect 7348 19798 7382 19832
rect 7416 19798 7450 19832
rect 7484 19798 7518 19832
rect 7552 19798 7586 19832
rect 7620 19798 7654 19832
rect 7688 19798 7722 19832
rect 7756 19798 7790 19832
rect 7824 19798 7858 19832
rect 7892 19798 7926 19832
rect 7960 19798 7994 19832
rect 8028 19798 8062 19832
rect 8096 19798 8130 19832
rect 8164 19798 8198 19832
rect 8232 19798 8266 19832
rect 8300 19798 8334 19832
rect 8368 19798 8402 19832
rect 8436 19798 8470 19832
rect 8504 19798 8538 19832
rect 8572 19798 8606 19832
rect 8640 19798 8674 19832
rect 8708 19798 8742 19832
rect 8776 19798 8810 19832
rect 8844 19798 8878 19832
rect 8912 19798 8946 19832
rect 8980 19798 9014 19832
rect 9048 19798 9082 19832
rect 9116 19798 9150 19832
rect 9184 19798 9218 19832
rect 9252 19798 9286 19832
rect 9320 19798 9354 19832
rect 9388 19798 9422 19832
rect 9456 19798 9490 19832
rect 9524 19798 9558 19832
rect 9592 19798 9626 19832
rect 9660 19798 9694 19832
rect 9728 19798 9762 19832
rect 9796 19798 9830 19832
rect 9864 19798 9898 19832
rect 9932 19798 9966 19832
rect 10000 19798 10034 19832
rect 10068 19798 10102 19832
rect 10136 19798 10170 19832
rect 10204 19798 10238 19832
rect 10272 19798 10306 19832
rect 10340 19798 10374 19832
rect 10408 19798 10442 19832
rect 10476 19798 10510 19832
rect 10544 19798 10578 19832
rect 10612 19798 10646 19832
rect 10680 19798 10714 19832
rect 10748 19798 10782 19832
rect 10816 19798 10850 19832
rect 10884 19798 10918 19832
rect 10952 19798 10986 19832
rect 11020 19798 11054 19832
rect 11088 19798 11122 19832
rect 11156 19798 11190 19832
rect 11224 19798 11258 19832
rect 11292 19798 11326 19832
rect 11360 19798 11394 19832
rect 11428 19798 11462 19832
rect 11496 19798 11530 19832
rect 11564 19798 11598 19832
rect 11632 19798 11666 19832
rect 11700 19798 11734 19832
rect 11768 19798 11802 19832
rect 11836 19798 11870 19832
rect 11904 19798 11938 19832
rect 11972 19798 12006 19832
rect 12040 19798 12074 19832
rect 12108 19798 12142 19832
rect 12176 19798 12210 19832
rect 12244 19798 12278 19832
rect 12312 19798 12346 19832
rect 12380 19798 12414 19832
rect 12448 19798 12482 19832
rect 12516 19798 12550 19832
rect 12584 19798 12618 19832
rect 12652 19798 12686 19832
rect 12720 19798 12754 19832
rect 12788 19798 12822 19832
rect 12856 19798 12890 19832
rect 12924 19798 12958 19832
rect 12992 19798 13026 19832
rect 13060 19798 13094 19832
rect 13128 19798 13162 19832
rect 13196 19798 13230 19832
rect 13264 19798 13298 19832
rect 13332 19798 13366 19832
rect 13400 19798 13434 19832
rect 13468 19798 13502 19832
rect 13536 19798 13570 19832
rect 13604 19798 13628 19832
rect 4554 19764 4656 19798
rect 13458 19701 13628 19798
rect 4656 18135 4754 18169
rect 4788 18135 4822 18169
rect 4856 18135 4890 18169
rect 4924 18135 4958 18169
rect 4992 18135 5026 18169
rect 5060 18135 5094 18169
rect 5128 18135 5162 18169
rect 5196 18135 5230 18169
rect 5264 18135 5298 18169
rect 5332 18135 5366 18169
rect 5400 18135 5434 18169
rect 5468 18135 5502 18169
rect 5536 18135 5570 18169
rect 5604 18135 5638 18169
rect 5672 18135 5706 18169
rect 5740 18135 5774 18169
rect 5808 18135 5842 18169
rect 5876 18135 5910 18169
rect 5944 18135 5978 18169
rect 6012 18135 6046 18169
rect 6080 18135 6114 18169
rect 6148 18135 6182 18169
rect 6216 18135 6250 18169
rect 6284 18135 6318 18169
rect 6352 18135 6386 18169
rect 6420 18135 6454 18169
rect 6488 18135 6522 18169
rect 6556 18135 6590 18169
rect 6624 18135 6658 18169
rect 6692 18135 6726 18169
rect 6760 18135 6794 18169
rect 6828 18135 6862 18169
rect 6896 18135 6930 18169
rect 6964 18135 6998 18169
rect 7032 18135 7066 18169
rect 7100 18135 7134 18169
rect 7168 18135 7202 18169
rect 7236 18135 7270 18169
rect 7304 18135 7338 18169
rect 7372 18135 7406 18169
rect 7440 18135 7474 18169
rect 7508 18135 7542 18169
rect 7576 18135 7610 18169
rect 7644 18135 7678 18169
rect 7712 18135 7746 18169
rect 7780 18135 7814 18169
rect 7848 18135 7882 18169
rect 7916 18135 7950 18169
rect 7984 18135 8018 18169
rect 8052 18135 8086 18169
rect 8120 18135 8154 18169
rect 8188 18135 8222 18169
rect 8256 18135 8290 18169
rect 8324 18135 8358 18169
rect 8392 18135 8426 18169
rect 8460 18135 8494 18169
rect 8528 18135 8562 18169
rect 8596 18135 8630 18169
rect 8664 18135 8698 18169
rect 8732 18135 8766 18169
rect 8800 18135 8834 18169
rect 8868 18135 8902 18169
rect 8936 18135 8970 18169
rect 9004 18135 9038 18169
rect 9072 18135 9106 18169
rect 9140 18135 9174 18169
rect 9208 18135 9242 18169
rect 9276 18135 9310 18169
rect 9344 18135 9378 18169
rect 9412 18135 9446 18169
rect 9480 18135 9514 18169
rect 9548 18135 9582 18169
rect 9616 18135 9650 18169
rect 9684 18135 9718 18169
rect 9752 18135 9786 18169
rect 9820 18135 9854 18169
rect 9888 18135 9922 18169
rect 9956 18135 9990 18169
rect 10024 18135 10058 18169
rect 10092 18135 10126 18169
rect 10160 18135 10194 18169
rect 10228 18135 10262 18169
rect 10296 18135 10330 18169
rect 10364 18135 10398 18169
rect 10432 18135 10466 18169
rect 10500 18135 10534 18169
rect 10568 18135 10602 18169
rect 10636 18135 10670 18169
rect 10704 18135 10738 18169
rect 10772 18135 10806 18169
rect 10840 18135 10874 18169
rect 10908 18135 10942 18169
rect 10976 18135 11010 18169
rect 11044 18135 11078 18169
rect 11112 18135 11146 18169
rect 11180 18135 11214 18169
rect 11248 18135 11282 18169
rect 11316 18135 11350 18169
rect 11384 18135 11418 18169
rect 11452 18135 11486 18169
rect 11520 18135 11554 18169
rect 11588 18135 11622 18169
rect 11656 18135 11690 18169
rect 11724 18135 11758 18169
rect 11792 18135 11826 18169
rect 11860 18135 11894 18169
rect 11928 18135 11962 18169
rect 11996 18135 12030 18169
rect 12064 18135 12098 18169
rect 12132 18135 12166 18169
rect 12200 18135 12234 18169
rect 12268 18135 12302 18169
rect 12336 18135 12370 18169
rect 12404 18135 12438 18169
rect 12472 18135 12506 18169
rect 12540 18135 12574 18169
rect 12608 18135 12642 18169
rect 12676 18135 12710 18169
rect 12744 18135 12778 18169
rect 12812 18135 12846 18169
rect 12880 18135 12914 18169
rect 12948 18135 12982 18169
rect 13016 18135 13050 18169
rect 13084 18135 13118 18169
rect 13152 18135 13186 18169
rect 13220 18135 13254 18169
rect 13288 18135 13322 18169
rect 13356 18135 13390 18169
rect 13424 18135 13458 18169
rect 4656 16466 4754 16470
rect 4554 16436 4754 16466
rect 4788 16436 4822 16470
rect 4856 16436 4890 16470
rect 4924 16436 4958 16470
rect 4992 16436 5026 16470
rect 5060 16436 5094 16470
rect 5128 16436 5162 16470
rect 5196 16436 5230 16470
rect 5264 16436 5298 16470
rect 5332 16436 5366 16470
rect 5400 16436 5434 16470
rect 5468 16436 5502 16470
rect 5536 16436 5570 16470
rect 5604 16436 5638 16470
rect 5672 16436 5706 16470
rect 5740 16436 5774 16470
rect 5808 16436 5842 16470
rect 5876 16436 5910 16470
rect 5944 16436 5978 16470
rect 6012 16436 6046 16470
rect 6080 16436 6114 16470
rect 6148 16436 6182 16470
rect 6216 16436 6250 16470
rect 6284 16436 6318 16470
rect 6352 16436 6386 16470
rect 6420 16436 6454 16470
rect 6488 16436 6522 16470
rect 6556 16436 6590 16470
rect 6624 16436 6658 16470
rect 6692 16436 6726 16470
rect 6760 16436 6794 16470
rect 6828 16436 6862 16470
rect 6896 16436 6930 16470
rect 6964 16436 6998 16470
rect 7032 16436 7066 16470
rect 7100 16436 7134 16470
rect 7168 16436 7202 16470
rect 7236 16436 7270 16470
rect 7304 16436 7338 16470
rect 7372 16436 7406 16470
rect 7440 16436 7474 16470
rect 7508 16436 7542 16470
rect 7576 16436 7610 16470
rect 7644 16436 7678 16470
rect 7712 16436 7746 16470
rect 7780 16436 7814 16470
rect 7848 16436 7882 16470
rect 7916 16436 7950 16470
rect 7984 16436 8018 16470
rect 8052 16436 8086 16470
rect 8120 16436 8154 16470
rect 8188 16436 8222 16470
rect 8256 16436 8290 16470
rect 8324 16436 8358 16470
rect 8392 16436 8426 16470
rect 8460 16436 8494 16470
rect 8528 16436 8562 16470
rect 8596 16436 8630 16470
rect 8664 16436 8698 16470
rect 8732 16436 8766 16470
rect 8800 16436 8834 16470
rect 8868 16436 8902 16470
rect 8936 16436 8970 16470
rect 9004 16436 9038 16470
rect 9072 16436 9106 16470
rect 9140 16436 9174 16470
rect 9208 16436 9242 16470
rect 9276 16436 9310 16470
rect 9344 16436 9378 16470
rect 9412 16436 9446 16470
rect 9480 16436 9514 16470
rect 9548 16436 9582 16470
rect 9616 16436 9650 16470
rect 9684 16436 9718 16470
rect 9752 16436 9786 16470
rect 9820 16436 9854 16470
rect 9888 16436 9922 16470
rect 9956 16436 9990 16470
rect 10024 16436 10058 16470
rect 10092 16436 10126 16470
rect 10160 16436 10194 16470
rect 10228 16436 10262 16470
rect 10296 16436 10330 16470
rect 10364 16436 10398 16470
rect 10432 16436 10466 16470
rect 10500 16436 10534 16470
rect 10568 16436 10602 16470
rect 10636 16436 10670 16470
rect 10704 16436 10738 16470
rect 10772 16436 10806 16470
rect 10840 16436 10874 16470
rect 10908 16436 10942 16470
rect 10976 16436 11010 16470
rect 11044 16436 11078 16470
rect 11112 16436 11146 16470
rect 11180 16436 11214 16470
rect 11248 16436 11282 16470
rect 11316 16436 11350 16470
rect 11384 16436 11418 16470
rect 11452 16436 11486 16470
rect 11520 16436 11554 16470
rect 11588 16436 11622 16470
rect 11656 16436 11690 16470
rect 11724 16436 11758 16470
rect 11792 16436 11826 16470
rect 11860 16436 11894 16470
rect 11928 16436 11962 16470
rect 11996 16436 12030 16470
rect 12064 16436 12098 16470
rect 12132 16436 12166 16470
rect 12200 16436 12234 16470
rect 12268 16436 12302 16470
rect 12336 16436 12370 16470
rect 12404 16436 12438 16470
rect 12472 16436 12506 16470
rect 12540 16436 12574 16470
rect 12608 16436 12642 16470
rect 12676 16436 12710 16470
rect 12744 16436 12778 16470
rect 12812 16436 12846 16470
rect 12880 16436 12914 16470
rect 12948 16436 12982 16470
rect 13016 16436 13050 16470
rect 13084 16436 13118 16470
rect 13152 16436 13186 16470
rect 13220 16436 13254 16470
rect 13288 16436 13322 16470
rect 13356 16436 13390 16470
rect 13424 16436 13458 16470
rect 4554 16432 4656 16436
rect 4554 16417 4622 16432
rect 2274 16383 2514 16417
rect 2444 16315 2514 16383
rect 4588 16398 4622 16417
rect 4588 16315 4656 16398
rect 2274 5081 2478 5129
rect 13392 5115 13458 5183
rect 13392 5081 13628 5115
rect 1669 3646 3413 3670
rect 1669 3612 1677 3646
rect 1711 3612 1747 3646
rect 1781 3612 1817 3646
rect 1851 3612 1887 3646
rect 1921 3612 1957 3646
rect 1991 3612 2027 3646
rect 2061 3612 2097 3646
rect 2131 3612 2167 3646
rect 2201 3612 2237 3646
rect 2271 3612 2307 3646
rect 2341 3612 2377 3646
rect 2411 3612 2447 3646
rect 2481 3612 2517 3646
rect 2551 3612 2587 3646
rect 2621 3612 2657 3646
rect 2691 3612 2727 3646
rect 2761 3612 2797 3646
rect 2831 3612 2867 3646
rect 2901 3612 2937 3646
rect 2971 3612 3007 3646
rect 3041 3612 3077 3646
rect 3111 3612 3147 3646
rect 3181 3612 3217 3646
rect 3251 3612 3287 3646
rect 3321 3612 3413 3646
rect 1669 3578 3413 3612
rect 1669 3544 1677 3578
rect 1711 3544 1747 3578
rect 1781 3544 1817 3578
rect 1851 3544 1887 3578
rect 1921 3544 1957 3578
rect 1991 3544 2027 3578
rect 2061 3544 2097 3578
rect 2131 3544 2167 3578
rect 2201 3544 2237 3578
rect 2271 3544 2307 3578
rect 2341 3544 2377 3578
rect 2411 3544 2447 3578
rect 2481 3544 2517 3578
rect 2551 3544 2587 3578
rect 2621 3544 2657 3578
rect 2691 3544 2727 3578
rect 2761 3544 2797 3578
rect 2831 3544 2867 3578
rect 2901 3544 2937 3578
rect 2971 3544 3007 3578
rect 3041 3544 3077 3578
rect 3111 3544 3147 3578
rect 3181 3544 3217 3578
rect 3251 3544 3287 3578
rect 3321 3544 3413 3578
rect 1669 3510 3413 3544
rect 1669 3476 1677 3510
rect 1711 3476 1747 3510
rect 1781 3476 1817 3510
rect 1851 3476 1887 3510
rect 1921 3476 1957 3510
rect 1991 3476 2027 3510
rect 2061 3476 2097 3510
rect 2131 3476 2167 3510
rect 2201 3476 2237 3510
rect 2271 3476 2307 3510
rect 2341 3476 2377 3510
rect 2411 3476 2447 3510
rect 2481 3476 2517 3510
rect 2551 3476 2587 3510
rect 2621 3476 2657 3510
rect 2691 3476 2727 3510
rect 2761 3476 2797 3510
rect 2831 3476 2867 3510
rect 2901 3476 2937 3510
rect 2971 3476 3007 3510
rect 3041 3476 3077 3510
rect 3111 3476 3147 3510
rect 3181 3476 3217 3510
rect 3251 3476 3287 3510
rect 3321 3476 3413 3510
rect 1669 3442 3413 3476
rect 1669 3408 1677 3442
rect 1711 3408 1747 3442
rect 1781 3408 1817 3442
rect 1851 3408 1887 3442
rect 1921 3408 1957 3442
rect 1991 3408 2027 3442
rect 2061 3408 2097 3442
rect 2131 3408 2167 3442
rect 2201 3408 2237 3442
rect 2271 3408 2307 3442
rect 2341 3408 2377 3442
rect 2411 3408 2447 3442
rect 2481 3408 2517 3442
rect 2551 3408 2587 3442
rect 2621 3408 2657 3442
rect 2691 3408 2727 3442
rect 2761 3408 2797 3442
rect 2831 3408 2867 3442
rect 2901 3408 2937 3442
rect 2971 3408 3007 3442
rect 3041 3408 3077 3442
rect 3111 3408 3147 3442
rect 3181 3408 3217 3442
rect 3251 3408 3287 3442
rect 3321 3408 3413 3442
rect 1669 3374 3413 3408
rect 1669 3340 1677 3374
rect 1711 3340 1747 3374
rect 1781 3340 1817 3374
rect 1851 3340 1887 3374
rect 1921 3340 1957 3374
rect 1991 3340 2027 3374
rect 2061 3340 2097 3374
rect 2131 3340 2167 3374
rect 2201 3340 2237 3374
rect 2271 3340 2307 3374
rect 2341 3340 2377 3374
rect 2411 3340 2447 3374
rect 2481 3340 2517 3374
rect 2551 3340 2587 3374
rect 2621 3340 2657 3374
rect 2691 3340 2727 3374
rect 2761 3340 2797 3374
rect 2831 3340 2867 3374
rect 2901 3340 2937 3374
rect 2971 3340 3007 3374
rect 3041 3340 3077 3374
rect 3111 3340 3147 3374
rect 3181 3340 3217 3374
rect 3251 3340 3287 3374
rect 3321 3340 3413 3374
rect 1669 3306 3413 3340
rect 1669 3272 1677 3306
rect 1711 3272 1747 3306
rect 1781 3272 1817 3306
rect 1851 3272 1887 3306
rect 1921 3272 1957 3306
rect 1991 3272 2027 3306
rect 2061 3272 2097 3306
rect 2131 3272 2167 3306
rect 2201 3272 2237 3306
rect 2271 3272 2307 3306
rect 2341 3272 2377 3306
rect 2411 3272 2447 3306
rect 2481 3272 2517 3306
rect 2551 3272 2587 3306
rect 2621 3272 2657 3306
rect 2691 3272 2727 3306
rect 2761 3272 2797 3306
rect 2831 3272 2867 3306
rect 2901 3272 2937 3306
rect 2971 3272 3007 3306
rect 3041 3272 3077 3306
rect 3111 3272 3147 3306
rect 3181 3272 3217 3306
rect 3251 3272 3287 3306
rect 3321 3272 3413 3306
rect 1669 3238 3413 3272
rect 1669 3204 1677 3238
rect 1711 3204 1747 3238
rect 1781 3204 1817 3238
rect 1851 3204 1887 3238
rect 1921 3204 1957 3238
rect 1991 3204 2027 3238
rect 2061 3204 2097 3238
rect 2131 3204 2167 3238
rect 2201 3204 2237 3238
rect 2271 3204 2307 3238
rect 2341 3204 2377 3238
rect 2411 3204 2447 3238
rect 2481 3204 2517 3238
rect 2551 3204 2587 3238
rect 2621 3204 2657 3238
rect 2691 3204 2727 3238
rect 2761 3204 2797 3238
rect 2831 3204 2867 3238
rect 2901 3204 2937 3238
rect 2971 3204 3007 3238
rect 3041 3204 3077 3238
rect 3111 3204 3147 3238
rect 3181 3204 3217 3238
rect 3251 3204 3287 3238
rect 3321 3204 3413 3238
rect 1669 3169 3413 3204
rect 1669 3135 1677 3169
rect 1711 3135 1747 3169
rect 1781 3135 1817 3169
rect 1851 3135 1887 3169
rect 1921 3135 1957 3169
rect 1991 3135 2027 3169
rect 2061 3135 2097 3169
rect 2131 3135 2167 3169
rect 2201 3135 2237 3169
rect 2271 3135 2307 3169
rect 2341 3135 2377 3169
rect 2411 3135 2447 3169
rect 2481 3135 2517 3169
rect 2551 3135 2587 3169
rect 2621 3135 2657 3169
rect 2691 3135 2727 3169
rect 2761 3135 2797 3169
rect 2831 3135 2867 3169
rect 2901 3135 2937 3169
rect 2971 3135 3007 3169
rect 3041 3135 3077 3169
rect 3111 3135 3147 3169
rect 3181 3135 3217 3169
rect 3251 3135 3287 3169
rect 3321 3135 3413 3169
rect 1669 3100 3413 3135
rect 1669 3066 1677 3100
rect 1711 3066 1747 3100
rect 1781 3066 1817 3100
rect 1851 3066 1887 3100
rect 1921 3066 1957 3100
rect 1991 3066 2027 3100
rect 2061 3066 2097 3100
rect 2131 3066 2167 3100
rect 2201 3066 2237 3100
rect 2271 3066 2307 3100
rect 2341 3066 2377 3100
rect 2411 3066 2447 3100
rect 2481 3066 2517 3100
rect 2551 3066 2587 3100
rect 2621 3066 2657 3100
rect 2691 3066 2727 3100
rect 2761 3066 2797 3100
rect 2831 3066 2867 3100
rect 2901 3066 2937 3100
rect 2971 3066 3007 3100
rect 3041 3066 3077 3100
rect 3111 3066 3147 3100
rect 3181 3066 3217 3100
rect 3251 3066 3287 3100
rect 3321 3066 3413 3100
rect 1669 3031 3413 3066
rect 1669 2997 1677 3031
rect 1711 2997 1747 3031
rect 1781 2997 1817 3031
rect 1851 2997 1887 3031
rect 1921 2997 1957 3031
rect 1991 2997 2027 3031
rect 2061 2997 2097 3031
rect 2131 2997 2167 3031
rect 2201 2997 2237 3031
rect 2271 2997 2307 3031
rect 2341 2997 2377 3031
rect 2411 2997 2447 3031
rect 2481 2997 2517 3031
rect 2551 2997 2587 3031
rect 2621 2997 2657 3031
rect 2691 2997 2727 3031
rect 2761 2997 2797 3031
rect 2831 2997 2867 3031
rect 2901 2997 2937 3031
rect 2971 2997 3007 3031
rect 3041 2997 3077 3031
rect 3111 2997 3147 3031
rect 3181 2997 3217 3031
rect 3251 2997 3287 3031
rect 3321 2997 3413 3031
rect 1669 2962 3413 2997
rect 1669 2928 1677 2962
rect 1711 2928 1747 2962
rect 1781 2928 1817 2962
rect 1851 2928 1887 2962
rect 1921 2928 1957 2962
rect 1991 2928 2027 2962
rect 2061 2928 2097 2962
rect 2131 2928 2167 2962
rect 2201 2928 2237 2962
rect 2271 2928 2307 2962
rect 2341 2928 2377 2962
rect 2411 2928 2447 2962
rect 2481 2928 2517 2962
rect 2551 2928 2587 2962
rect 2621 2928 2657 2962
rect 2691 2928 2727 2962
rect 2761 2928 2797 2962
rect 2831 2928 2867 2962
rect 2901 2928 2937 2962
rect 2971 2928 3007 2962
rect 3041 2928 3077 2962
rect 3111 2928 3147 2962
rect 3181 2928 3217 2962
rect 3251 2928 3287 2962
rect 3321 2928 3413 2962
rect 1669 2893 3413 2928
rect 1669 2859 1677 2893
rect 1711 2859 1747 2893
rect 1781 2859 1817 2893
rect 1851 2859 1887 2893
rect 1921 2859 1957 2893
rect 1991 2859 2027 2893
rect 2061 2859 2097 2893
rect 2131 2859 2167 2893
rect 2201 2859 2237 2893
rect 2271 2859 2307 2893
rect 2341 2859 2377 2893
rect 2411 2859 2447 2893
rect 2481 2859 2517 2893
rect 2551 2859 2587 2893
rect 2621 2859 2657 2893
rect 2691 2859 2727 2893
rect 2761 2859 2797 2893
rect 2831 2859 2867 2893
rect 2901 2859 2937 2893
rect 2971 2859 3007 2893
rect 3041 2859 3077 2893
rect 3111 2859 3147 2893
rect 3181 2859 3217 2893
rect 3251 2859 3287 2893
rect 3321 2859 3413 2893
rect 1669 2824 3413 2859
rect 1669 2790 1677 2824
rect 1711 2790 1747 2824
rect 1781 2790 1817 2824
rect 1851 2790 1887 2824
rect 1921 2790 1957 2824
rect 1991 2790 2027 2824
rect 2061 2790 2097 2824
rect 2131 2790 2167 2824
rect 2201 2790 2237 2824
rect 2271 2790 2307 2824
rect 2341 2790 2377 2824
rect 2411 2790 2447 2824
rect 2481 2790 2517 2824
rect 2551 2790 2587 2824
rect 2621 2790 2657 2824
rect 2691 2790 2727 2824
rect 2761 2790 2797 2824
rect 2831 2790 2867 2824
rect 2901 2790 2937 2824
rect 2971 2790 3007 2824
rect 3041 2790 3077 2824
rect 3111 2790 3147 2824
rect 3181 2790 3217 2824
rect 3251 2790 3287 2824
rect 3321 2790 3413 2824
rect 1669 2755 3413 2790
rect 1669 2721 1677 2755
rect 1711 2721 1747 2755
rect 1781 2721 1817 2755
rect 1851 2721 1887 2755
rect 1921 2721 1957 2755
rect 1991 2721 2027 2755
rect 2061 2721 2097 2755
rect 2131 2721 2167 2755
rect 2201 2721 2237 2755
rect 2271 2721 2307 2755
rect 2341 2721 2377 2755
rect 2411 2721 2447 2755
rect 2481 2721 2517 2755
rect 2551 2721 2587 2755
rect 2621 2721 2657 2755
rect 2691 2721 2727 2755
rect 2761 2721 2797 2755
rect 2831 2721 2867 2755
rect 2901 2721 2937 2755
rect 2971 2721 3007 2755
rect 3041 2721 3077 2755
rect 3111 2721 3147 2755
rect 3181 2721 3217 2755
rect 3251 2721 3287 2755
rect 3321 2721 3413 2755
rect 1669 2686 3413 2721
rect 1669 2652 1677 2686
rect 1711 2652 1747 2686
rect 1781 2652 1817 2686
rect 1851 2652 1887 2686
rect 1921 2652 1957 2686
rect 1991 2652 2027 2686
rect 2061 2652 2097 2686
rect 2131 2652 2167 2686
rect 2201 2652 2237 2686
rect 2271 2652 2307 2686
rect 2341 2652 2377 2686
rect 2411 2652 2447 2686
rect 2481 2652 2517 2686
rect 2551 2652 2587 2686
rect 2621 2652 2657 2686
rect 2691 2652 2727 2686
rect 2761 2652 2797 2686
rect 2831 2652 2867 2686
rect 2901 2652 2937 2686
rect 2971 2652 3007 2686
rect 3041 2652 3077 2686
rect 3111 2652 3147 2686
rect 3181 2652 3217 2686
rect 3251 2652 3287 2686
rect 3321 2652 3413 2686
rect 1669 2617 3413 2652
rect 1669 2583 1677 2617
rect 1711 2583 1747 2617
rect 1781 2583 1817 2617
rect 1851 2583 1887 2617
rect 1921 2583 1957 2617
rect 1991 2583 2027 2617
rect 2061 2583 2097 2617
rect 2131 2583 2167 2617
rect 2201 2583 2237 2617
rect 2271 2583 2307 2617
rect 2341 2583 2377 2617
rect 2411 2583 2447 2617
rect 2481 2583 2517 2617
rect 2551 2583 2587 2617
rect 2621 2583 2657 2617
rect 2691 2583 2727 2617
rect 2761 2583 2797 2617
rect 2831 2583 2867 2617
rect 2901 2583 2937 2617
rect 2971 2583 3007 2617
rect 3041 2583 3077 2617
rect 3111 2583 3147 2617
rect 3181 2583 3217 2617
rect 3251 2583 3287 2617
rect 3321 2583 3413 2617
rect 1669 2548 3413 2583
rect 1669 2514 1677 2548
rect 1711 2514 1747 2548
rect 1781 2514 1817 2548
rect 1851 2514 1887 2548
rect 1921 2514 1957 2548
rect 1991 2514 2027 2548
rect 2061 2514 2097 2548
rect 2131 2514 2167 2548
rect 2201 2514 2237 2548
rect 2271 2514 2307 2548
rect 2341 2514 2377 2548
rect 2411 2514 2447 2548
rect 2481 2514 2517 2548
rect 2551 2514 2587 2548
rect 2621 2514 2657 2548
rect 2691 2514 2727 2548
rect 2761 2514 2797 2548
rect 2831 2514 2867 2548
rect 2901 2514 2937 2548
rect 2971 2514 3007 2548
rect 3041 2514 3077 2548
rect 3111 2514 3147 2548
rect 3181 2514 3217 2548
rect 3251 2514 3287 2548
rect 3321 2514 3413 2548
rect 1669 2479 3413 2514
rect 1669 2445 1677 2479
rect 1711 2445 1747 2479
rect 1781 2445 1817 2479
rect 1851 2445 1887 2479
rect 1921 2445 1957 2479
rect 1991 2445 2027 2479
rect 2061 2445 2097 2479
rect 2131 2445 2167 2479
rect 2201 2445 2237 2479
rect 2271 2445 2307 2479
rect 2341 2445 2377 2479
rect 2411 2445 2447 2479
rect 2481 2445 2517 2479
rect 2551 2445 2587 2479
rect 2621 2445 2657 2479
rect 2691 2445 2727 2479
rect 2761 2445 2797 2479
rect 2831 2445 2867 2479
rect 2901 2445 2937 2479
rect 2971 2445 3007 2479
rect 3041 2445 3077 2479
rect 3111 2445 3147 2479
rect 3181 2445 3217 2479
rect 3251 2445 3287 2479
rect 3321 2445 3413 2479
rect 1669 2410 3413 2445
rect 1669 2376 1677 2410
rect 1711 2376 1747 2410
rect 1781 2376 1817 2410
rect 1851 2376 1887 2410
rect 1921 2376 1957 2410
rect 1991 2376 2027 2410
rect 2061 2376 2097 2410
rect 2131 2376 2167 2410
rect 2201 2376 2237 2410
rect 2271 2376 2307 2410
rect 2341 2376 2377 2410
rect 2411 2376 2447 2410
rect 2481 2376 2517 2410
rect 2551 2376 2587 2410
rect 2621 2376 2657 2410
rect 2691 2376 2727 2410
rect 2761 2376 2797 2410
rect 2831 2376 2867 2410
rect 2901 2376 2937 2410
rect 2971 2376 3007 2410
rect 3041 2376 3077 2410
rect 3111 2376 3147 2410
rect 3181 2376 3217 2410
rect 3251 2376 3287 2410
rect 3321 2376 3413 2410
rect 1669 2341 3413 2376
rect 1669 2307 1677 2341
rect 1711 2307 1747 2341
rect 1781 2307 1817 2341
rect 1851 2307 1887 2341
rect 1921 2307 1957 2341
rect 1991 2307 2027 2341
rect 2061 2307 2097 2341
rect 2131 2307 2167 2341
rect 2201 2307 2237 2341
rect 2271 2307 2307 2341
rect 2341 2307 2377 2341
rect 2411 2307 2447 2341
rect 2481 2307 2517 2341
rect 2551 2307 2587 2341
rect 2621 2307 2657 2341
rect 2691 2307 2727 2341
rect 2761 2307 2797 2341
rect 2831 2307 2867 2341
rect 2901 2307 2937 2341
rect 2971 2307 3007 2341
rect 3041 2307 3077 2341
rect 3111 2307 3147 2341
rect 3181 2307 3217 2341
rect 3251 2307 3287 2341
rect 3321 2307 3413 2341
rect 1669 2272 3413 2307
rect 1669 2238 1677 2272
rect 1711 2238 1747 2272
rect 1781 2238 1817 2272
rect 1851 2238 1887 2272
rect 1921 2238 1957 2272
rect 1991 2238 2027 2272
rect 2061 2238 2097 2272
rect 2131 2238 2167 2272
rect 2201 2238 2237 2272
rect 2271 2238 2307 2272
rect 2341 2238 2377 2272
rect 2411 2238 2447 2272
rect 2481 2238 2517 2272
rect 2551 2238 2587 2272
rect 2621 2238 2657 2272
rect 2691 2238 2727 2272
rect 2761 2238 2797 2272
rect 2831 2238 2867 2272
rect 2901 2238 2937 2272
rect 2971 2238 3007 2272
rect 3041 2238 3077 2272
rect 3111 2238 3147 2272
rect 3181 2238 3217 2272
rect 3251 2238 3287 2272
rect 3321 2238 3413 2272
rect 1669 2203 3413 2238
rect 1669 2169 1677 2203
rect 1711 2169 1747 2203
rect 1781 2169 1817 2203
rect 1851 2169 1887 2203
rect 1921 2169 1957 2203
rect 1991 2169 2027 2203
rect 2061 2169 2097 2203
rect 2131 2169 2167 2203
rect 2201 2169 2237 2203
rect 2271 2169 2307 2203
rect 2341 2169 2377 2203
rect 2411 2169 2447 2203
rect 2481 2169 2517 2203
rect 2551 2169 2587 2203
rect 2621 2169 2657 2203
rect 2691 2169 2727 2203
rect 2761 2169 2797 2203
rect 2831 2169 2867 2203
rect 2901 2169 2937 2203
rect 2971 2169 3007 2203
rect 3041 2169 3077 2203
rect 3111 2169 3147 2203
rect 3181 2169 3217 2203
rect 3251 2169 3287 2203
rect 3321 2169 3413 2203
rect 1669 2134 3413 2169
rect 1669 2100 1677 2134
rect 1711 2100 1747 2134
rect 1781 2100 1817 2134
rect 1851 2100 1887 2134
rect 1921 2100 1957 2134
rect 1991 2100 2027 2134
rect 2061 2100 2097 2134
rect 2131 2100 2167 2134
rect 2201 2100 2237 2134
rect 2271 2100 2307 2134
rect 2341 2100 2377 2134
rect 2411 2100 2447 2134
rect 2481 2100 2517 2134
rect 2551 2100 2587 2134
rect 2621 2100 2657 2134
rect 2691 2100 2727 2134
rect 2761 2100 2797 2134
rect 2831 2100 2867 2134
rect 2901 2100 2937 2134
rect 2971 2100 3007 2134
rect 3041 2100 3077 2134
rect 3111 2100 3147 2134
rect 3181 2100 3217 2134
rect 3251 2100 3287 2134
rect 3321 2100 3413 2134
rect 1669 2065 3413 2100
rect 1669 2031 1677 2065
rect 1711 2031 1747 2065
rect 1781 2031 1817 2065
rect 1851 2031 1887 2065
rect 1921 2031 1957 2065
rect 1991 2031 2027 2065
rect 2061 2031 2097 2065
rect 2131 2031 2167 2065
rect 2201 2031 2237 2065
rect 2271 2031 2307 2065
rect 2341 2031 2377 2065
rect 2411 2031 2447 2065
rect 2481 2031 2517 2065
rect 2551 2031 2587 2065
rect 2621 2031 2657 2065
rect 2691 2031 2727 2065
rect 2761 2031 2797 2065
rect 2831 2031 2867 2065
rect 2901 2031 2937 2065
rect 2971 2031 3007 2065
rect 3041 2031 3077 2065
rect 3111 2031 3147 2065
rect 3181 2031 3217 2065
rect 3251 2031 3287 2065
rect 3321 2031 3413 2065
rect 1669 1996 3413 2031
rect 1669 1962 1677 1996
rect 1711 1962 1747 1996
rect 1781 1962 1817 1996
rect 1851 1962 1887 1996
rect 1921 1962 1957 1996
rect 1991 1962 2027 1996
rect 2061 1962 2097 1996
rect 2131 1962 2167 1996
rect 2201 1962 2237 1996
rect 2271 1962 2307 1996
rect 2341 1962 2377 1996
rect 2411 1962 2447 1996
rect 2481 1962 2517 1996
rect 2551 1962 2587 1996
rect 2621 1962 2657 1996
rect 2691 1962 2727 1996
rect 2761 1962 2797 1996
rect 2831 1962 2867 1996
rect 2901 1962 2937 1996
rect 2971 1962 3007 1996
rect 3041 1962 3077 1996
rect 3111 1962 3147 1996
rect 3181 1962 3217 1996
rect 3251 1962 3287 1996
rect 3321 1962 3413 1996
rect 1669 1927 3413 1962
rect 1669 1893 1677 1927
rect 1711 1893 1747 1927
rect 1781 1893 1817 1927
rect 1851 1893 1887 1927
rect 1921 1893 1957 1927
rect 1991 1893 2027 1927
rect 2061 1893 2097 1927
rect 2131 1893 2167 1927
rect 2201 1893 2237 1927
rect 2271 1893 2307 1927
rect 2341 1893 2377 1927
rect 2411 1893 2447 1927
rect 2481 1893 2517 1927
rect 2551 1893 2587 1927
rect 2621 1893 2657 1927
rect 2691 1893 2727 1927
rect 2761 1893 2797 1927
rect 2831 1893 2867 1927
rect 2901 1893 2937 1927
rect 2971 1893 3007 1927
rect 3041 1893 3077 1927
rect 3111 1893 3147 1927
rect 3181 1893 3217 1927
rect 3251 1893 3287 1927
rect 3321 1893 3413 1927
rect 1669 1858 3413 1893
rect 1669 1824 1677 1858
rect 1711 1824 1747 1858
rect 1781 1824 1817 1858
rect 1851 1824 1887 1858
rect 1921 1824 1957 1858
rect 1991 1824 2027 1858
rect 2061 1824 2097 1858
rect 2131 1824 2167 1858
rect 2201 1824 2237 1858
rect 2271 1824 2307 1858
rect 2341 1824 2377 1858
rect 2411 1824 2447 1858
rect 2481 1824 2517 1858
rect 2551 1824 2587 1858
rect 2621 1824 2657 1858
rect 2691 1824 2727 1858
rect 2761 1824 2797 1858
rect 2831 1824 2867 1858
rect 2901 1824 2937 1858
rect 2971 1824 3007 1858
rect 3041 1824 3077 1858
rect 3111 1824 3147 1858
rect 3181 1824 3217 1858
rect 3251 1824 3287 1858
rect 3321 1824 3413 1858
rect 1669 1789 3413 1824
rect 1669 1755 1677 1789
rect 1711 1755 1747 1789
rect 1781 1755 1817 1789
rect 1851 1755 1887 1789
rect 1921 1755 1957 1789
rect 1991 1755 2027 1789
rect 2061 1755 2097 1789
rect 2131 1755 2167 1789
rect 2201 1755 2237 1789
rect 2271 1755 2307 1789
rect 2341 1755 2377 1789
rect 2411 1755 2447 1789
rect 2481 1755 2517 1789
rect 2551 1755 2587 1789
rect 2621 1755 2657 1789
rect 2691 1755 2727 1789
rect 2761 1755 2797 1789
rect 2831 1755 2867 1789
rect 2901 1755 2937 1789
rect 2971 1755 3007 1789
rect 3041 1755 3077 1789
rect 3111 1755 3147 1789
rect 3181 1755 3217 1789
rect 3251 1755 3287 1789
rect 3321 1755 3413 1789
rect 1669 1720 3413 1755
rect 1669 1686 1677 1720
rect 1711 1686 1747 1720
rect 1781 1686 1817 1720
rect 1851 1686 1887 1720
rect 1921 1686 1957 1720
rect 1991 1686 2027 1720
rect 2061 1686 2097 1720
rect 2131 1686 2167 1720
rect 2201 1686 2237 1720
rect 2271 1686 2307 1720
rect 2341 1686 2377 1720
rect 2411 1686 2447 1720
rect 2481 1686 2517 1720
rect 2551 1686 2587 1720
rect 2621 1686 2657 1720
rect 2691 1686 2727 1720
rect 2761 1686 2797 1720
rect 2831 1686 2867 1720
rect 2901 1686 2937 1720
rect 2971 1686 3007 1720
rect 3041 1686 3077 1720
rect 3111 1686 3147 1720
rect 3181 1686 3217 1720
rect 3251 1686 3287 1720
rect 3321 1686 3413 1720
rect 1669 1651 3413 1686
rect 1669 1617 1677 1651
rect 1711 1617 1747 1651
rect 1781 1617 1817 1651
rect 1851 1617 1887 1651
rect 1921 1617 1957 1651
rect 1991 1617 2027 1651
rect 2061 1617 2097 1651
rect 2131 1617 2167 1651
rect 2201 1617 2237 1651
rect 2271 1617 2307 1651
rect 2341 1617 2377 1651
rect 2411 1617 2447 1651
rect 2481 1617 2517 1651
rect 2551 1617 2587 1651
rect 2621 1617 2657 1651
rect 2691 1617 2727 1651
rect 2761 1617 2797 1651
rect 2831 1617 2867 1651
rect 2901 1617 2937 1651
rect 2971 1617 3007 1651
rect 3041 1617 3077 1651
rect 3111 1617 3147 1651
rect 3181 1617 3217 1651
rect 3251 1617 3287 1651
rect 3321 1617 3413 1651
rect 1669 1582 3413 1617
rect 1669 1548 1677 1582
rect 1711 1548 1747 1582
rect 1781 1548 1817 1582
rect 1851 1548 1887 1582
rect 1921 1548 1957 1582
rect 1991 1548 2027 1582
rect 2061 1548 2097 1582
rect 2131 1548 2167 1582
rect 2201 1548 2237 1582
rect 2271 1548 2307 1582
rect 2341 1548 2377 1582
rect 2411 1548 2447 1582
rect 2481 1548 2517 1582
rect 2551 1548 2587 1582
rect 2621 1548 2657 1582
rect 2691 1548 2727 1582
rect 2761 1548 2797 1582
rect 2831 1548 2867 1582
rect 2901 1548 2937 1582
rect 2971 1548 3007 1582
rect 3041 1548 3077 1582
rect 3111 1548 3147 1582
rect 3181 1548 3217 1582
rect 3251 1548 3287 1582
rect 3321 1548 3413 1582
rect 1669 1513 3413 1548
rect 1669 1479 1677 1513
rect 1711 1479 1747 1513
rect 1781 1479 1817 1513
rect 1851 1479 1887 1513
rect 1921 1479 1957 1513
rect 1991 1479 2027 1513
rect 2061 1479 2097 1513
rect 2131 1479 2167 1513
rect 2201 1479 2237 1513
rect 2271 1479 2307 1513
rect 2341 1479 2377 1513
rect 2411 1479 2447 1513
rect 2481 1479 2517 1513
rect 2551 1479 2587 1513
rect 2621 1479 2657 1513
rect 2691 1479 2727 1513
rect 2761 1479 2797 1513
rect 2831 1479 2867 1513
rect 2901 1479 2937 1513
rect 2971 1479 3007 1513
rect 3041 1479 3077 1513
rect 3111 1479 3147 1513
rect 3181 1479 3217 1513
rect 3251 1479 3287 1513
rect 3321 1479 3413 1513
rect 1669 1444 3413 1479
rect 1669 1410 1677 1444
rect 1711 1410 1747 1444
rect 1781 1410 1817 1444
rect 1851 1410 1887 1444
rect 1921 1410 1957 1444
rect 1991 1410 2027 1444
rect 2061 1410 2097 1444
rect 2131 1410 2167 1444
rect 2201 1410 2237 1444
rect 2271 1410 2307 1444
rect 2341 1410 2377 1444
rect 2411 1410 2447 1444
rect 2481 1410 2517 1444
rect 2551 1410 2587 1444
rect 2621 1410 2657 1444
rect 2691 1410 2727 1444
rect 2761 1410 2797 1444
rect 2831 1410 2867 1444
rect 2901 1410 2937 1444
rect 2971 1410 3007 1444
rect 3041 1410 3077 1444
rect 3111 1410 3147 1444
rect 3181 1410 3217 1444
rect 3251 1410 3287 1444
rect 3321 1410 3413 1444
rect 1669 1375 3413 1410
rect 1669 1341 1677 1375
rect 1711 1341 1747 1375
rect 1781 1341 1817 1375
rect 1851 1341 1887 1375
rect 1921 1341 1957 1375
rect 1991 1341 2027 1375
rect 2061 1341 2097 1375
rect 2131 1341 2167 1375
rect 2201 1341 2237 1375
rect 2271 1341 2307 1375
rect 2341 1341 2377 1375
rect 2411 1341 2447 1375
rect 2481 1341 2517 1375
rect 2551 1341 2587 1375
rect 2621 1341 2657 1375
rect 2691 1341 2727 1375
rect 2761 1341 2797 1375
rect 2831 1341 2867 1375
rect 2901 1341 2937 1375
rect 2971 1341 3007 1375
rect 3041 1341 3077 1375
rect 3111 1341 3147 1375
rect 3181 1341 3217 1375
rect 3251 1341 3287 1375
rect 3321 1341 3413 1375
rect 1669 1306 3413 1341
rect 1669 1272 1677 1306
rect 1711 1272 1747 1306
rect 1781 1272 1817 1306
rect 1851 1272 1887 1306
rect 1921 1272 1957 1306
rect 1991 1272 2027 1306
rect 2061 1272 2097 1306
rect 2131 1272 2167 1306
rect 2201 1272 2237 1306
rect 2271 1272 2307 1306
rect 2341 1272 2377 1306
rect 2411 1272 2447 1306
rect 2481 1272 2517 1306
rect 2551 1272 2587 1306
rect 2621 1272 2657 1306
rect 2691 1272 2727 1306
rect 2761 1272 2797 1306
rect 2831 1272 2867 1306
rect 2901 1272 2937 1306
rect 2971 1272 3007 1306
rect 3041 1272 3077 1306
rect 3111 1272 3147 1306
rect 3181 1272 3217 1306
rect 3251 1272 3287 1306
rect 3321 1272 3413 1306
rect 1669 1237 3413 1272
rect 1669 1203 1677 1237
rect 1711 1203 1747 1237
rect 1781 1203 1817 1237
rect 1851 1203 1887 1237
rect 1921 1203 1957 1237
rect 1991 1203 2027 1237
rect 2061 1203 2097 1237
rect 2131 1203 2167 1237
rect 2201 1203 2237 1237
rect 2271 1203 2307 1237
rect 2341 1203 2377 1237
rect 2411 1203 2447 1237
rect 2481 1203 2517 1237
rect 2551 1203 2587 1237
rect 2621 1203 2657 1237
rect 2691 1203 2727 1237
rect 2761 1203 2797 1237
rect 2831 1203 2867 1237
rect 2901 1203 2937 1237
rect 2971 1203 3007 1237
rect 3041 1203 3077 1237
rect 3111 1203 3147 1237
rect 3181 1203 3217 1237
rect 3251 1203 3287 1237
rect 3321 1203 3413 1237
rect 1669 1168 3413 1203
rect 1669 1134 1677 1168
rect 1711 1134 1747 1168
rect 1781 1134 1817 1168
rect 1851 1134 1887 1168
rect 1921 1134 1957 1168
rect 1991 1134 2027 1168
rect 2061 1134 2097 1168
rect 2131 1134 2167 1168
rect 2201 1134 2237 1168
rect 2271 1134 2307 1168
rect 2341 1134 2377 1168
rect 2411 1134 2447 1168
rect 2481 1134 2517 1168
rect 2551 1134 2587 1168
rect 2621 1134 2657 1168
rect 2691 1134 2727 1168
rect 2761 1134 2797 1168
rect 2831 1134 2867 1168
rect 2901 1134 2937 1168
rect 2971 1134 3007 1168
rect 3041 1134 3077 1168
rect 3111 1134 3147 1168
rect 3181 1134 3217 1168
rect 3251 1134 3287 1168
rect 3321 1134 3413 1168
rect 1669 1099 3413 1134
rect 1669 1065 1677 1099
rect 1711 1065 1747 1099
rect 1781 1065 1817 1099
rect 1851 1065 1887 1099
rect 1921 1065 1957 1099
rect 1991 1065 2027 1099
rect 2061 1065 2097 1099
rect 2131 1065 2167 1099
rect 2201 1065 2237 1099
rect 2271 1065 2307 1099
rect 2341 1065 2377 1099
rect 2411 1065 2447 1099
rect 2481 1065 2517 1099
rect 2551 1065 2587 1099
rect 2621 1065 2657 1099
rect 2691 1065 2727 1099
rect 2761 1065 2797 1099
rect 2831 1065 2867 1099
rect 2901 1065 2937 1099
rect 2971 1065 3007 1099
rect 3041 1065 3077 1099
rect 3111 1065 3147 1099
rect 3181 1065 3217 1099
rect 3251 1065 3287 1099
rect 3321 1065 3413 1099
rect 1669 1030 3413 1065
rect 1669 996 1677 1030
rect 1711 996 1747 1030
rect 1781 996 1817 1030
rect 1851 996 1887 1030
rect 1921 996 1957 1030
rect 1991 996 2027 1030
rect 2061 996 2097 1030
rect 2131 996 2167 1030
rect 2201 996 2237 1030
rect 2271 996 2307 1030
rect 2341 996 2377 1030
rect 2411 996 2447 1030
rect 2481 996 2517 1030
rect 2551 996 2587 1030
rect 2621 996 2657 1030
rect 2691 996 2727 1030
rect 2761 996 2797 1030
rect 2831 996 2867 1030
rect 2901 996 2937 1030
rect 2971 996 3007 1030
rect 3041 996 3077 1030
rect 3111 996 3147 1030
rect 3181 996 3217 1030
rect 3251 996 3287 1030
rect 3321 996 3413 1030
rect 1669 961 3413 996
rect 1669 927 1677 961
rect 1711 927 1747 961
rect 1781 927 1817 961
rect 1851 927 1887 961
rect 1921 927 1957 961
rect 1991 927 2027 961
rect 2061 927 2097 961
rect 2131 927 2167 961
rect 2201 927 2237 961
rect 2271 927 2307 961
rect 2341 927 2377 961
rect 2411 927 2447 961
rect 2481 927 2517 961
rect 2551 927 2587 961
rect 2621 927 2657 961
rect 2691 927 2727 961
rect 2761 927 2797 961
rect 2831 927 2867 961
rect 2901 927 2937 961
rect 2971 927 3007 961
rect 3041 927 3077 961
rect 3111 927 3147 961
rect 3181 927 3217 961
rect 3251 927 3287 961
rect 3321 927 3413 961
rect 1669 892 3413 927
rect 1669 858 1677 892
rect 1711 858 1747 892
rect 1781 858 1817 892
rect 1851 858 1887 892
rect 1921 858 1957 892
rect 1991 858 2027 892
rect 2061 858 2097 892
rect 2131 858 2167 892
rect 2201 858 2237 892
rect 2271 858 2307 892
rect 2341 858 2377 892
rect 2411 858 2447 892
rect 2481 858 2517 892
rect 2551 858 2587 892
rect 2621 858 2657 892
rect 2691 858 2727 892
rect 2761 858 2797 892
rect 2831 858 2867 892
rect 2901 858 2937 892
rect 2971 858 3007 892
rect 3041 858 3077 892
rect 3111 858 3147 892
rect 3181 858 3217 892
rect 3251 858 3287 892
rect 3321 858 3413 892
rect 1669 823 3413 858
rect 1669 789 1677 823
rect 1711 789 1747 823
rect 1781 789 1817 823
rect 1851 789 1887 823
rect 1921 789 1957 823
rect 1991 789 2027 823
rect 2061 789 2097 823
rect 2131 789 2167 823
rect 2201 789 2237 823
rect 2271 789 2307 823
rect 2341 789 2377 823
rect 2411 789 2447 823
rect 2481 789 2517 823
rect 2551 789 2587 823
rect 2621 789 2657 823
rect 2691 789 2727 823
rect 2761 789 2797 823
rect 2831 789 2867 823
rect 2901 789 2937 823
rect 2971 789 3007 823
rect 3041 789 3077 823
rect 3111 789 3147 823
rect 3181 789 3217 823
rect 3251 789 3287 823
rect 3321 789 3413 823
rect 1669 754 3413 789
rect 1669 720 1677 754
rect 1711 720 1747 754
rect 1781 720 1817 754
rect 1851 720 1887 754
rect 1921 720 1957 754
rect 1991 720 2027 754
rect 2061 720 2097 754
rect 2131 720 2167 754
rect 2201 720 2237 754
rect 2271 720 2307 754
rect 2341 720 2377 754
rect 2411 720 2447 754
rect 2481 720 2517 754
rect 2551 720 2587 754
rect 2621 720 2657 754
rect 2691 720 2727 754
rect 2761 720 2797 754
rect 2831 720 2867 754
rect 2901 720 2937 754
rect 2971 720 3007 754
rect 3041 720 3077 754
rect 3111 720 3147 754
rect 3181 720 3217 754
rect 3251 720 3287 754
rect 3321 720 3413 754
rect 1669 685 3413 720
rect 1669 651 1677 685
rect 1711 651 1747 685
rect 1781 651 1817 685
rect 1851 651 1887 685
rect 1921 651 1957 685
rect 1991 651 2027 685
rect 2061 651 2097 685
rect 2131 651 2167 685
rect 2201 651 2237 685
rect 2271 651 2307 685
rect 2341 651 2377 685
rect 2411 651 2447 685
rect 2481 651 2517 685
rect 2551 651 2587 685
rect 2621 651 2657 685
rect 2691 651 2727 685
rect 2761 651 2797 685
rect 2831 651 2867 685
rect 2901 651 2937 685
rect 2971 651 3007 685
rect 3041 651 3077 685
rect 3111 651 3147 685
rect 3181 651 3217 685
rect 3251 651 3287 685
rect 3321 651 3413 685
rect 1669 616 3413 651
rect 1669 582 1677 616
rect 1711 582 1747 616
rect 1781 582 1817 616
rect 1851 582 1887 616
rect 1921 582 1957 616
rect 1991 582 2027 616
rect 2061 582 2097 616
rect 2131 582 2167 616
rect 2201 582 2237 616
rect 2271 582 2307 616
rect 2341 582 2377 616
rect 2411 582 2447 616
rect 2481 582 2517 616
rect 2551 582 2587 616
rect 2621 582 2657 616
rect 2691 582 2727 616
rect 2761 582 2797 616
rect 2831 582 2867 616
rect 2901 582 2937 616
rect 2971 582 3007 616
rect 3041 582 3077 616
rect 3111 582 3147 616
rect 3181 582 3217 616
rect 3251 582 3287 616
rect 3321 582 3413 616
rect 1669 547 3413 582
rect 1669 513 1677 547
rect 1711 513 1747 547
rect 1781 513 1817 547
rect 1851 513 1887 547
rect 1921 513 1957 547
rect 1991 513 2027 547
rect 2061 513 2097 547
rect 2131 513 2167 547
rect 2201 513 2237 547
rect 2271 513 2307 547
rect 2341 513 2377 547
rect 2411 513 2447 547
rect 2481 513 2517 547
rect 2551 513 2587 547
rect 2621 513 2657 547
rect 2691 513 2727 547
rect 2761 513 2797 547
rect 2831 513 2867 547
rect 2901 513 2937 547
rect 2971 513 3007 547
rect 3041 513 3077 547
rect 3111 513 3147 547
rect 3181 513 3217 547
rect 3251 513 3287 547
rect 3321 513 3413 547
rect 1669 478 3413 513
rect 1669 444 1677 478
rect 1711 444 1747 478
rect 1781 444 1817 478
rect 1851 444 1887 478
rect 1921 444 1957 478
rect 1991 444 2027 478
rect 2061 444 2097 478
rect 2131 444 2167 478
rect 2201 444 2237 478
rect 2271 444 2307 478
rect 2341 444 2377 478
rect 2411 444 2447 478
rect 2481 444 2517 478
rect 2551 444 2587 478
rect 2621 444 2657 478
rect 2691 444 2727 478
rect 2761 444 2797 478
rect 2831 444 2867 478
rect 2901 444 2937 478
rect 2971 444 3007 478
rect 3041 444 3077 478
rect 3111 444 3147 478
rect 3181 444 3217 478
rect 3251 444 3287 478
rect 3321 444 3413 478
rect 1669 409 3413 444
rect 1669 375 1677 409
rect 1711 375 1747 409
rect 1781 375 1817 409
rect 1851 375 1887 409
rect 1921 375 1957 409
rect 1991 375 2027 409
rect 2061 375 2097 409
rect 2131 375 2167 409
rect 2201 375 2237 409
rect 2271 375 2307 409
rect 2341 375 2377 409
rect 2411 375 2447 409
rect 2481 375 2517 409
rect 2551 375 2587 409
rect 2621 375 2657 409
rect 2691 375 2727 409
rect 2761 375 2797 409
rect 2831 375 2867 409
rect 2901 375 2937 409
rect 2971 375 3007 409
rect 3041 375 3077 409
rect 3111 375 3147 409
rect 3181 375 3217 409
rect 3251 375 3287 409
rect 3321 375 3413 409
rect 1669 340 3413 375
rect 1669 306 1677 340
rect 1711 306 1747 340
rect 1781 306 1817 340
rect 1851 306 1887 340
rect 1921 306 1957 340
rect 1991 306 2027 340
rect 2061 306 2097 340
rect 2131 306 2167 340
rect 2201 306 2237 340
rect 2271 306 2307 340
rect 2341 306 2377 340
rect 2411 306 2447 340
rect 2481 306 2517 340
rect 2551 306 2587 340
rect 2621 306 2657 340
rect 2691 306 2727 340
rect 2761 306 2797 340
rect 2831 306 2867 340
rect 2901 306 2937 340
rect 2971 306 3007 340
rect 3041 306 3077 340
rect 3111 306 3147 340
rect 3181 306 3217 340
rect 3251 306 3287 340
rect 3321 306 3413 340
rect 1669 282 3413 306
<< nsubdiff >>
rect 270 3408 368 3442
rect 402 3408 436 3442
rect 470 3408 504 3442
rect 538 3408 572 3442
rect 606 3408 640 3442
rect 674 3408 708 3442
rect 742 3408 776 3442
rect 810 3408 844 3442
rect 878 3408 912 3442
rect 946 3408 980 3442
rect 1014 3408 1048 3442
rect 1082 3408 1116 3442
rect 1150 3408 1184 3442
rect 1218 3408 1252 3442
rect 1286 3408 1320 3442
rect 1354 3408 1422 3442
rect 270 3374 304 3408
rect 270 3306 304 3340
rect 270 3238 304 3272
rect 270 3170 304 3204
rect 270 3102 304 3136
rect 270 3034 304 3068
rect 270 2966 304 3000
rect 270 2898 304 2932
rect 270 2830 304 2864
rect 270 2762 304 2796
rect 270 2694 304 2728
rect 270 2626 304 2660
rect 270 2558 304 2592
rect 270 2490 304 2524
rect 270 2422 304 2456
rect 270 2354 304 2388
rect 270 2286 304 2320
rect 270 2218 304 2252
rect 270 2150 304 2184
rect 270 2082 304 2116
rect 270 2014 304 2048
rect 270 1946 304 1980
rect 270 1878 304 1912
rect 1388 3366 1422 3408
rect 1388 3298 1422 3332
rect 1388 3230 1422 3264
rect 1388 3162 1422 3196
rect 1388 3094 1422 3128
rect 1388 3026 1422 3060
rect 1388 2958 1422 2992
rect 1388 2890 1422 2924
rect 1388 2822 1422 2856
rect 1388 2754 1422 2788
rect 1388 2686 1422 2720
rect 1388 2618 1422 2652
rect 1388 2550 1422 2584
rect 1388 2482 1422 2516
rect 1388 2414 1422 2448
rect 1388 2346 1422 2380
rect 1388 2278 1422 2312
rect 1388 2210 1422 2244
rect 1388 2142 1422 2176
rect 1388 2074 1422 2108
rect 1388 2006 1422 2040
rect 1388 1938 1422 1972
rect 270 1810 304 1844
rect 1388 1870 1422 1904
rect 270 1742 304 1776
rect 270 1674 304 1708
rect 270 1606 304 1640
rect 270 1538 304 1572
rect 270 1470 304 1504
rect 270 1402 304 1436
rect 270 1334 304 1368
rect 270 1266 304 1300
rect 270 1198 304 1232
rect 270 1130 304 1164
rect 270 1062 304 1096
rect 270 994 304 1028
rect 270 926 304 960
rect 270 858 304 892
rect 270 790 304 824
rect 270 722 304 756
rect 270 654 304 688
rect 270 586 304 620
rect 270 518 304 552
rect 270 450 304 484
rect 270 382 304 416
rect 1388 1802 1422 1836
rect 1388 1734 1422 1768
rect 1388 1666 1422 1700
rect 1388 1598 1422 1632
rect 1388 1530 1422 1564
rect 1388 1462 1422 1496
rect 1388 1394 1422 1428
rect 1388 1326 1422 1360
rect 1388 1258 1422 1292
rect 1388 1190 1422 1224
rect 1388 1122 1422 1156
rect 1388 1054 1422 1088
rect 1388 986 1422 1020
rect 1388 918 1422 952
rect 1388 850 1422 884
rect 1388 782 1422 816
rect 1388 714 1422 748
rect 1388 646 1422 680
rect 1388 578 1422 612
rect 1388 510 1422 544
rect 1388 442 1422 476
rect 1388 374 1422 408
rect 270 238 304 348
rect 1388 306 1422 340
rect 13523 3420 13621 3454
rect 13655 3420 13689 3454
rect 13723 3420 13757 3454
rect 13791 3420 13825 3454
rect 13859 3420 13893 3454
rect 13927 3420 13961 3454
rect 13995 3420 14029 3454
rect 14063 3420 14097 3454
rect 14131 3420 14165 3454
rect 14199 3420 14233 3454
rect 14267 3420 14301 3454
rect 14335 3420 14369 3454
rect 14403 3420 14437 3454
rect 14471 3420 14505 3454
rect 14539 3420 14573 3454
rect 14607 3420 14675 3454
rect 13523 3386 13557 3420
rect 13523 3318 13557 3352
rect 13523 3250 13557 3284
rect 13523 3182 13557 3216
rect 13523 3114 13557 3148
rect 13523 3046 13557 3080
rect 13523 2978 13557 3012
rect 13523 2910 13557 2944
rect 13523 2842 13557 2876
rect 13523 2774 13557 2808
rect 13523 2706 13557 2740
rect 13523 2638 13557 2672
rect 13523 2570 13557 2604
rect 13523 2502 13557 2536
rect 13523 2434 13557 2468
rect 13523 2366 13557 2400
rect 13523 2298 13557 2332
rect 13523 2230 13557 2264
rect 13523 2162 13557 2196
rect 13523 2094 13557 2128
rect 13523 2026 13557 2060
rect 13523 1958 13557 1992
rect 13523 1890 13557 1924
rect 14641 3378 14675 3420
rect 14641 3310 14675 3344
rect 14641 3242 14675 3276
rect 14641 3174 14675 3208
rect 14641 3106 14675 3140
rect 14641 3038 14675 3072
rect 14641 2970 14675 3004
rect 14641 2902 14675 2936
rect 14641 2834 14675 2868
rect 14641 2766 14675 2800
rect 14641 2698 14675 2732
rect 14641 2630 14675 2664
rect 14641 2562 14675 2596
rect 14641 2494 14675 2528
rect 14641 2426 14675 2460
rect 14641 2358 14675 2392
rect 14641 2290 14675 2324
rect 14641 2222 14675 2256
rect 14641 2154 14675 2188
rect 14641 2086 14675 2120
rect 14641 2018 14675 2052
rect 14641 1950 14675 1984
rect 13523 1822 13557 1856
rect 14641 1882 14675 1916
rect 13523 1754 13557 1788
rect 13523 1686 13557 1720
rect 13523 1618 13557 1652
rect 13523 1550 13557 1584
rect 13523 1482 13557 1516
rect 13523 1414 13557 1448
rect 13523 1346 13557 1380
rect 13523 1278 13557 1312
rect 13523 1210 13557 1244
rect 13523 1142 13557 1176
rect 13523 1074 13557 1108
rect 13523 1006 13557 1040
rect 13523 938 13557 972
rect 13523 870 13557 904
rect 13523 802 13557 836
rect 13523 734 13557 768
rect 13523 666 13557 700
rect 13523 598 13557 632
rect 13523 530 13557 564
rect 13523 462 13557 496
rect 13523 394 13557 428
rect 14641 1814 14675 1848
rect 14641 1746 14675 1780
rect 14641 1678 14675 1712
rect 14641 1610 14675 1644
rect 14641 1542 14675 1576
rect 14641 1474 14675 1508
rect 14641 1406 14675 1440
rect 14641 1338 14675 1372
rect 14641 1270 14675 1304
rect 14641 1202 14675 1236
rect 14641 1134 14675 1168
rect 14641 1066 14675 1100
rect 14641 998 14675 1032
rect 14641 930 14675 964
rect 14641 862 14675 896
rect 14641 794 14675 828
rect 14641 726 14675 760
rect 14641 658 14675 692
rect 14641 590 14675 624
rect 14641 522 14675 556
rect 14641 454 14675 488
rect 14641 386 14675 420
rect 1388 238 1422 272
rect 270 204 338 238
rect 372 204 406 238
rect 440 204 474 238
rect 508 204 542 238
rect 576 204 610 238
rect 644 204 678 238
rect 712 204 746 238
rect 780 204 814 238
rect 848 204 882 238
rect 916 204 950 238
rect 984 204 1018 238
rect 1052 204 1086 238
rect 1120 204 1154 238
rect 1188 204 1222 238
rect 1256 204 1290 238
rect 1324 204 1422 238
rect 13523 250 13557 360
rect 14641 318 14675 352
rect 14641 250 14675 284
rect 13523 216 13591 250
rect 13625 216 13659 250
rect 13693 216 13727 250
rect 13761 216 13795 250
rect 13829 216 13863 250
rect 13897 216 13931 250
rect 13965 216 13999 250
rect 14033 216 14067 250
rect 14101 216 14135 250
rect 14169 216 14203 250
rect 14237 216 14271 250
rect 14305 216 14339 250
rect 14373 216 14407 250
rect 14441 216 14475 250
rect 14509 216 14543 250
rect 14577 216 14675 250
<< mvnsubdiff >>
rect 1946 39440 2076 39474
rect 2110 39440 2144 39474
rect 1946 39406 2144 39440
rect 2048 39372 2144 39406
rect 13874 39372 13942 39474
rect 13840 39355 13942 39372
rect 13840 39321 13908 39355
rect 13840 39287 13942 39321
rect 4314 19985 4382 20019
rect 4416 19985 4450 20019
rect 4484 19985 4518 20019
rect 4552 19985 4586 20019
rect 4620 19985 4654 20019
rect 4688 19985 4722 20019
rect 4756 19985 4790 20019
rect 4824 19985 4858 20019
rect 4892 19985 4926 20019
rect 4960 19985 4994 20019
rect 5028 19985 5062 20019
rect 5096 19985 5130 20019
rect 5164 19985 5198 20019
rect 5232 19985 5266 20019
rect 5300 19985 5334 20019
rect 5368 19985 5402 20019
rect 5436 19985 5470 20019
rect 5504 19985 5538 20019
rect 5572 19985 5606 20019
rect 5640 19985 5674 20019
rect 5708 19985 5742 20019
rect 5776 19985 5810 20019
rect 5844 19985 5878 20019
rect 5912 19985 5946 20019
rect 5980 19985 6014 20019
rect 6048 19985 6082 20019
rect 6116 19985 6150 20019
rect 6184 19985 6218 20019
rect 6252 19985 6286 20019
rect 6320 19985 6354 20019
rect 6388 19985 6422 20019
rect 6456 19985 6490 20019
rect 6524 19985 6558 20019
rect 6592 19985 6626 20019
rect 6660 19985 6694 20019
rect 6728 19985 6762 20019
rect 6796 19985 6830 20019
rect 6864 19985 6898 20019
rect 6932 19985 6966 20019
rect 7000 19985 7034 20019
rect 7068 19985 7102 20019
rect 7136 19985 7170 20019
rect 7204 19985 7238 20019
rect 7272 19985 7306 20019
rect 7340 19985 7374 20019
rect 7408 19985 7442 20019
rect 7476 19985 7510 20019
rect 7544 19985 7578 20019
rect 7612 19985 7646 20019
rect 7680 19985 7714 20019
rect 7748 19985 7782 20019
rect 7816 19985 7850 20019
rect 7884 19985 7918 20019
rect 7952 19985 7986 20019
rect 8020 19985 8054 20019
rect 8088 19985 8122 20019
rect 8156 19985 8190 20019
rect 8224 19985 8258 20019
rect 8292 19985 8326 20019
rect 8360 19985 8394 20019
rect 8428 19985 8462 20019
rect 8496 19985 8530 20019
rect 8564 19985 8598 20019
rect 8632 19985 8666 20019
rect 8700 19985 8734 20019
rect 8768 19985 8802 20019
rect 8836 19985 8870 20019
rect 8904 19985 8938 20019
rect 8972 19985 9006 20019
rect 9040 19985 9074 20019
rect 9108 19985 9142 20019
rect 9176 19985 9210 20019
rect 9244 19985 9278 20019
rect 9312 19985 9346 20019
rect 9380 19985 9414 20019
rect 9448 19985 9482 20019
rect 9516 19985 9550 20019
rect 9584 19985 9618 20019
rect 9652 19985 9686 20019
rect 9720 19985 9754 20019
rect 9788 19985 9822 20019
rect 9856 19985 9890 20019
rect 9924 19985 9958 20019
rect 9992 19985 10026 20019
rect 10060 19985 10094 20019
rect 10128 19985 10162 20019
rect 10196 19985 10230 20019
rect 10264 19985 10298 20019
rect 10332 19985 10366 20019
rect 10400 19985 10434 20019
rect 10468 19985 10502 20019
rect 10536 19985 10570 20019
rect 10604 19985 10638 20019
rect 10672 19985 10706 20019
rect 10740 19985 10774 20019
rect 10808 19985 10842 20019
rect 10876 19985 10910 20019
rect 10944 19985 10978 20019
rect 11012 19985 11046 20019
rect 11080 19985 11114 20019
rect 11148 19985 11182 20019
rect 11216 19985 11250 20019
rect 11284 19985 11318 20019
rect 11352 19985 11386 20019
rect 11420 19985 11454 20019
rect 11488 19985 11522 20019
rect 11556 19985 11590 20019
rect 11624 19985 11658 20019
rect 11692 19985 11726 20019
rect 11760 19985 11794 20019
rect 11828 19985 11862 20019
rect 11896 19985 11930 20019
rect 11964 19985 11998 20019
rect 12032 19985 12066 20019
rect 12100 19985 12134 20019
rect 12168 19985 12202 20019
rect 12236 19985 12270 20019
rect 12304 19985 12338 20019
rect 12372 19985 12406 20019
rect 12440 19985 12474 20019
rect 12508 19985 12542 20019
rect 12576 19985 12610 20019
rect 12644 19985 12678 20019
rect 12712 19985 12746 20019
rect 12780 19985 12814 20019
rect 12848 19985 12882 20019
rect 12916 19985 12950 20019
rect 12984 19985 13018 20019
rect 13052 19985 13086 20019
rect 13120 19985 13154 20019
rect 13188 19985 13222 20019
rect 13256 19985 13290 20019
rect 13324 19985 13358 20019
rect 13392 19985 13426 20019
rect 13460 19985 13494 20019
rect 13528 19985 13562 20019
rect 13596 19985 13630 20019
rect 13664 19985 13840 20019
rect 4314 19894 4348 19985
rect 4314 19826 4348 19860
rect 4314 19758 4348 19792
rect 4314 19690 4348 19724
rect 4314 19622 4348 19656
rect 4314 19554 4348 19588
rect 4314 19486 4348 19520
rect 4314 19418 4348 19452
rect 4314 19350 4348 19384
rect 4314 19282 4348 19316
rect 4314 19214 4348 19248
rect 4314 19146 4348 19180
rect 4314 19078 4348 19112
rect 4314 19010 4348 19044
rect 4314 18942 4348 18976
rect 4314 18874 4348 18908
rect 4314 18806 4348 18840
rect 4314 18738 4348 18772
rect 4314 18670 4348 18704
rect 4314 18602 4348 18636
rect 4314 18534 4348 18568
rect 4314 18466 4348 18500
rect 4314 18398 4348 18432
rect 4314 18330 4348 18364
rect 4314 18262 4348 18296
rect 4314 18194 4348 18228
rect 4314 18126 4348 18160
rect 4314 18058 4348 18092
rect 4314 17990 4348 18024
rect 4314 17922 4348 17956
rect 4314 17854 4348 17888
rect 4314 17786 4348 17820
rect 4314 17718 4348 17752
rect 4314 17650 4348 17684
rect 4314 17582 4348 17616
rect 4314 17514 4348 17548
rect 4314 17446 4348 17480
rect 4314 17378 4348 17412
rect 4314 17310 4348 17344
rect 4314 17242 4348 17276
rect 4314 17174 4348 17208
rect 4314 17106 4348 17140
rect 4314 17038 4348 17072
rect 4314 16970 4348 17004
rect 4314 16902 4348 16936
rect 4314 16834 4348 16868
rect 4314 16766 4348 16800
rect 4314 16698 4348 16732
rect 4314 16630 4348 16664
rect 2048 16596 2208 16630
rect 2242 16596 2276 16630
rect 2310 16596 2344 16630
rect 2378 16596 2412 16630
rect 2446 16596 2480 16630
rect 2514 16596 2548 16630
rect 2582 16596 2616 16630
rect 2650 16596 2684 16630
rect 2718 16596 2752 16630
rect 2786 16596 2820 16630
rect 2854 16596 2888 16630
rect 2922 16596 2956 16630
rect 2990 16596 3024 16630
rect 3058 16596 3092 16630
rect 3126 16596 3160 16630
rect 3194 16596 3228 16630
rect 3262 16596 3296 16630
rect 3330 16596 3364 16630
rect 3398 16596 3432 16630
rect 3466 16596 3500 16630
rect 3534 16596 3568 16630
rect 3602 16596 3636 16630
rect 3670 16596 3704 16630
rect 3738 16596 3772 16630
rect 3806 16596 3840 16630
rect 3874 16596 3908 16630
rect 3942 16596 3976 16630
rect 4010 16596 4044 16630
rect 4078 16596 4112 16630
rect 4146 16596 4180 16630
rect 4214 16596 4348 16630
rect 1946 5345 2048 5508
rect 13840 5481 13942 5593
rect 2048 4835 2088 4869
rect 1946 4801 2088 4835
rect 1946 4767 2020 4801
rect 2054 4767 2088 4801
rect 2598 4767 2666 4869
rect 13240 4767 13340 4869
rect 13782 4835 13840 4869
rect 13782 4801 13942 4835
rect 13782 4767 13816 4801
rect 13850 4767 13942 4801
<< psubdiffcont >>
rect 2482 39119 2516 39153
rect 2550 39119 2584 39153
rect 2618 39119 2652 39153
rect 2686 39119 2720 39153
rect 2754 39119 2788 39153
rect 2822 39119 2856 39153
rect 2890 39119 2924 39153
rect 2958 39119 2992 39153
rect 3026 39119 3060 39153
rect 3094 39119 3128 39153
rect 3162 39119 3196 39153
rect 3230 39119 3264 39153
rect 3298 39119 3332 39153
rect 3366 39119 3400 39153
rect 3434 39119 3468 39153
rect 3502 39119 3536 39153
rect 3570 39119 3604 39153
rect 3638 39119 3672 39153
rect 3706 39119 3740 39153
rect 3774 39119 3808 39153
rect 3842 39119 3876 39153
rect 3910 39119 3944 39153
rect 3978 39119 4012 39153
rect 4046 39119 4080 39153
rect 4114 39119 4148 39153
rect 4182 39119 4216 39153
rect 4250 39119 4284 39153
rect 4318 39119 4352 39153
rect 4386 39119 4420 39153
rect 4454 39119 4488 39153
rect 4522 39119 4556 39153
rect 4590 39119 4624 39153
rect 4658 39119 4692 39153
rect 4726 39119 4760 39153
rect 4794 39119 4828 39153
rect 4862 39119 4896 39153
rect 4930 39119 4964 39153
rect 4998 39119 5032 39153
rect 5066 39119 5100 39153
rect 5134 39119 5168 39153
rect 5202 39119 5236 39153
rect 5270 39119 5304 39153
rect 5338 39119 5372 39153
rect 5406 39119 5440 39153
rect 5474 39119 5508 39153
rect 5542 39119 5576 39153
rect 5610 39119 5644 39153
rect 5678 39119 5712 39153
rect 5746 39119 5780 39153
rect 5814 39119 5848 39153
rect 5882 39119 5916 39153
rect 5950 39119 5984 39153
rect 6018 39119 6052 39153
rect 6086 39119 6120 39153
rect 6154 39119 6188 39153
rect 6222 39119 6256 39153
rect 6290 39119 6324 39153
rect 6358 39119 6392 39153
rect 6426 39119 6460 39153
rect 6494 39119 6528 39153
rect 6562 39119 6596 39153
rect 6630 39119 6664 39153
rect 6698 39119 6732 39153
rect 6766 39119 6800 39153
rect 6834 39119 6868 39153
rect 6902 39119 6936 39153
rect 6970 39119 7004 39153
rect 7038 39119 7072 39153
rect 7106 39119 7140 39153
rect 7174 39119 7208 39153
rect 7242 39119 7276 39153
rect 7310 39119 7344 39153
rect 7378 39119 7412 39153
rect 7446 39119 7480 39153
rect 7514 39119 7548 39153
rect 7582 39119 7616 39153
rect 7650 39119 7684 39153
rect 7718 39119 7752 39153
rect 7786 39119 7820 39153
rect 7854 39119 7888 39153
rect 7922 39119 7956 39153
rect 7990 39119 8024 39153
rect 8058 39119 8092 39153
rect 8126 39119 8160 39153
rect 8194 39119 8228 39153
rect 8262 39119 8296 39153
rect 8330 39119 8364 39153
rect 8398 39119 8432 39153
rect 8466 39119 8500 39153
rect 8534 39119 8568 39153
rect 8602 39119 8636 39153
rect 8670 39119 8704 39153
rect 8738 39119 8772 39153
rect 8806 39119 8840 39153
rect 8874 39119 8908 39153
rect 8943 39119 8977 39153
rect 9012 39119 9046 39153
rect 9081 39119 9115 39153
rect 9150 39119 9184 39153
rect 9219 39119 9253 39153
rect 9288 39119 9322 39153
rect 9357 39119 9391 39153
rect 9426 39119 9460 39153
rect 9495 39119 9529 39153
rect 9564 39119 9598 39153
rect 9633 39119 9667 39153
rect 9702 39119 9736 39153
rect 9771 39119 9805 39153
rect 9840 39119 9874 39153
rect 9909 39119 9943 39153
rect 9978 39119 10012 39153
rect 10047 39119 10081 39153
rect 10116 39119 10150 39153
rect 10185 39119 10219 39153
rect 10254 39119 10288 39153
rect 10323 39119 10357 39153
rect 10392 39119 10426 39153
rect 10461 39119 10495 39153
rect 10530 39119 10564 39153
rect 10599 39119 10633 39153
rect 10668 39119 10702 39153
rect 10737 39119 10771 39153
rect 10806 39119 10840 39153
rect 10875 39119 10909 39153
rect 10944 39119 10978 39153
rect 11013 39119 11047 39153
rect 11082 39119 11116 39153
rect 11151 39119 11185 39153
rect 11220 39119 11254 39153
rect 11289 39119 11323 39153
rect 11358 39119 11392 39153
rect 11427 39119 11461 39153
rect 11496 39119 11530 39153
rect 11565 39119 11599 39153
rect 11634 39119 11668 39153
rect 11703 39119 11737 39153
rect 11772 39119 11806 39153
rect 11841 39119 11875 39153
rect 11910 39119 11944 39153
rect 11979 39119 12013 39153
rect 12048 39119 12082 39153
rect 12117 39119 12151 39153
rect 12186 39119 12220 39153
rect 12255 39119 12289 39153
rect 12324 39119 12358 39153
rect 12393 39119 12427 39153
rect 12462 39119 12496 39153
rect 12531 39119 12565 39153
rect 12600 39119 12634 39153
rect 12669 39119 12703 39153
rect 12738 39119 12772 39153
rect 12807 39119 12841 39153
rect 12876 39119 12910 39153
rect 12945 39119 12979 39153
rect 13014 39119 13048 39153
rect 13083 39119 13117 39153
rect 13152 39119 13186 39153
rect 13221 39119 13255 39153
rect 13290 39119 13324 39153
rect 13359 39119 13393 39153
rect 13428 39119 13462 39153
rect 2274 29157 2444 39119
rect 2482 38993 2516 39027
rect 2550 38993 2584 39027
rect 2618 38993 2652 39027
rect 2686 38993 2720 39027
rect 2754 38993 2788 39027
rect 2822 38993 2856 39027
rect 2890 38993 2924 39027
rect 2958 38993 2992 39027
rect 3026 38993 3060 39027
rect 3094 38993 3128 39027
rect 3162 38993 3196 39027
rect 3230 38993 3264 39027
rect 3298 38993 3332 39027
rect 3366 38993 3400 39027
rect 3434 38993 3468 39027
rect 3502 38993 3536 39027
rect 3570 38993 3604 39027
rect 3638 38993 3672 39027
rect 3706 38993 3740 39027
rect 3774 38993 3808 39027
rect 3842 38993 3876 39027
rect 3910 38993 3944 39027
rect 3978 38993 4012 39027
rect 4046 38993 4080 39027
rect 4114 38993 4148 39027
rect 4182 38993 4216 39027
rect 4250 38993 4284 39027
rect 4318 38993 4352 39027
rect 4386 38993 4420 39027
rect 4454 38993 4488 39027
rect 4522 38993 4556 39027
rect 4590 38993 4624 39027
rect 4658 38993 4692 39027
rect 4726 38993 4760 39027
rect 4794 38993 4828 39027
rect 4862 38993 4896 39027
rect 4930 38993 4964 39027
rect 4998 38993 5032 39027
rect 5066 38993 5100 39027
rect 5134 38993 5168 39027
rect 5202 38993 5236 39027
rect 5270 38993 5304 39027
rect 5338 38993 5372 39027
rect 5406 38993 5440 39027
rect 5474 38993 5508 39027
rect 5542 38993 5576 39027
rect 5610 38993 5644 39027
rect 5678 38993 5712 39027
rect 5746 38993 5780 39027
rect 5814 38993 5848 39027
rect 5882 38993 5916 39027
rect 5950 38993 5984 39027
rect 6018 38993 6052 39027
rect 6086 38993 6120 39027
rect 6154 38993 6188 39027
rect 6222 38993 6256 39027
rect 6290 38993 6324 39027
rect 6358 38993 6392 39027
rect 6426 38993 6460 39027
rect 6494 38993 6528 39027
rect 6562 38993 6596 39027
rect 6630 38993 6664 39027
rect 6698 38993 6732 39027
rect 6766 38993 6800 39027
rect 6834 38993 6868 39027
rect 6902 38993 6936 39027
rect 6970 38993 7004 39027
rect 7038 38993 7072 39027
rect 7106 38993 7140 39027
rect 7174 38993 7208 39027
rect 7242 38993 7276 39027
rect 7310 38993 7344 39027
rect 7378 38993 7412 39027
rect 7446 38993 7480 39027
rect 7514 38993 7548 39027
rect 7582 38993 7616 39027
rect 7650 38993 7684 39027
rect 7718 38993 7752 39027
rect 7786 38993 7820 39027
rect 7854 38993 7888 39027
rect 7922 38993 7956 39027
rect 7990 38993 8024 39027
rect 8058 38993 8092 39027
rect 8126 38993 8160 39027
rect 8194 38993 8228 39027
rect 8262 38993 8296 39027
rect 8330 38993 8364 39027
rect 8398 38993 8432 39027
rect 8466 38993 8500 39027
rect 8534 38993 8568 39027
rect 8602 38993 8636 39027
rect 8670 38993 8704 39027
rect 8738 38993 8772 39027
rect 8806 38993 8840 39027
rect 8874 38993 8908 39027
rect 8943 38993 8977 39027
rect 9012 38993 9046 39027
rect 9081 38993 9115 39027
rect 9150 38993 9184 39027
rect 9219 38993 9253 39027
rect 9288 38993 9322 39027
rect 9357 38993 9391 39027
rect 9426 38993 9460 39027
rect 9495 38993 9529 39027
rect 9564 38993 9598 39027
rect 9633 38993 9667 39027
rect 9702 38993 9736 39027
rect 9771 38993 9805 39027
rect 9840 38993 9874 39027
rect 9909 38993 9943 39027
rect 9978 38993 10012 39027
rect 10047 38993 10081 39027
rect 10116 38993 10150 39027
rect 10185 38993 10219 39027
rect 10254 38993 10288 39027
rect 10323 38993 10357 39027
rect 10392 38993 10426 39027
rect 10461 38993 10495 39027
rect 10530 38993 10564 39027
rect 10599 38993 10633 39027
rect 10668 38993 10702 39027
rect 10737 38993 10771 39027
rect 10806 38993 10840 39027
rect 10875 38993 10909 39027
rect 10944 38993 10978 39027
rect 11013 38993 11047 39027
rect 11082 38993 11116 39027
rect 11151 38993 11185 39027
rect 11220 38993 11254 39027
rect 11289 38993 11323 39027
rect 11358 38993 11392 39027
rect 11427 38993 11461 39027
rect 11496 38993 11530 39027
rect 11565 38993 11599 39027
rect 11634 38993 11668 39027
rect 11703 38993 11737 39027
rect 11772 38993 11806 39027
rect 11841 38993 11875 39027
rect 11910 38993 11944 39027
rect 11979 38993 12013 39027
rect 12048 38993 12082 39027
rect 12117 38993 12151 39027
rect 12186 38993 12220 39027
rect 12255 38993 12289 39027
rect 12324 38993 12358 39027
rect 12393 38993 12427 39027
rect 12462 38993 12496 39027
rect 12531 38993 12565 39027
rect 12600 38993 12634 39027
rect 12669 38993 12703 39027
rect 12738 38993 12772 39027
rect 12807 38993 12841 39027
rect 12876 38993 12910 39027
rect 12945 38993 12979 39027
rect 13014 38993 13048 39027
rect 13083 38993 13117 39027
rect 13152 38993 13186 39027
rect 13221 38993 13255 39027
rect 13290 38993 13324 39027
rect 13359 38993 13393 39027
rect 13428 38993 13462 39027
rect 2274 29089 2376 29157
rect 2274 29021 2308 29055
rect 2410 28995 4144 29063
rect 4178 29029 4212 29063
rect 2342 28961 4144 28995
rect 2342 28893 4076 28961
rect 4196 28927 4298 28995
rect 4128 20257 4298 28927
rect 4335 23554 4369 23588
rect 4403 23554 4437 23588
rect 4471 23554 4505 23588
rect 4539 23554 4573 23588
rect 4607 23554 4641 23588
rect 4675 23554 4709 23588
rect 4743 23554 4777 23588
rect 4811 23554 4845 23588
rect 4879 23554 4913 23588
rect 4947 23554 4981 23588
rect 5015 23554 5049 23588
rect 5083 23554 5117 23588
rect 5151 23554 5185 23588
rect 5219 23554 5253 23588
rect 5287 23554 5321 23588
rect 5355 23554 5389 23588
rect 5423 23554 5457 23588
rect 5491 23554 5525 23588
rect 5559 23554 5593 23588
rect 5627 23554 5661 23588
rect 5695 23554 5729 23588
rect 5763 23554 5797 23588
rect 5831 23554 5865 23588
rect 5899 23554 5933 23588
rect 5967 23554 6001 23588
rect 6035 23554 6069 23588
rect 6103 23554 6137 23588
rect 6171 23554 6205 23588
rect 6239 23554 6273 23588
rect 6307 23554 6341 23588
rect 6375 23554 6409 23588
rect 6443 23554 6477 23588
rect 6511 23554 6545 23588
rect 6579 23554 6613 23588
rect 6647 23554 6681 23588
rect 6715 23554 6749 23588
rect 6783 23554 6817 23588
rect 6851 23554 6885 23588
rect 6919 23554 6953 23588
rect 6987 23554 7021 23588
rect 7055 23554 7089 23588
rect 7123 23554 7157 23588
rect 7191 23554 7225 23588
rect 7259 23554 7293 23588
rect 7327 23554 7361 23588
rect 7395 23554 7429 23588
rect 7463 23554 7497 23588
rect 7531 23554 7565 23588
rect 7599 23554 7633 23588
rect 7667 23554 7701 23588
rect 7735 23554 7769 23588
rect 7803 23554 7837 23588
rect 7871 23554 7905 23588
rect 7939 23554 7973 23588
rect 8007 23554 8041 23588
rect 8075 23554 8109 23588
rect 8143 23554 8177 23588
rect 8211 23554 8245 23588
rect 8279 23554 8313 23588
rect 8347 23554 8381 23588
rect 8415 23554 8449 23588
rect 8483 23554 8517 23588
rect 8551 23554 8585 23588
rect 8619 23554 8653 23588
rect 8687 23554 8721 23588
rect 8755 23554 8789 23588
rect 8823 23554 8857 23588
rect 8891 23554 8925 23588
rect 8959 23554 8993 23588
rect 9027 23554 9061 23588
rect 9095 23554 9129 23588
rect 9163 23554 9197 23588
rect 9231 23554 9265 23588
rect 9299 23554 9333 23588
rect 9367 23554 9401 23588
rect 9435 23554 9469 23588
rect 9503 23554 9537 23588
rect 9571 23554 9605 23588
rect 9639 23554 9673 23588
rect 9707 23554 9741 23588
rect 9775 23554 9809 23588
rect 9843 23554 9877 23588
rect 9911 23554 9945 23588
rect 9979 23554 10013 23588
rect 10047 23554 10081 23588
rect 10115 23554 10149 23588
rect 10183 23554 10217 23588
rect 10251 23554 10285 23588
rect 10319 23554 10353 23588
rect 10387 23554 10421 23588
rect 10455 23554 10489 23588
rect 10523 23554 10557 23588
rect 10591 23554 10625 23588
rect 10659 23554 10693 23588
rect 10727 23554 10761 23588
rect 10795 23554 10829 23588
rect 10863 23554 10897 23588
rect 10931 23554 10965 23588
rect 10999 23554 11033 23588
rect 11067 23554 11101 23588
rect 11135 23554 11169 23588
rect 11203 23554 11237 23588
rect 11271 23554 11305 23588
rect 11339 23554 11373 23588
rect 11407 23554 11441 23588
rect 11475 23554 11509 23588
rect 11543 23554 11577 23588
rect 11611 23554 11645 23588
rect 11679 23554 11713 23588
rect 11747 23554 11781 23588
rect 11815 23554 11849 23588
rect 11883 23554 11917 23588
rect 11951 23554 11985 23588
rect 12019 23554 12053 23588
rect 12087 23554 12121 23588
rect 12155 23554 12189 23588
rect 12223 23554 12257 23588
rect 12291 23554 12325 23588
rect 12359 23554 12393 23588
rect 12427 23554 12461 23588
rect 12495 23554 12529 23588
rect 12563 23554 12597 23588
rect 12631 23554 12665 23588
rect 12699 23554 12733 23588
rect 12767 23554 12801 23588
rect 12835 23554 12869 23588
rect 12903 23554 12937 23588
rect 12971 23554 13005 23588
rect 13039 23554 13073 23588
rect 13107 23554 13141 23588
rect 13175 23554 13209 23588
rect 13243 23554 13277 23588
rect 13311 23554 13345 23588
rect 13379 23554 13413 23588
rect 13447 23554 13481 23588
rect 4335 21855 4369 21889
rect 4403 21855 4437 21889
rect 4471 21855 4505 21889
rect 4539 21855 4573 21889
rect 4607 21855 4641 21889
rect 4675 21855 4709 21889
rect 4743 21855 4777 21889
rect 4811 21855 4845 21889
rect 4879 21855 4913 21889
rect 4947 21855 4981 21889
rect 5015 21855 5049 21889
rect 5083 21855 5117 21889
rect 5151 21855 5185 21889
rect 5219 21855 5253 21889
rect 5287 21855 5321 21889
rect 5355 21855 5389 21889
rect 5423 21855 5457 21889
rect 5491 21855 5525 21889
rect 5559 21855 5593 21889
rect 5627 21855 5661 21889
rect 5695 21855 5729 21889
rect 5763 21855 5797 21889
rect 5831 21855 5865 21889
rect 5899 21855 5933 21889
rect 5967 21855 6001 21889
rect 6035 21855 6069 21889
rect 6103 21855 6137 21889
rect 6171 21855 6205 21889
rect 6239 21855 6273 21889
rect 6307 21855 6341 21889
rect 6375 21855 6409 21889
rect 6443 21855 6477 21889
rect 6511 21855 6545 21889
rect 6579 21855 6613 21889
rect 6647 21855 6681 21889
rect 6715 21855 6749 21889
rect 6783 21855 6817 21889
rect 6851 21855 6885 21889
rect 6919 21855 6953 21889
rect 6987 21855 7021 21889
rect 7055 21855 7089 21889
rect 7123 21855 7157 21889
rect 7191 21855 7225 21889
rect 7259 21855 7293 21889
rect 7327 21855 7361 21889
rect 7395 21855 7429 21889
rect 7463 21855 7497 21889
rect 7531 21855 7565 21889
rect 7599 21855 7633 21889
rect 7667 21855 7701 21889
rect 7735 21855 7769 21889
rect 7803 21855 7837 21889
rect 7871 21855 7905 21889
rect 7939 21855 7973 21889
rect 8007 21855 8041 21889
rect 8075 21855 8109 21889
rect 8143 21855 8177 21889
rect 8211 21855 8245 21889
rect 8279 21855 8313 21889
rect 8347 21855 8381 21889
rect 8415 21855 8449 21889
rect 8483 21855 8517 21889
rect 8551 21855 8585 21889
rect 8619 21855 8653 21889
rect 8687 21855 8721 21889
rect 8755 21855 8789 21889
rect 8823 21855 8857 21889
rect 8891 21855 8925 21889
rect 8959 21855 8993 21889
rect 9027 21855 9061 21889
rect 9095 21855 9129 21889
rect 9163 21855 9197 21889
rect 9231 21855 9265 21889
rect 9299 21855 9333 21889
rect 9367 21855 9401 21889
rect 9435 21855 9469 21889
rect 9503 21855 9537 21889
rect 9571 21855 9605 21889
rect 9639 21855 9673 21889
rect 9707 21855 9741 21889
rect 9775 21855 9809 21889
rect 9843 21855 9877 21889
rect 9911 21855 9945 21889
rect 9979 21855 10013 21889
rect 10047 21855 10081 21889
rect 10115 21855 10149 21889
rect 10183 21855 10217 21889
rect 10251 21855 10285 21889
rect 10319 21855 10353 21889
rect 10387 21855 10421 21889
rect 10455 21855 10489 21889
rect 10523 21855 10557 21889
rect 10591 21855 10625 21889
rect 10659 21855 10693 21889
rect 10727 21855 10761 21889
rect 10795 21855 10829 21889
rect 10863 21855 10897 21889
rect 10931 21855 10965 21889
rect 10999 21855 11033 21889
rect 11067 21855 11101 21889
rect 11135 21855 11169 21889
rect 11203 21855 11237 21889
rect 11271 21855 11305 21889
rect 11339 21855 11373 21889
rect 11407 21855 11441 21889
rect 11475 21855 11509 21889
rect 11543 21855 11577 21889
rect 11611 21855 11645 21889
rect 11679 21855 11713 21889
rect 11747 21855 11781 21889
rect 11815 21855 11849 21889
rect 11883 21855 11917 21889
rect 11951 21855 11985 21889
rect 12019 21855 12053 21889
rect 12087 21855 12121 21889
rect 12155 21855 12189 21889
rect 12223 21855 12257 21889
rect 12291 21855 12325 21889
rect 12359 21855 12393 21889
rect 12427 21855 12461 21889
rect 12495 21855 12529 21889
rect 12563 21855 12597 21889
rect 12631 21855 12665 21889
rect 12699 21855 12733 21889
rect 12767 21855 12801 21889
rect 12835 21855 12869 21889
rect 12903 21855 12937 21889
rect 12971 21855 13005 21889
rect 13039 21855 13073 21889
rect 13107 21855 13141 21889
rect 13175 21855 13209 21889
rect 13243 21855 13277 21889
rect 13311 21855 13345 21889
rect 13379 21855 13413 21889
rect 13447 21855 13481 21889
rect 13515 20531 13617 39129
rect 13515 20462 13549 20496
rect 13583 20462 13617 20496
rect 13515 20393 13549 20427
rect 13583 20393 13617 20427
rect 13515 20324 13549 20358
rect 13583 20324 13617 20358
rect 13515 20255 13549 20289
rect 13583 20255 13617 20289
rect 4152 20173 4186 20207
rect 4221 20173 4255 20207
rect 4290 20173 4324 20207
rect 4359 20173 4393 20207
rect 4428 20173 4462 20207
rect 4497 20173 4531 20207
rect 4566 20173 4600 20207
rect 4635 20173 4669 20207
rect 4704 20173 4738 20207
rect 4773 20173 4807 20207
rect 4842 20173 4876 20207
rect 4911 20173 4945 20207
rect 4980 20173 5014 20207
rect 5049 20173 5083 20207
rect 5118 20173 5152 20207
rect 5187 20173 5221 20207
rect 5256 20173 5290 20207
rect 5325 20173 5359 20207
rect 5394 20173 5428 20207
rect 5463 20173 5497 20207
rect 5532 20173 5566 20207
rect 5601 20173 5635 20207
rect 5670 20173 5704 20207
rect 5739 20173 5773 20207
rect 5807 20173 5841 20207
rect 5875 20173 5909 20207
rect 5943 20173 5977 20207
rect 6011 20173 6045 20207
rect 6079 20173 6113 20207
rect 6147 20173 6181 20207
rect 6215 20173 6249 20207
rect 6283 20173 6317 20207
rect 6351 20173 6385 20207
rect 6419 20173 6453 20207
rect 6487 20173 6521 20207
rect 6555 20173 6589 20207
rect 6623 20173 6657 20207
rect 6691 20173 6725 20207
rect 6759 20173 6793 20207
rect 6827 20173 6861 20207
rect 6895 20173 6929 20207
rect 6963 20173 6997 20207
rect 7031 20173 7065 20207
rect 7099 20173 7133 20207
rect 7167 20173 7201 20207
rect 7235 20173 7269 20207
rect 7303 20173 7337 20207
rect 7371 20173 7405 20207
rect 7439 20173 7473 20207
rect 7507 20173 7541 20207
rect 7575 20173 7609 20207
rect 7643 20173 7677 20207
rect 7711 20173 7745 20207
rect 7779 20173 7813 20207
rect 7847 20173 7881 20207
rect 7915 20173 7949 20207
rect 7983 20173 8017 20207
rect 8051 20173 8085 20207
rect 8119 20173 8153 20207
rect 8187 20173 8221 20207
rect 8255 20173 8289 20207
rect 8323 20173 8357 20207
rect 8391 20173 8425 20207
rect 8459 20173 8493 20207
rect 8527 20173 8561 20207
rect 8595 20173 8629 20207
rect 8663 20173 8697 20207
rect 8731 20173 8765 20207
rect 8799 20173 8833 20207
rect 8867 20173 8901 20207
rect 8935 20173 8969 20207
rect 9003 20173 9037 20207
rect 9071 20173 9105 20207
rect 9139 20173 9173 20207
rect 9207 20173 9241 20207
rect 9275 20173 9309 20207
rect 9343 20173 9377 20207
rect 9411 20173 9445 20207
rect 9479 20173 9513 20207
rect 9547 20173 9581 20207
rect 9615 20173 9649 20207
rect 9683 20173 9717 20207
rect 9751 20173 9785 20207
rect 9819 20173 9853 20207
rect 9887 20173 9921 20207
rect 9955 20173 9989 20207
rect 10023 20173 10057 20207
rect 10091 20173 10125 20207
rect 10159 20173 10193 20207
rect 10227 20173 10261 20207
rect 10295 20173 10329 20207
rect 10363 20173 10397 20207
rect 10431 20173 10465 20207
rect 10499 20173 10533 20207
rect 10567 20173 10601 20207
rect 10635 20173 10669 20207
rect 10703 20173 10737 20207
rect 10771 20173 10805 20207
rect 10839 20173 10873 20207
rect 10907 20173 10941 20207
rect 10975 20173 11009 20207
rect 11043 20173 11077 20207
rect 11111 20173 11145 20207
rect 11179 20173 11213 20207
rect 11247 20173 11281 20207
rect 11315 20173 11349 20207
rect 11383 20173 11417 20207
rect 11451 20173 11485 20207
rect 11519 20173 11553 20207
rect 11587 20173 11621 20207
rect 11655 20173 11689 20207
rect 11723 20173 11757 20207
rect 11791 20173 11825 20207
rect 11859 20173 11893 20207
rect 11927 20173 11961 20207
rect 11995 20173 12029 20207
rect 12063 20173 12097 20207
rect 12131 20173 12165 20207
rect 12199 20173 12233 20207
rect 12267 20173 12301 20207
rect 12335 20173 12369 20207
rect 12403 20173 12437 20207
rect 12471 20173 12505 20207
rect 12539 20173 12573 20207
rect 12607 20173 12641 20207
rect 12675 20173 12709 20207
rect 12743 20173 12777 20207
rect 12811 20173 12845 20207
rect 12879 20173 12913 20207
rect 12947 20173 12981 20207
rect 13015 20173 13049 20207
rect 13083 20173 13117 20207
rect 13151 20173 13185 20207
rect 13219 20173 13253 20207
rect 13287 20173 13321 20207
rect 13355 20173 13389 20207
rect 13423 20173 13457 20207
rect 13491 20173 13525 20207
rect 13559 20173 13593 20207
rect 4578 19798 4612 19832
rect 4647 19798 4681 19832
rect 4716 19798 4750 19832
rect 4785 19798 4819 19832
rect 4854 19798 4888 19832
rect 4923 19798 4957 19832
rect 4992 19798 5026 19832
rect 5061 19798 5095 19832
rect 5130 19798 5164 19832
rect 5199 19798 5233 19832
rect 5268 19798 5302 19832
rect 5337 19798 5371 19832
rect 5406 19798 5440 19832
rect 5475 19798 5509 19832
rect 5544 19798 5578 19832
rect 5613 19798 5647 19832
rect 5682 19798 5716 19832
rect 5750 19798 5784 19832
rect 5818 19798 5852 19832
rect 5886 19798 5920 19832
rect 5954 19798 5988 19832
rect 6022 19798 6056 19832
rect 6090 19798 6124 19832
rect 6158 19798 6192 19832
rect 6226 19798 6260 19832
rect 6294 19798 6328 19832
rect 6362 19798 6396 19832
rect 6430 19798 6464 19832
rect 6498 19798 6532 19832
rect 6566 19798 6600 19832
rect 6634 19798 6668 19832
rect 6702 19798 6736 19832
rect 6770 19798 6804 19832
rect 6838 19798 6872 19832
rect 6906 19798 6940 19832
rect 6974 19798 7008 19832
rect 7042 19798 7076 19832
rect 7110 19798 7144 19832
rect 7178 19798 7212 19832
rect 7246 19798 7280 19832
rect 7314 19798 7348 19832
rect 7382 19798 7416 19832
rect 7450 19798 7484 19832
rect 7518 19798 7552 19832
rect 7586 19798 7620 19832
rect 7654 19798 7688 19832
rect 7722 19798 7756 19832
rect 7790 19798 7824 19832
rect 7858 19798 7892 19832
rect 7926 19798 7960 19832
rect 7994 19798 8028 19832
rect 8062 19798 8096 19832
rect 8130 19798 8164 19832
rect 8198 19798 8232 19832
rect 8266 19798 8300 19832
rect 8334 19798 8368 19832
rect 8402 19798 8436 19832
rect 8470 19798 8504 19832
rect 8538 19798 8572 19832
rect 8606 19798 8640 19832
rect 8674 19798 8708 19832
rect 8742 19798 8776 19832
rect 8810 19798 8844 19832
rect 8878 19798 8912 19832
rect 8946 19798 8980 19832
rect 9014 19798 9048 19832
rect 9082 19798 9116 19832
rect 9150 19798 9184 19832
rect 9218 19798 9252 19832
rect 9286 19798 9320 19832
rect 9354 19798 9388 19832
rect 9422 19798 9456 19832
rect 9490 19798 9524 19832
rect 9558 19798 9592 19832
rect 9626 19798 9660 19832
rect 9694 19798 9728 19832
rect 9762 19798 9796 19832
rect 9830 19798 9864 19832
rect 9898 19798 9932 19832
rect 9966 19798 10000 19832
rect 10034 19798 10068 19832
rect 10102 19798 10136 19832
rect 10170 19798 10204 19832
rect 10238 19798 10272 19832
rect 10306 19798 10340 19832
rect 10374 19798 10408 19832
rect 10442 19798 10476 19832
rect 10510 19798 10544 19832
rect 10578 19798 10612 19832
rect 10646 19798 10680 19832
rect 10714 19798 10748 19832
rect 10782 19798 10816 19832
rect 10850 19798 10884 19832
rect 10918 19798 10952 19832
rect 10986 19798 11020 19832
rect 11054 19798 11088 19832
rect 11122 19798 11156 19832
rect 11190 19798 11224 19832
rect 11258 19798 11292 19832
rect 11326 19798 11360 19832
rect 11394 19798 11428 19832
rect 11462 19798 11496 19832
rect 11530 19798 11564 19832
rect 11598 19798 11632 19832
rect 11666 19798 11700 19832
rect 11734 19798 11768 19832
rect 11802 19798 11836 19832
rect 11870 19798 11904 19832
rect 11938 19798 11972 19832
rect 12006 19798 12040 19832
rect 12074 19798 12108 19832
rect 12142 19798 12176 19832
rect 12210 19798 12244 19832
rect 12278 19798 12312 19832
rect 12346 19798 12380 19832
rect 12414 19798 12448 19832
rect 12482 19798 12516 19832
rect 12550 19798 12584 19832
rect 12618 19798 12652 19832
rect 12686 19798 12720 19832
rect 12754 19798 12788 19832
rect 12822 19798 12856 19832
rect 12890 19798 12924 19832
rect 12958 19798 12992 19832
rect 13026 19798 13060 19832
rect 13094 19798 13128 19832
rect 13162 19798 13196 19832
rect 13230 19798 13264 19832
rect 13298 19798 13332 19832
rect 13366 19798 13400 19832
rect 13434 19798 13468 19832
rect 13502 19798 13536 19832
rect 13570 19798 13604 19832
rect 4554 16466 4656 19764
rect 4754 18135 4788 18169
rect 4822 18135 4856 18169
rect 4890 18135 4924 18169
rect 4958 18135 4992 18169
rect 5026 18135 5060 18169
rect 5094 18135 5128 18169
rect 5162 18135 5196 18169
rect 5230 18135 5264 18169
rect 5298 18135 5332 18169
rect 5366 18135 5400 18169
rect 5434 18135 5468 18169
rect 5502 18135 5536 18169
rect 5570 18135 5604 18169
rect 5638 18135 5672 18169
rect 5706 18135 5740 18169
rect 5774 18135 5808 18169
rect 5842 18135 5876 18169
rect 5910 18135 5944 18169
rect 5978 18135 6012 18169
rect 6046 18135 6080 18169
rect 6114 18135 6148 18169
rect 6182 18135 6216 18169
rect 6250 18135 6284 18169
rect 6318 18135 6352 18169
rect 6386 18135 6420 18169
rect 6454 18135 6488 18169
rect 6522 18135 6556 18169
rect 6590 18135 6624 18169
rect 6658 18135 6692 18169
rect 6726 18135 6760 18169
rect 6794 18135 6828 18169
rect 6862 18135 6896 18169
rect 6930 18135 6964 18169
rect 6998 18135 7032 18169
rect 7066 18135 7100 18169
rect 7134 18135 7168 18169
rect 7202 18135 7236 18169
rect 7270 18135 7304 18169
rect 7338 18135 7372 18169
rect 7406 18135 7440 18169
rect 7474 18135 7508 18169
rect 7542 18135 7576 18169
rect 7610 18135 7644 18169
rect 7678 18135 7712 18169
rect 7746 18135 7780 18169
rect 7814 18135 7848 18169
rect 7882 18135 7916 18169
rect 7950 18135 7984 18169
rect 8018 18135 8052 18169
rect 8086 18135 8120 18169
rect 8154 18135 8188 18169
rect 8222 18135 8256 18169
rect 8290 18135 8324 18169
rect 8358 18135 8392 18169
rect 8426 18135 8460 18169
rect 8494 18135 8528 18169
rect 8562 18135 8596 18169
rect 8630 18135 8664 18169
rect 8698 18135 8732 18169
rect 8766 18135 8800 18169
rect 8834 18135 8868 18169
rect 8902 18135 8936 18169
rect 8970 18135 9004 18169
rect 9038 18135 9072 18169
rect 9106 18135 9140 18169
rect 9174 18135 9208 18169
rect 9242 18135 9276 18169
rect 9310 18135 9344 18169
rect 9378 18135 9412 18169
rect 9446 18135 9480 18169
rect 9514 18135 9548 18169
rect 9582 18135 9616 18169
rect 9650 18135 9684 18169
rect 9718 18135 9752 18169
rect 9786 18135 9820 18169
rect 9854 18135 9888 18169
rect 9922 18135 9956 18169
rect 9990 18135 10024 18169
rect 10058 18135 10092 18169
rect 10126 18135 10160 18169
rect 10194 18135 10228 18169
rect 10262 18135 10296 18169
rect 10330 18135 10364 18169
rect 10398 18135 10432 18169
rect 10466 18135 10500 18169
rect 10534 18135 10568 18169
rect 10602 18135 10636 18169
rect 10670 18135 10704 18169
rect 10738 18135 10772 18169
rect 10806 18135 10840 18169
rect 10874 18135 10908 18169
rect 10942 18135 10976 18169
rect 11010 18135 11044 18169
rect 11078 18135 11112 18169
rect 11146 18135 11180 18169
rect 11214 18135 11248 18169
rect 11282 18135 11316 18169
rect 11350 18135 11384 18169
rect 11418 18135 11452 18169
rect 11486 18135 11520 18169
rect 11554 18135 11588 18169
rect 11622 18135 11656 18169
rect 11690 18135 11724 18169
rect 11758 18135 11792 18169
rect 11826 18135 11860 18169
rect 11894 18135 11928 18169
rect 11962 18135 11996 18169
rect 12030 18135 12064 18169
rect 12098 18135 12132 18169
rect 12166 18135 12200 18169
rect 12234 18135 12268 18169
rect 12302 18135 12336 18169
rect 12370 18135 12404 18169
rect 12438 18135 12472 18169
rect 12506 18135 12540 18169
rect 12574 18135 12608 18169
rect 12642 18135 12676 18169
rect 12710 18135 12744 18169
rect 12778 18135 12812 18169
rect 12846 18135 12880 18169
rect 12914 18135 12948 18169
rect 12982 18135 13016 18169
rect 13050 18135 13084 18169
rect 13118 18135 13152 18169
rect 13186 18135 13220 18169
rect 13254 18135 13288 18169
rect 13322 18135 13356 18169
rect 13390 18135 13424 18169
rect 4754 16436 4788 16470
rect 4822 16436 4856 16470
rect 4890 16436 4924 16470
rect 4958 16436 4992 16470
rect 5026 16436 5060 16470
rect 5094 16436 5128 16470
rect 5162 16436 5196 16470
rect 5230 16436 5264 16470
rect 5298 16436 5332 16470
rect 5366 16436 5400 16470
rect 5434 16436 5468 16470
rect 5502 16436 5536 16470
rect 5570 16436 5604 16470
rect 5638 16436 5672 16470
rect 5706 16436 5740 16470
rect 5774 16436 5808 16470
rect 5842 16436 5876 16470
rect 5910 16436 5944 16470
rect 5978 16436 6012 16470
rect 6046 16436 6080 16470
rect 6114 16436 6148 16470
rect 6182 16436 6216 16470
rect 6250 16436 6284 16470
rect 6318 16436 6352 16470
rect 6386 16436 6420 16470
rect 6454 16436 6488 16470
rect 6522 16436 6556 16470
rect 6590 16436 6624 16470
rect 6658 16436 6692 16470
rect 6726 16436 6760 16470
rect 6794 16436 6828 16470
rect 6862 16436 6896 16470
rect 6930 16436 6964 16470
rect 6998 16436 7032 16470
rect 7066 16436 7100 16470
rect 7134 16436 7168 16470
rect 7202 16436 7236 16470
rect 7270 16436 7304 16470
rect 7338 16436 7372 16470
rect 7406 16436 7440 16470
rect 7474 16436 7508 16470
rect 7542 16436 7576 16470
rect 7610 16436 7644 16470
rect 7678 16436 7712 16470
rect 7746 16436 7780 16470
rect 7814 16436 7848 16470
rect 7882 16436 7916 16470
rect 7950 16436 7984 16470
rect 8018 16436 8052 16470
rect 8086 16436 8120 16470
rect 8154 16436 8188 16470
rect 8222 16436 8256 16470
rect 8290 16436 8324 16470
rect 8358 16436 8392 16470
rect 8426 16436 8460 16470
rect 8494 16436 8528 16470
rect 8562 16436 8596 16470
rect 8630 16436 8664 16470
rect 8698 16436 8732 16470
rect 8766 16436 8800 16470
rect 8834 16436 8868 16470
rect 8902 16436 8936 16470
rect 8970 16436 9004 16470
rect 9038 16436 9072 16470
rect 9106 16436 9140 16470
rect 9174 16436 9208 16470
rect 9242 16436 9276 16470
rect 9310 16436 9344 16470
rect 9378 16436 9412 16470
rect 9446 16436 9480 16470
rect 9514 16436 9548 16470
rect 9582 16436 9616 16470
rect 9650 16436 9684 16470
rect 9718 16436 9752 16470
rect 9786 16436 9820 16470
rect 9854 16436 9888 16470
rect 9922 16436 9956 16470
rect 9990 16436 10024 16470
rect 10058 16436 10092 16470
rect 10126 16436 10160 16470
rect 10194 16436 10228 16470
rect 10262 16436 10296 16470
rect 10330 16436 10364 16470
rect 10398 16436 10432 16470
rect 10466 16436 10500 16470
rect 10534 16436 10568 16470
rect 10602 16436 10636 16470
rect 10670 16436 10704 16470
rect 10738 16436 10772 16470
rect 10806 16436 10840 16470
rect 10874 16436 10908 16470
rect 10942 16436 10976 16470
rect 11010 16436 11044 16470
rect 11078 16436 11112 16470
rect 11146 16436 11180 16470
rect 11214 16436 11248 16470
rect 11282 16436 11316 16470
rect 11350 16436 11384 16470
rect 11418 16436 11452 16470
rect 11486 16436 11520 16470
rect 11554 16436 11588 16470
rect 11622 16436 11656 16470
rect 11690 16436 11724 16470
rect 11758 16436 11792 16470
rect 11826 16436 11860 16470
rect 11894 16436 11928 16470
rect 11962 16436 11996 16470
rect 12030 16436 12064 16470
rect 12098 16436 12132 16470
rect 12166 16436 12200 16470
rect 12234 16436 12268 16470
rect 12302 16436 12336 16470
rect 12370 16436 12404 16470
rect 12438 16436 12472 16470
rect 12506 16436 12540 16470
rect 12574 16436 12608 16470
rect 12642 16436 12676 16470
rect 12710 16436 12744 16470
rect 12778 16436 12812 16470
rect 12846 16436 12880 16470
rect 12914 16436 12948 16470
rect 12982 16436 13016 16470
rect 13050 16436 13084 16470
rect 13118 16436 13152 16470
rect 13186 16436 13220 16470
rect 13254 16436 13288 16470
rect 13322 16436 13356 16470
rect 13390 16436 13424 16470
rect 2274 5183 2444 16383
rect 2514 16315 4588 16417
rect 4622 16398 4656 16432
rect 2274 5129 13392 5183
rect 2478 5081 13392 5129
rect 13458 5115 13628 19701
rect 1677 3612 1711 3646
rect 1747 3612 1781 3646
rect 1817 3612 1851 3646
rect 1887 3612 1921 3646
rect 1957 3612 1991 3646
rect 2027 3612 2061 3646
rect 2097 3612 2131 3646
rect 2167 3612 2201 3646
rect 2237 3612 2271 3646
rect 2307 3612 2341 3646
rect 2377 3612 2411 3646
rect 2447 3612 2481 3646
rect 2517 3612 2551 3646
rect 2587 3612 2621 3646
rect 2657 3612 2691 3646
rect 2727 3612 2761 3646
rect 2797 3612 2831 3646
rect 2867 3612 2901 3646
rect 2937 3612 2971 3646
rect 3007 3612 3041 3646
rect 3077 3612 3111 3646
rect 3147 3612 3181 3646
rect 3217 3612 3251 3646
rect 3287 3612 3321 3646
rect 1677 3544 1711 3578
rect 1747 3544 1781 3578
rect 1817 3544 1851 3578
rect 1887 3544 1921 3578
rect 1957 3544 1991 3578
rect 2027 3544 2061 3578
rect 2097 3544 2131 3578
rect 2167 3544 2201 3578
rect 2237 3544 2271 3578
rect 2307 3544 2341 3578
rect 2377 3544 2411 3578
rect 2447 3544 2481 3578
rect 2517 3544 2551 3578
rect 2587 3544 2621 3578
rect 2657 3544 2691 3578
rect 2727 3544 2761 3578
rect 2797 3544 2831 3578
rect 2867 3544 2901 3578
rect 2937 3544 2971 3578
rect 3007 3544 3041 3578
rect 3077 3544 3111 3578
rect 3147 3544 3181 3578
rect 3217 3544 3251 3578
rect 3287 3544 3321 3578
rect 1677 3476 1711 3510
rect 1747 3476 1781 3510
rect 1817 3476 1851 3510
rect 1887 3476 1921 3510
rect 1957 3476 1991 3510
rect 2027 3476 2061 3510
rect 2097 3476 2131 3510
rect 2167 3476 2201 3510
rect 2237 3476 2271 3510
rect 2307 3476 2341 3510
rect 2377 3476 2411 3510
rect 2447 3476 2481 3510
rect 2517 3476 2551 3510
rect 2587 3476 2621 3510
rect 2657 3476 2691 3510
rect 2727 3476 2761 3510
rect 2797 3476 2831 3510
rect 2867 3476 2901 3510
rect 2937 3476 2971 3510
rect 3007 3476 3041 3510
rect 3077 3476 3111 3510
rect 3147 3476 3181 3510
rect 3217 3476 3251 3510
rect 3287 3476 3321 3510
rect 1677 3408 1711 3442
rect 1747 3408 1781 3442
rect 1817 3408 1851 3442
rect 1887 3408 1921 3442
rect 1957 3408 1991 3442
rect 2027 3408 2061 3442
rect 2097 3408 2131 3442
rect 2167 3408 2201 3442
rect 2237 3408 2271 3442
rect 2307 3408 2341 3442
rect 2377 3408 2411 3442
rect 2447 3408 2481 3442
rect 2517 3408 2551 3442
rect 2587 3408 2621 3442
rect 2657 3408 2691 3442
rect 2727 3408 2761 3442
rect 2797 3408 2831 3442
rect 2867 3408 2901 3442
rect 2937 3408 2971 3442
rect 3007 3408 3041 3442
rect 3077 3408 3111 3442
rect 3147 3408 3181 3442
rect 3217 3408 3251 3442
rect 3287 3408 3321 3442
rect 1677 3340 1711 3374
rect 1747 3340 1781 3374
rect 1817 3340 1851 3374
rect 1887 3340 1921 3374
rect 1957 3340 1991 3374
rect 2027 3340 2061 3374
rect 2097 3340 2131 3374
rect 2167 3340 2201 3374
rect 2237 3340 2271 3374
rect 2307 3340 2341 3374
rect 2377 3340 2411 3374
rect 2447 3340 2481 3374
rect 2517 3340 2551 3374
rect 2587 3340 2621 3374
rect 2657 3340 2691 3374
rect 2727 3340 2761 3374
rect 2797 3340 2831 3374
rect 2867 3340 2901 3374
rect 2937 3340 2971 3374
rect 3007 3340 3041 3374
rect 3077 3340 3111 3374
rect 3147 3340 3181 3374
rect 3217 3340 3251 3374
rect 3287 3340 3321 3374
rect 1677 3272 1711 3306
rect 1747 3272 1781 3306
rect 1817 3272 1851 3306
rect 1887 3272 1921 3306
rect 1957 3272 1991 3306
rect 2027 3272 2061 3306
rect 2097 3272 2131 3306
rect 2167 3272 2201 3306
rect 2237 3272 2271 3306
rect 2307 3272 2341 3306
rect 2377 3272 2411 3306
rect 2447 3272 2481 3306
rect 2517 3272 2551 3306
rect 2587 3272 2621 3306
rect 2657 3272 2691 3306
rect 2727 3272 2761 3306
rect 2797 3272 2831 3306
rect 2867 3272 2901 3306
rect 2937 3272 2971 3306
rect 3007 3272 3041 3306
rect 3077 3272 3111 3306
rect 3147 3272 3181 3306
rect 3217 3272 3251 3306
rect 3287 3272 3321 3306
rect 1677 3204 1711 3238
rect 1747 3204 1781 3238
rect 1817 3204 1851 3238
rect 1887 3204 1921 3238
rect 1957 3204 1991 3238
rect 2027 3204 2061 3238
rect 2097 3204 2131 3238
rect 2167 3204 2201 3238
rect 2237 3204 2271 3238
rect 2307 3204 2341 3238
rect 2377 3204 2411 3238
rect 2447 3204 2481 3238
rect 2517 3204 2551 3238
rect 2587 3204 2621 3238
rect 2657 3204 2691 3238
rect 2727 3204 2761 3238
rect 2797 3204 2831 3238
rect 2867 3204 2901 3238
rect 2937 3204 2971 3238
rect 3007 3204 3041 3238
rect 3077 3204 3111 3238
rect 3147 3204 3181 3238
rect 3217 3204 3251 3238
rect 3287 3204 3321 3238
rect 1677 3135 1711 3169
rect 1747 3135 1781 3169
rect 1817 3135 1851 3169
rect 1887 3135 1921 3169
rect 1957 3135 1991 3169
rect 2027 3135 2061 3169
rect 2097 3135 2131 3169
rect 2167 3135 2201 3169
rect 2237 3135 2271 3169
rect 2307 3135 2341 3169
rect 2377 3135 2411 3169
rect 2447 3135 2481 3169
rect 2517 3135 2551 3169
rect 2587 3135 2621 3169
rect 2657 3135 2691 3169
rect 2727 3135 2761 3169
rect 2797 3135 2831 3169
rect 2867 3135 2901 3169
rect 2937 3135 2971 3169
rect 3007 3135 3041 3169
rect 3077 3135 3111 3169
rect 3147 3135 3181 3169
rect 3217 3135 3251 3169
rect 3287 3135 3321 3169
rect 1677 3066 1711 3100
rect 1747 3066 1781 3100
rect 1817 3066 1851 3100
rect 1887 3066 1921 3100
rect 1957 3066 1991 3100
rect 2027 3066 2061 3100
rect 2097 3066 2131 3100
rect 2167 3066 2201 3100
rect 2237 3066 2271 3100
rect 2307 3066 2341 3100
rect 2377 3066 2411 3100
rect 2447 3066 2481 3100
rect 2517 3066 2551 3100
rect 2587 3066 2621 3100
rect 2657 3066 2691 3100
rect 2727 3066 2761 3100
rect 2797 3066 2831 3100
rect 2867 3066 2901 3100
rect 2937 3066 2971 3100
rect 3007 3066 3041 3100
rect 3077 3066 3111 3100
rect 3147 3066 3181 3100
rect 3217 3066 3251 3100
rect 3287 3066 3321 3100
rect 1677 2997 1711 3031
rect 1747 2997 1781 3031
rect 1817 2997 1851 3031
rect 1887 2997 1921 3031
rect 1957 2997 1991 3031
rect 2027 2997 2061 3031
rect 2097 2997 2131 3031
rect 2167 2997 2201 3031
rect 2237 2997 2271 3031
rect 2307 2997 2341 3031
rect 2377 2997 2411 3031
rect 2447 2997 2481 3031
rect 2517 2997 2551 3031
rect 2587 2997 2621 3031
rect 2657 2997 2691 3031
rect 2727 2997 2761 3031
rect 2797 2997 2831 3031
rect 2867 2997 2901 3031
rect 2937 2997 2971 3031
rect 3007 2997 3041 3031
rect 3077 2997 3111 3031
rect 3147 2997 3181 3031
rect 3217 2997 3251 3031
rect 3287 2997 3321 3031
rect 1677 2928 1711 2962
rect 1747 2928 1781 2962
rect 1817 2928 1851 2962
rect 1887 2928 1921 2962
rect 1957 2928 1991 2962
rect 2027 2928 2061 2962
rect 2097 2928 2131 2962
rect 2167 2928 2201 2962
rect 2237 2928 2271 2962
rect 2307 2928 2341 2962
rect 2377 2928 2411 2962
rect 2447 2928 2481 2962
rect 2517 2928 2551 2962
rect 2587 2928 2621 2962
rect 2657 2928 2691 2962
rect 2727 2928 2761 2962
rect 2797 2928 2831 2962
rect 2867 2928 2901 2962
rect 2937 2928 2971 2962
rect 3007 2928 3041 2962
rect 3077 2928 3111 2962
rect 3147 2928 3181 2962
rect 3217 2928 3251 2962
rect 3287 2928 3321 2962
rect 1677 2859 1711 2893
rect 1747 2859 1781 2893
rect 1817 2859 1851 2893
rect 1887 2859 1921 2893
rect 1957 2859 1991 2893
rect 2027 2859 2061 2893
rect 2097 2859 2131 2893
rect 2167 2859 2201 2893
rect 2237 2859 2271 2893
rect 2307 2859 2341 2893
rect 2377 2859 2411 2893
rect 2447 2859 2481 2893
rect 2517 2859 2551 2893
rect 2587 2859 2621 2893
rect 2657 2859 2691 2893
rect 2727 2859 2761 2893
rect 2797 2859 2831 2893
rect 2867 2859 2901 2893
rect 2937 2859 2971 2893
rect 3007 2859 3041 2893
rect 3077 2859 3111 2893
rect 3147 2859 3181 2893
rect 3217 2859 3251 2893
rect 3287 2859 3321 2893
rect 1677 2790 1711 2824
rect 1747 2790 1781 2824
rect 1817 2790 1851 2824
rect 1887 2790 1921 2824
rect 1957 2790 1991 2824
rect 2027 2790 2061 2824
rect 2097 2790 2131 2824
rect 2167 2790 2201 2824
rect 2237 2790 2271 2824
rect 2307 2790 2341 2824
rect 2377 2790 2411 2824
rect 2447 2790 2481 2824
rect 2517 2790 2551 2824
rect 2587 2790 2621 2824
rect 2657 2790 2691 2824
rect 2727 2790 2761 2824
rect 2797 2790 2831 2824
rect 2867 2790 2901 2824
rect 2937 2790 2971 2824
rect 3007 2790 3041 2824
rect 3077 2790 3111 2824
rect 3147 2790 3181 2824
rect 3217 2790 3251 2824
rect 3287 2790 3321 2824
rect 1677 2721 1711 2755
rect 1747 2721 1781 2755
rect 1817 2721 1851 2755
rect 1887 2721 1921 2755
rect 1957 2721 1991 2755
rect 2027 2721 2061 2755
rect 2097 2721 2131 2755
rect 2167 2721 2201 2755
rect 2237 2721 2271 2755
rect 2307 2721 2341 2755
rect 2377 2721 2411 2755
rect 2447 2721 2481 2755
rect 2517 2721 2551 2755
rect 2587 2721 2621 2755
rect 2657 2721 2691 2755
rect 2727 2721 2761 2755
rect 2797 2721 2831 2755
rect 2867 2721 2901 2755
rect 2937 2721 2971 2755
rect 3007 2721 3041 2755
rect 3077 2721 3111 2755
rect 3147 2721 3181 2755
rect 3217 2721 3251 2755
rect 3287 2721 3321 2755
rect 1677 2652 1711 2686
rect 1747 2652 1781 2686
rect 1817 2652 1851 2686
rect 1887 2652 1921 2686
rect 1957 2652 1991 2686
rect 2027 2652 2061 2686
rect 2097 2652 2131 2686
rect 2167 2652 2201 2686
rect 2237 2652 2271 2686
rect 2307 2652 2341 2686
rect 2377 2652 2411 2686
rect 2447 2652 2481 2686
rect 2517 2652 2551 2686
rect 2587 2652 2621 2686
rect 2657 2652 2691 2686
rect 2727 2652 2761 2686
rect 2797 2652 2831 2686
rect 2867 2652 2901 2686
rect 2937 2652 2971 2686
rect 3007 2652 3041 2686
rect 3077 2652 3111 2686
rect 3147 2652 3181 2686
rect 3217 2652 3251 2686
rect 3287 2652 3321 2686
rect 1677 2583 1711 2617
rect 1747 2583 1781 2617
rect 1817 2583 1851 2617
rect 1887 2583 1921 2617
rect 1957 2583 1991 2617
rect 2027 2583 2061 2617
rect 2097 2583 2131 2617
rect 2167 2583 2201 2617
rect 2237 2583 2271 2617
rect 2307 2583 2341 2617
rect 2377 2583 2411 2617
rect 2447 2583 2481 2617
rect 2517 2583 2551 2617
rect 2587 2583 2621 2617
rect 2657 2583 2691 2617
rect 2727 2583 2761 2617
rect 2797 2583 2831 2617
rect 2867 2583 2901 2617
rect 2937 2583 2971 2617
rect 3007 2583 3041 2617
rect 3077 2583 3111 2617
rect 3147 2583 3181 2617
rect 3217 2583 3251 2617
rect 3287 2583 3321 2617
rect 1677 2514 1711 2548
rect 1747 2514 1781 2548
rect 1817 2514 1851 2548
rect 1887 2514 1921 2548
rect 1957 2514 1991 2548
rect 2027 2514 2061 2548
rect 2097 2514 2131 2548
rect 2167 2514 2201 2548
rect 2237 2514 2271 2548
rect 2307 2514 2341 2548
rect 2377 2514 2411 2548
rect 2447 2514 2481 2548
rect 2517 2514 2551 2548
rect 2587 2514 2621 2548
rect 2657 2514 2691 2548
rect 2727 2514 2761 2548
rect 2797 2514 2831 2548
rect 2867 2514 2901 2548
rect 2937 2514 2971 2548
rect 3007 2514 3041 2548
rect 3077 2514 3111 2548
rect 3147 2514 3181 2548
rect 3217 2514 3251 2548
rect 3287 2514 3321 2548
rect 1677 2445 1711 2479
rect 1747 2445 1781 2479
rect 1817 2445 1851 2479
rect 1887 2445 1921 2479
rect 1957 2445 1991 2479
rect 2027 2445 2061 2479
rect 2097 2445 2131 2479
rect 2167 2445 2201 2479
rect 2237 2445 2271 2479
rect 2307 2445 2341 2479
rect 2377 2445 2411 2479
rect 2447 2445 2481 2479
rect 2517 2445 2551 2479
rect 2587 2445 2621 2479
rect 2657 2445 2691 2479
rect 2727 2445 2761 2479
rect 2797 2445 2831 2479
rect 2867 2445 2901 2479
rect 2937 2445 2971 2479
rect 3007 2445 3041 2479
rect 3077 2445 3111 2479
rect 3147 2445 3181 2479
rect 3217 2445 3251 2479
rect 3287 2445 3321 2479
rect 1677 2376 1711 2410
rect 1747 2376 1781 2410
rect 1817 2376 1851 2410
rect 1887 2376 1921 2410
rect 1957 2376 1991 2410
rect 2027 2376 2061 2410
rect 2097 2376 2131 2410
rect 2167 2376 2201 2410
rect 2237 2376 2271 2410
rect 2307 2376 2341 2410
rect 2377 2376 2411 2410
rect 2447 2376 2481 2410
rect 2517 2376 2551 2410
rect 2587 2376 2621 2410
rect 2657 2376 2691 2410
rect 2727 2376 2761 2410
rect 2797 2376 2831 2410
rect 2867 2376 2901 2410
rect 2937 2376 2971 2410
rect 3007 2376 3041 2410
rect 3077 2376 3111 2410
rect 3147 2376 3181 2410
rect 3217 2376 3251 2410
rect 3287 2376 3321 2410
rect 1677 2307 1711 2341
rect 1747 2307 1781 2341
rect 1817 2307 1851 2341
rect 1887 2307 1921 2341
rect 1957 2307 1991 2341
rect 2027 2307 2061 2341
rect 2097 2307 2131 2341
rect 2167 2307 2201 2341
rect 2237 2307 2271 2341
rect 2307 2307 2341 2341
rect 2377 2307 2411 2341
rect 2447 2307 2481 2341
rect 2517 2307 2551 2341
rect 2587 2307 2621 2341
rect 2657 2307 2691 2341
rect 2727 2307 2761 2341
rect 2797 2307 2831 2341
rect 2867 2307 2901 2341
rect 2937 2307 2971 2341
rect 3007 2307 3041 2341
rect 3077 2307 3111 2341
rect 3147 2307 3181 2341
rect 3217 2307 3251 2341
rect 3287 2307 3321 2341
rect 1677 2238 1711 2272
rect 1747 2238 1781 2272
rect 1817 2238 1851 2272
rect 1887 2238 1921 2272
rect 1957 2238 1991 2272
rect 2027 2238 2061 2272
rect 2097 2238 2131 2272
rect 2167 2238 2201 2272
rect 2237 2238 2271 2272
rect 2307 2238 2341 2272
rect 2377 2238 2411 2272
rect 2447 2238 2481 2272
rect 2517 2238 2551 2272
rect 2587 2238 2621 2272
rect 2657 2238 2691 2272
rect 2727 2238 2761 2272
rect 2797 2238 2831 2272
rect 2867 2238 2901 2272
rect 2937 2238 2971 2272
rect 3007 2238 3041 2272
rect 3077 2238 3111 2272
rect 3147 2238 3181 2272
rect 3217 2238 3251 2272
rect 3287 2238 3321 2272
rect 1677 2169 1711 2203
rect 1747 2169 1781 2203
rect 1817 2169 1851 2203
rect 1887 2169 1921 2203
rect 1957 2169 1991 2203
rect 2027 2169 2061 2203
rect 2097 2169 2131 2203
rect 2167 2169 2201 2203
rect 2237 2169 2271 2203
rect 2307 2169 2341 2203
rect 2377 2169 2411 2203
rect 2447 2169 2481 2203
rect 2517 2169 2551 2203
rect 2587 2169 2621 2203
rect 2657 2169 2691 2203
rect 2727 2169 2761 2203
rect 2797 2169 2831 2203
rect 2867 2169 2901 2203
rect 2937 2169 2971 2203
rect 3007 2169 3041 2203
rect 3077 2169 3111 2203
rect 3147 2169 3181 2203
rect 3217 2169 3251 2203
rect 3287 2169 3321 2203
rect 1677 2100 1711 2134
rect 1747 2100 1781 2134
rect 1817 2100 1851 2134
rect 1887 2100 1921 2134
rect 1957 2100 1991 2134
rect 2027 2100 2061 2134
rect 2097 2100 2131 2134
rect 2167 2100 2201 2134
rect 2237 2100 2271 2134
rect 2307 2100 2341 2134
rect 2377 2100 2411 2134
rect 2447 2100 2481 2134
rect 2517 2100 2551 2134
rect 2587 2100 2621 2134
rect 2657 2100 2691 2134
rect 2727 2100 2761 2134
rect 2797 2100 2831 2134
rect 2867 2100 2901 2134
rect 2937 2100 2971 2134
rect 3007 2100 3041 2134
rect 3077 2100 3111 2134
rect 3147 2100 3181 2134
rect 3217 2100 3251 2134
rect 3287 2100 3321 2134
rect 1677 2031 1711 2065
rect 1747 2031 1781 2065
rect 1817 2031 1851 2065
rect 1887 2031 1921 2065
rect 1957 2031 1991 2065
rect 2027 2031 2061 2065
rect 2097 2031 2131 2065
rect 2167 2031 2201 2065
rect 2237 2031 2271 2065
rect 2307 2031 2341 2065
rect 2377 2031 2411 2065
rect 2447 2031 2481 2065
rect 2517 2031 2551 2065
rect 2587 2031 2621 2065
rect 2657 2031 2691 2065
rect 2727 2031 2761 2065
rect 2797 2031 2831 2065
rect 2867 2031 2901 2065
rect 2937 2031 2971 2065
rect 3007 2031 3041 2065
rect 3077 2031 3111 2065
rect 3147 2031 3181 2065
rect 3217 2031 3251 2065
rect 3287 2031 3321 2065
rect 1677 1962 1711 1996
rect 1747 1962 1781 1996
rect 1817 1962 1851 1996
rect 1887 1962 1921 1996
rect 1957 1962 1991 1996
rect 2027 1962 2061 1996
rect 2097 1962 2131 1996
rect 2167 1962 2201 1996
rect 2237 1962 2271 1996
rect 2307 1962 2341 1996
rect 2377 1962 2411 1996
rect 2447 1962 2481 1996
rect 2517 1962 2551 1996
rect 2587 1962 2621 1996
rect 2657 1962 2691 1996
rect 2727 1962 2761 1996
rect 2797 1962 2831 1996
rect 2867 1962 2901 1996
rect 2937 1962 2971 1996
rect 3007 1962 3041 1996
rect 3077 1962 3111 1996
rect 3147 1962 3181 1996
rect 3217 1962 3251 1996
rect 3287 1962 3321 1996
rect 1677 1893 1711 1927
rect 1747 1893 1781 1927
rect 1817 1893 1851 1927
rect 1887 1893 1921 1927
rect 1957 1893 1991 1927
rect 2027 1893 2061 1927
rect 2097 1893 2131 1927
rect 2167 1893 2201 1927
rect 2237 1893 2271 1927
rect 2307 1893 2341 1927
rect 2377 1893 2411 1927
rect 2447 1893 2481 1927
rect 2517 1893 2551 1927
rect 2587 1893 2621 1927
rect 2657 1893 2691 1927
rect 2727 1893 2761 1927
rect 2797 1893 2831 1927
rect 2867 1893 2901 1927
rect 2937 1893 2971 1927
rect 3007 1893 3041 1927
rect 3077 1893 3111 1927
rect 3147 1893 3181 1927
rect 3217 1893 3251 1927
rect 3287 1893 3321 1927
rect 1677 1824 1711 1858
rect 1747 1824 1781 1858
rect 1817 1824 1851 1858
rect 1887 1824 1921 1858
rect 1957 1824 1991 1858
rect 2027 1824 2061 1858
rect 2097 1824 2131 1858
rect 2167 1824 2201 1858
rect 2237 1824 2271 1858
rect 2307 1824 2341 1858
rect 2377 1824 2411 1858
rect 2447 1824 2481 1858
rect 2517 1824 2551 1858
rect 2587 1824 2621 1858
rect 2657 1824 2691 1858
rect 2727 1824 2761 1858
rect 2797 1824 2831 1858
rect 2867 1824 2901 1858
rect 2937 1824 2971 1858
rect 3007 1824 3041 1858
rect 3077 1824 3111 1858
rect 3147 1824 3181 1858
rect 3217 1824 3251 1858
rect 3287 1824 3321 1858
rect 1677 1755 1711 1789
rect 1747 1755 1781 1789
rect 1817 1755 1851 1789
rect 1887 1755 1921 1789
rect 1957 1755 1991 1789
rect 2027 1755 2061 1789
rect 2097 1755 2131 1789
rect 2167 1755 2201 1789
rect 2237 1755 2271 1789
rect 2307 1755 2341 1789
rect 2377 1755 2411 1789
rect 2447 1755 2481 1789
rect 2517 1755 2551 1789
rect 2587 1755 2621 1789
rect 2657 1755 2691 1789
rect 2727 1755 2761 1789
rect 2797 1755 2831 1789
rect 2867 1755 2901 1789
rect 2937 1755 2971 1789
rect 3007 1755 3041 1789
rect 3077 1755 3111 1789
rect 3147 1755 3181 1789
rect 3217 1755 3251 1789
rect 3287 1755 3321 1789
rect 1677 1686 1711 1720
rect 1747 1686 1781 1720
rect 1817 1686 1851 1720
rect 1887 1686 1921 1720
rect 1957 1686 1991 1720
rect 2027 1686 2061 1720
rect 2097 1686 2131 1720
rect 2167 1686 2201 1720
rect 2237 1686 2271 1720
rect 2307 1686 2341 1720
rect 2377 1686 2411 1720
rect 2447 1686 2481 1720
rect 2517 1686 2551 1720
rect 2587 1686 2621 1720
rect 2657 1686 2691 1720
rect 2727 1686 2761 1720
rect 2797 1686 2831 1720
rect 2867 1686 2901 1720
rect 2937 1686 2971 1720
rect 3007 1686 3041 1720
rect 3077 1686 3111 1720
rect 3147 1686 3181 1720
rect 3217 1686 3251 1720
rect 3287 1686 3321 1720
rect 1677 1617 1711 1651
rect 1747 1617 1781 1651
rect 1817 1617 1851 1651
rect 1887 1617 1921 1651
rect 1957 1617 1991 1651
rect 2027 1617 2061 1651
rect 2097 1617 2131 1651
rect 2167 1617 2201 1651
rect 2237 1617 2271 1651
rect 2307 1617 2341 1651
rect 2377 1617 2411 1651
rect 2447 1617 2481 1651
rect 2517 1617 2551 1651
rect 2587 1617 2621 1651
rect 2657 1617 2691 1651
rect 2727 1617 2761 1651
rect 2797 1617 2831 1651
rect 2867 1617 2901 1651
rect 2937 1617 2971 1651
rect 3007 1617 3041 1651
rect 3077 1617 3111 1651
rect 3147 1617 3181 1651
rect 3217 1617 3251 1651
rect 3287 1617 3321 1651
rect 1677 1548 1711 1582
rect 1747 1548 1781 1582
rect 1817 1548 1851 1582
rect 1887 1548 1921 1582
rect 1957 1548 1991 1582
rect 2027 1548 2061 1582
rect 2097 1548 2131 1582
rect 2167 1548 2201 1582
rect 2237 1548 2271 1582
rect 2307 1548 2341 1582
rect 2377 1548 2411 1582
rect 2447 1548 2481 1582
rect 2517 1548 2551 1582
rect 2587 1548 2621 1582
rect 2657 1548 2691 1582
rect 2727 1548 2761 1582
rect 2797 1548 2831 1582
rect 2867 1548 2901 1582
rect 2937 1548 2971 1582
rect 3007 1548 3041 1582
rect 3077 1548 3111 1582
rect 3147 1548 3181 1582
rect 3217 1548 3251 1582
rect 3287 1548 3321 1582
rect 1677 1479 1711 1513
rect 1747 1479 1781 1513
rect 1817 1479 1851 1513
rect 1887 1479 1921 1513
rect 1957 1479 1991 1513
rect 2027 1479 2061 1513
rect 2097 1479 2131 1513
rect 2167 1479 2201 1513
rect 2237 1479 2271 1513
rect 2307 1479 2341 1513
rect 2377 1479 2411 1513
rect 2447 1479 2481 1513
rect 2517 1479 2551 1513
rect 2587 1479 2621 1513
rect 2657 1479 2691 1513
rect 2727 1479 2761 1513
rect 2797 1479 2831 1513
rect 2867 1479 2901 1513
rect 2937 1479 2971 1513
rect 3007 1479 3041 1513
rect 3077 1479 3111 1513
rect 3147 1479 3181 1513
rect 3217 1479 3251 1513
rect 3287 1479 3321 1513
rect 1677 1410 1711 1444
rect 1747 1410 1781 1444
rect 1817 1410 1851 1444
rect 1887 1410 1921 1444
rect 1957 1410 1991 1444
rect 2027 1410 2061 1444
rect 2097 1410 2131 1444
rect 2167 1410 2201 1444
rect 2237 1410 2271 1444
rect 2307 1410 2341 1444
rect 2377 1410 2411 1444
rect 2447 1410 2481 1444
rect 2517 1410 2551 1444
rect 2587 1410 2621 1444
rect 2657 1410 2691 1444
rect 2727 1410 2761 1444
rect 2797 1410 2831 1444
rect 2867 1410 2901 1444
rect 2937 1410 2971 1444
rect 3007 1410 3041 1444
rect 3077 1410 3111 1444
rect 3147 1410 3181 1444
rect 3217 1410 3251 1444
rect 3287 1410 3321 1444
rect 1677 1341 1711 1375
rect 1747 1341 1781 1375
rect 1817 1341 1851 1375
rect 1887 1341 1921 1375
rect 1957 1341 1991 1375
rect 2027 1341 2061 1375
rect 2097 1341 2131 1375
rect 2167 1341 2201 1375
rect 2237 1341 2271 1375
rect 2307 1341 2341 1375
rect 2377 1341 2411 1375
rect 2447 1341 2481 1375
rect 2517 1341 2551 1375
rect 2587 1341 2621 1375
rect 2657 1341 2691 1375
rect 2727 1341 2761 1375
rect 2797 1341 2831 1375
rect 2867 1341 2901 1375
rect 2937 1341 2971 1375
rect 3007 1341 3041 1375
rect 3077 1341 3111 1375
rect 3147 1341 3181 1375
rect 3217 1341 3251 1375
rect 3287 1341 3321 1375
rect 1677 1272 1711 1306
rect 1747 1272 1781 1306
rect 1817 1272 1851 1306
rect 1887 1272 1921 1306
rect 1957 1272 1991 1306
rect 2027 1272 2061 1306
rect 2097 1272 2131 1306
rect 2167 1272 2201 1306
rect 2237 1272 2271 1306
rect 2307 1272 2341 1306
rect 2377 1272 2411 1306
rect 2447 1272 2481 1306
rect 2517 1272 2551 1306
rect 2587 1272 2621 1306
rect 2657 1272 2691 1306
rect 2727 1272 2761 1306
rect 2797 1272 2831 1306
rect 2867 1272 2901 1306
rect 2937 1272 2971 1306
rect 3007 1272 3041 1306
rect 3077 1272 3111 1306
rect 3147 1272 3181 1306
rect 3217 1272 3251 1306
rect 3287 1272 3321 1306
rect 1677 1203 1711 1237
rect 1747 1203 1781 1237
rect 1817 1203 1851 1237
rect 1887 1203 1921 1237
rect 1957 1203 1991 1237
rect 2027 1203 2061 1237
rect 2097 1203 2131 1237
rect 2167 1203 2201 1237
rect 2237 1203 2271 1237
rect 2307 1203 2341 1237
rect 2377 1203 2411 1237
rect 2447 1203 2481 1237
rect 2517 1203 2551 1237
rect 2587 1203 2621 1237
rect 2657 1203 2691 1237
rect 2727 1203 2761 1237
rect 2797 1203 2831 1237
rect 2867 1203 2901 1237
rect 2937 1203 2971 1237
rect 3007 1203 3041 1237
rect 3077 1203 3111 1237
rect 3147 1203 3181 1237
rect 3217 1203 3251 1237
rect 3287 1203 3321 1237
rect 1677 1134 1711 1168
rect 1747 1134 1781 1168
rect 1817 1134 1851 1168
rect 1887 1134 1921 1168
rect 1957 1134 1991 1168
rect 2027 1134 2061 1168
rect 2097 1134 2131 1168
rect 2167 1134 2201 1168
rect 2237 1134 2271 1168
rect 2307 1134 2341 1168
rect 2377 1134 2411 1168
rect 2447 1134 2481 1168
rect 2517 1134 2551 1168
rect 2587 1134 2621 1168
rect 2657 1134 2691 1168
rect 2727 1134 2761 1168
rect 2797 1134 2831 1168
rect 2867 1134 2901 1168
rect 2937 1134 2971 1168
rect 3007 1134 3041 1168
rect 3077 1134 3111 1168
rect 3147 1134 3181 1168
rect 3217 1134 3251 1168
rect 3287 1134 3321 1168
rect 1677 1065 1711 1099
rect 1747 1065 1781 1099
rect 1817 1065 1851 1099
rect 1887 1065 1921 1099
rect 1957 1065 1991 1099
rect 2027 1065 2061 1099
rect 2097 1065 2131 1099
rect 2167 1065 2201 1099
rect 2237 1065 2271 1099
rect 2307 1065 2341 1099
rect 2377 1065 2411 1099
rect 2447 1065 2481 1099
rect 2517 1065 2551 1099
rect 2587 1065 2621 1099
rect 2657 1065 2691 1099
rect 2727 1065 2761 1099
rect 2797 1065 2831 1099
rect 2867 1065 2901 1099
rect 2937 1065 2971 1099
rect 3007 1065 3041 1099
rect 3077 1065 3111 1099
rect 3147 1065 3181 1099
rect 3217 1065 3251 1099
rect 3287 1065 3321 1099
rect 1677 996 1711 1030
rect 1747 996 1781 1030
rect 1817 996 1851 1030
rect 1887 996 1921 1030
rect 1957 996 1991 1030
rect 2027 996 2061 1030
rect 2097 996 2131 1030
rect 2167 996 2201 1030
rect 2237 996 2271 1030
rect 2307 996 2341 1030
rect 2377 996 2411 1030
rect 2447 996 2481 1030
rect 2517 996 2551 1030
rect 2587 996 2621 1030
rect 2657 996 2691 1030
rect 2727 996 2761 1030
rect 2797 996 2831 1030
rect 2867 996 2901 1030
rect 2937 996 2971 1030
rect 3007 996 3041 1030
rect 3077 996 3111 1030
rect 3147 996 3181 1030
rect 3217 996 3251 1030
rect 3287 996 3321 1030
rect 1677 927 1711 961
rect 1747 927 1781 961
rect 1817 927 1851 961
rect 1887 927 1921 961
rect 1957 927 1991 961
rect 2027 927 2061 961
rect 2097 927 2131 961
rect 2167 927 2201 961
rect 2237 927 2271 961
rect 2307 927 2341 961
rect 2377 927 2411 961
rect 2447 927 2481 961
rect 2517 927 2551 961
rect 2587 927 2621 961
rect 2657 927 2691 961
rect 2727 927 2761 961
rect 2797 927 2831 961
rect 2867 927 2901 961
rect 2937 927 2971 961
rect 3007 927 3041 961
rect 3077 927 3111 961
rect 3147 927 3181 961
rect 3217 927 3251 961
rect 3287 927 3321 961
rect 1677 858 1711 892
rect 1747 858 1781 892
rect 1817 858 1851 892
rect 1887 858 1921 892
rect 1957 858 1991 892
rect 2027 858 2061 892
rect 2097 858 2131 892
rect 2167 858 2201 892
rect 2237 858 2271 892
rect 2307 858 2341 892
rect 2377 858 2411 892
rect 2447 858 2481 892
rect 2517 858 2551 892
rect 2587 858 2621 892
rect 2657 858 2691 892
rect 2727 858 2761 892
rect 2797 858 2831 892
rect 2867 858 2901 892
rect 2937 858 2971 892
rect 3007 858 3041 892
rect 3077 858 3111 892
rect 3147 858 3181 892
rect 3217 858 3251 892
rect 3287 858 3321 892
rect 1677 789 1711 823
rect 1747 789 1781 823
rect 1817 789 1851 823
rect 1887 789 1921 823
rect 1957 789 1991 823
rect 2027 789 2061 823
rect 2097 789 2131 823
rect 2167 789 2201 823
rect 2237 789 2271 823
rect 2307 789 2341 823
rect 2377 789 2411 823
rect 2447 789 2481 823
rect 2517 789 2551 823
rect 2587 789 2621 823
rect 2657 789 2691 823
rect 2727 789 2761 823
rect 2797 789 2831 823
rect 2867 789 2901 823
rect 2937 789 2971 823
rect 3007 789 3041 823
rect 3077 789 3111 823
rect 3147 789 3181 823
rect 3217 789 3251 823
rect 3287 789 3321 823
rect 1677 720 1711 754
rect 1747 720 1781 754
rect 1817 720 1851 754
rect 1887 720 1921 754
rect 1957 720 1991 754
rect 2027 720 2061 754
rect 2097 720 2131 754
rect 2167 720 2201 754
rect 2237 720 2271 754
rect 2307 720 2341 754
rect 2377 720 2411 754
rect 2447 720 2481 754
rect 2517 720 2551 754
rect 2587 720 2621 754
rect 2657 720 2691 754
rect 2727 720 2761 754
rect 2797 720 2831 754
rect 2867 720 2901 754
rect 2937 720 2971 754
rect 3007 720 3041 754
rect 3077 720 3111 754
rect 3147 720 3181 754
rect 3217 720 3251 754
rect 3287 720 3321 754
rect 1677 651 1711 685
rect 1747 651 1781 685
rect 1817 651 1851 685
rect 1887 651 1921 685
rect 1957 651 1991 685
rect 2027 651 2061 685
rect 2097 651 2131 685
rect 2167 651 2201 685
rect 2237 651 2271 685
rect 2307 651 2341 685
rect 2377 651 2411 685
rect 2447 651 2481 685
rect 2517 651 2551 685
rect 2587 651 2621 685
rect 2657 651 2691 685
rect 2727 651 2761 685
rect 2797 651 2831 685
rect 2867 651 2901 685
rect 2937 651 2971 685
rect 3007 651 3041 685
rect 3077 651 3111 685
rect 3147 651 3181 685
rect 3217 651 3251 685
rect 3287 651 3321 685
rect 1677 582 1711 616
rect 1747 582 1781 616
rect 1817 582 1851 616
rect 1887 582 1921 616
rect 1957 582 1991 616
rect 2027 582 2061 616
rect 2097 582 2131 616
rect 2167 582 2201 616
rect 2237 582 2271 616
rect 2307 582 2341 616
rect 2377 582 2411 616
rect 2447 582 2481 616
rect 2517 582 2551 616
rect 2587 582 2621 616
rect 2657 582 2691 616
rect 2727 582 2761 616
rect 2797 582 2831 616
rect 2867 582 2901 616
rect 2937 582 2971 616
rect 3007 582 3041 616
rect 3077 582 3111 616
rect 3147 582 3181 616
rect 3217 582 3251 616
rect 3287 582 3321 616
rect 1677 513 1711 547
rect 1747 513 1781 547
rect 1817 513 1851 547
rect 1887 513 1921 547
rect 1957 513 1991 547
rect 2027 513 2061 547
rect 2097 513 2131 547
rect 2167 513 2201 547
rect 2237 513 2271 547
rect 2307 513 2341 547
rect 2377 513 2411 547
rect 2447 513 2481 547
rect 2517 513 2551 547
rect 2587 513 2621 547
rect 2657 513 2691 547
rect 2727 513 2761 547
rect 2797 513 2831 547
rect 2867 513 2901 547
rect 2937 513 2971 547
rect 3007 513 3041 547
rect 3077 513 3111 547
rect 3147 513 3181 547
rect 3217 513 3251 547
rect 3287 513 3321 547
rect 1677 444 1711 478
rect 1747 444 1781 478
rect 1817 444 1851 478
rect 1887 444 1921 478
rect 1957 444 1991 478
rect 2027 444 2061 478
rect 2097 444 2131 478
rect 2167 444 2201 478
rect 2237 444 2271 478
rect 2307 444 2341 478
rect 2377 444 2411 478
rect 2447 444 2481 478
rect 2517 444 2551 478
rect 2587 444 2621 478
rect 2657 444 2691 478
rect 2727 444 2761 478
rect 2797 444 2831 478
rect 2867 444 2901 478
rect 2937 444 2971 478
rect 3007 444 3041 478
rect 3077 444 3111 478
rect 3147 444 3181 478
rect 3217 444 3251 478
rect 3287 444 3321 478
rect 1677 375 1711 409
rect 1747 375 1781 409
rect 1817 375 1851 409
rect 1887 375 1921 409
rect 1957 375 1991 409
rect 2027 375 2061 409
rect 2097 375 2131 409
rect 2167 375 2201 409
rect 2237 375 2271 409
rect 2307 375 2341 409
rect 2377 375 2411 409
rect 2447 375 2481 409
rect 2517 375 2551 409
rect 2587 375 2621 409
rect 2657 375 2691 409
rect 2727 375 2761 409
rect 2797 375 2831 409
rect 2867 375 2901 409
rect 2937 375 2971 409
rect 3007 375 3041 409
rect 3077 375 3111 409
rect 3147 375 3181 409
rect 3217 375 3251 409
rect 3287 375 3321 409
rect 1677 306 1711 340
rect 1747 306 1781 340
rect 1817 306 1851 340
rect 1887 306 1921 340
rect 1957 306 1991 340
rect 2027 306 2061 340
rect 2097 306 2131 340
rect 2167 306 2201 340
rect 2237 306 2271 340
rect 2307 306 2341 340
rect 2377 306 2411 340
rect 2447 306 2481 340
rect 2517 306 2551 340
rect 2587 306 2621 340
rect 2657 306 2691 340
rect 2727 306 2761 340
rect 2797 306 2831 340
rect 2867 306 2901 340
rect 2937 306 2971 340
rect 3007 306 3041 340
rect 3077 306 3111 340
rect 3147 306 3181 340
rect 3217 306 3251 340
rect 3287 306 3321 340
<< nsubdiffcont >>
rect 368 3408 402 3442
rect 436 3408 470 3442
rect 504 3408 538 3442
rect 572 3408 606 3442
rect 640 3408 674 3442
rect 708 3408 742 3442
rect 776 3408 810 3442
rect 844 3408 878 3442
rect 912 3408 946 3442
rect 980 3408 1014 3442
rect 1048 3408 1082 3442
rect 1116 3408 1150 3442
rect 1184 3408 1218 3442
rect 1252 3408 1286 3442
rect 1320 3408 1354 3442
rect 270 3340 304 3374
rect 270 3272 304 3306
rect 270 3204 304 3238
rect 270 3136 304 3170
rect 270 3068 304 3102
rect 270 3000 304 3034
rect 270 2932 304 2966
rect 270 2864 304 2898
rect 270 2796 304 2830
rect 270 2728 304 2762
rect 270 2660 304 2694
rect 270 2592 304 2626
rect 270 2524 304 2558
rect 270 2456 304 2490
rect 270 2388 304 2422
rect 270 2320 304 2354
rect 270 2252 304 2286
rect 270 2184 304 2218
rect 270 2116 304 2150
rect 270 2048 304 2082
rect 270 1980 304 2014
rect 270 1912 304 1946
rect 1388 3332 1422 3366
rect 1388 3264 1422 3298
rect 1388 3196 1422 3230
rect 1388 3128 1422 3162
rect 1388 3060 1422 3094
rect 1388 2992 1422 3026
rect 1388 2924 1422 2958
rect 1388 2856 1422 2890
rect 1388 2788 1422 2822
rect 1388 2720 1422 2754
rect 1388 2652 1422 2686
rect 1388 2584 1422 2618
rect 1388 2516 1422 2550
rect 1388 2448 1422 2482
rect 1388 2380 1422 2414
rect 1388 2312 1422 2346
rect 1388 2244 1422 2278
rect 1388 2176 1422 2210
rect 1388 2108 1422 2142
rect 1388 2040 1422 2074
rect 1388 1972 1422 2006
rect 1388 1904 1422 1938
rect 270 1844 304 1878
rect 1388 1836 1422 1870
rect 270 1776 304 1810
rect 270 1708 304 1742
rect 270 1640 304 1674
rect 270 1572 304 1606
rect 270 1504 304 1538
rect 270 1436 304 1470
rect 270 1368 304 1402
rect 270 1300 304 1334
rect 270 1232 304 1266
rect 270 1164 304 1198
rect 270 1096 304 1130
rect 270 1028 304 1062
rect 270 960 304 994
rect 270 892 304 926
rect 270 824 304 858
rect 270 756 304 790
rect 270 688 304 722
rect 270 620 304 654
rect 270 552 304 586
rect 270 484 304 518
rect 270 416 304 450
rect 270 348 304 382
rect 1388 1768 1422 1802
rect 1388 1700 1422 1734
rect 1388 1632 1422 1666
rect 1388 1564 1422 1598
rect 1388 1496 1422 1530
rect 1388 1428 1422 1462
rect 1388 1360 1422 1394
rect 1388 1292 1422 1326
rect 1388 1224 1422 1258
rect 1388 1156 1422 1190
rect 1388 1088 1422 1122
rect 1388 1020 1422 1054
rect 1388 952 1422 986
rect 1388 884 1422 918
rect 1388 816 1422 850
rect 1388 748 1422 782
rect 1388 680 1422 714
rect 1388 612 1422 646
rect 1388 544 1422 578
rect 1388 476 1422 510
rect 1388 408 1422 442
rect 1388 340 1422 374
rect 1388 272 1422 306
rect 13621 3420 13655 3454
rect 13689 3420 13723 3454
rect 13757 3420 13791 3454
rect 13825 3420 13859 3454
rect 13893 3420 13927 3454
rect 13961 3420 13995 3454
rect 14029 3420 14063 3454
rect 14097 3420 14131 3454
rect 14165 3420 14199 3454
rect 14233 3420 14267 3454
rect 14301 3420 14335 3454
rect 14369 3420 14403 3454
rect 14437 3420 14471 3454
rect 14505 3420 14539 3454
rect 14573 3420 14607 3454
rect 13523 3352 13557 3386
rect 13523 3284 13557 3318
rect 13523 3216 13557 3250
rect 13523 3148 13557 3182
rect 13523 3080 13557 3114
rect 13523 3012 13557 3046
rect 13523 2944 13557 2978
rect 13523 2876 13557 2910
rect 13523 2808 13557 2842
rect 13523 2740 13557 2774
rect 13523 2672 13557 2706
rect 13523 2604 13557 2638
rect 13523 2536 13557 2570
rect 13523 2468 13557 2502
rect 13523 2400 13557 2434
rect 13523 2332 13557 2366
rect 13523 2264 13557 2298
rect 13523 2196 13557 2230
rect 13523 2128 13557 2162
rect 13523 2060 13557 2094
rect 13523 1992 13557 2026
rect 13523 1924 13557 1958
rect 14641 3344 14675 3378
rect 14641 3276 14675 3310
rect 14641 3208 14675 3242
rect 14641 3140 14675 3174
rect 14641 3072 14675 3106
rect 14641 3004 14675 3038
rect 14641 2936 14675 2970
rect 14641 2868 14675 2902
rect 14641 2800 14675 2834
rect 14641 2732 14675 2766
rect 14641 2664 14675 2698
rect 14641 2596 14675 2630
rect 14641 2528 14675 2562
rect 14641 2460 14675 2494
rect 14641 2392 14675 2426
rect 14641 2324 14675 2358
rect 14641 2256 14675 2290
rect 14641 2188 14675 2222
rect 14641 2120 14675 2154
rect 14641 2052 14675 2086
rect 14641 1984 14675 2018
rect 14641 1916 14675 1950
rect 13523 1856 13557 1890
rect 14641 1848 14675 1882
rect 13523 1788 13557 1822
rect 13523 1720 13557 1754
rect 13523 1652 13557 1686
rect 13523 1584 13557 1618
rect 13523 1516 13557 1550
rect 13523 1448 13557 1482
rect 13523 1380 13557 1414
rect 13523 1312 13557 1346
rect 13523 1244 13557 1278
rect 13523 1176 13557 1210
rect 13523 1108 13557 1142
rect 13523 1040 13557 1074
rect 13523 972 13557 1006
rect 13523 904 13557 938
rect 13523 836 13557 870
rect 13523 768 13557 802
rect 13523 700 13557 734
rect 13523 632 13557 666
rect 13523 564 13557 598
rect 13523 496 13557 530
rect 13523 428 13557 462
rect 13523 360 13557 394
rect 14641 1780 14675 1814
rect 14641 1712 14675 1746
rect 14641 1644 14675 1678
rect 14641 1576 14675 1610
rect 14641 1508 14675 1542
rect 14641 1440 14675 1474
rect 14641 1372 14675 1406
rect 14641 1304 14675 1338
rect 14641 1236 14675 1270
rect 14641 1168 14675 1202
rect 14641 1100 14675 1134
rect 14641 1032 14675 1066
rect 14641 964 14675 998
rect 14641 896 14675 930
rect 14641 828 14675 862
rect 14641 760 14675 794
rect 14641 692 14675 726
rect 14641 624 14675 658
rect 14641 556 14675 590
rect 14641 488 14675 522
rect 14641 420 14675 454
rect 338 204 372 238
rect 406 204 440 238
rect 474 204 508 238
rect 542 204 576 238
rect 610 204 644 238
rect 678 204 712 238
rect 746 204 780 238
rect 814 204 848 238
rect 882 204 916 238
rect 950 204 984 238
rect 1018 204 1052 238
rect 1086 204 1120 238
rect 1154 204 1188 238
rect 1222 204 1256 238
rect 1290 204 1324 238
rect 14641 352 14675 386
rect 14641 284 14675 318
rect 13591 216 13625 250
rect 13659 216 13693 250
rect 13727 216 13761 250
rect 13795 216 13829 250
rect 13863 216 13897 250
rect 13931 216 13965 250
rect 13999 216 14033 250
rect 14067 216 14101 250
rect 14135 216 14169 250
rect 14203 216 14237 250
rect 14271 216 14305 250
rect 14339 216 14373 250
rect 14407 216 14441 250
rect 14475 216 14509 250
rect 14543 216 14577 250
<< mvnsubdiffcont >>
rect 2076 39440 2110 39474
rect 1946 5508 2048 39406
rect 2144 39372 13874 39474
rect 13908 39321 13942 39355
rect 4382 19985 4416 20019
rect 4450 19985 4484 20019
rect 4518 19985 4552 20019
rect 4586 19985 4620 20019
rect 4654 19985 4688 20019
rect 4722 19985 4756 20019
rect 4790 19985 4824 20019
rect 4858 19985 4892 20019
rect 4926 19985 4960 20019
rect 4994 19985 5028 20019
rect 5062 19985 5096 20019
rect 5130 19985 5164 20019
rect 5198 19985 5232 20019
rect 5266 19985 5300 20019
rect 5334 19985 5368 20019
rect 5402 19985 5436 20019
rect 5470 19985 5504 20019
rect 5538 19985 5572 20019
rect 5606 19985 5640 20019
rect 5674 19985 5708 20019
rect 5742 19985 5776 20019
rect 5810 19985 5844 20019
rect 5878 19985 5912 20019
rect 5946 19985 5980 20019
rect 6014 19985 6048 20019
rect 6082 19985 6116 20019
rect 6150 19985 6184 20019
rect 6218 19985 6252 20019
rect 6286 19985 6320 20019
rect 6354 19985 6388 20019
rect 6422 19985 6456 20019
rect 6490 19985 6524 20019
rect 6558 19985 6592 20019
rect 6626 19985 6660 20019
rect 6694 19985 6728 20019
rect 6762 19985 6796 20019
rect 6830 19985 6864 20019
rect 6898 19985 6932 20019
rect 6966 19985 7000 20019
rect 7034 19985 7068 20019
rect 7102 19985 7136 20019
rect 7170 19985 7204 20019
rect 7238 19985 7272 20019
rect 7306 19985 7340 20019
rect 7374 19985 7408 20019
rect 7442 19985 7476 20019
rect 7510 19985 7544 20019
rect 7578 19985 7612 20019
rect 7646 19985 7680 20019
rect 7714 19985 7748 20019
rect 7782 19985 7816 20019
rect 7850 19985 7884 20019
rect 7918 19985 7952 20019
rect 7986 19985 8020 20019
rect 8054 19985 8088 20019
rect 8122 19985 8156 20019
rect 8190 19985 8224 20019
rect 8258 19985 8292 20019
rect 8326 19985 8360 20019
rect 8394 19985 8428 20019
rect 8462 19985 8496 20019
rect 8530 19985 8564 20019
rect 8598 19985 8632 20019
rect 8666 19985 8700 20019
rect 8734 19985 8768 20019
rect 8802 19985 8836 20019
rect 8870 19985 8904 20019
rect 8938 19985 8972 20019
rect 9006 19985 9040 20019
rect 9074 19985 9108 20019
rect 9142 19985 9176 20019
rect 9210 19985 9244 20019
rect 9278 19985 9312 20019
rect 9346 19985 9380 20019
rect 9414 19985 9448 20019
rect 9482 19985 9516 20019
rect 9550 19985 9584 20019
rect 9618 19985 9652 20019
rect 9686 19985 9720 20019
rect 9754 19985 9788 20019
rect 9822 19985 9856 20019
rect 9890 19985 9924 20019
rect 9958 19985 9992 20019
rect 10026 19985 10060 20019
rect 10094 19985 10128 20019
rect 10162 19985 10196 20019
rect 10230 19985 10264 20019
rect 10298 19985 10332 20019
rect 10366 19985 10400 20019
rect 10434 19985 10468 20019
rect 10502 19985 10536 20019
rect 10570 19985 10604 20019
rect 10638 19985 10672 20019
rect 10706 19985 10740 20019
rect 10774 19985 10808 20019
rect 10842 19985 10876 20019
rect 10910 19985 10944 20019
rect 10978 19985 11012 20019
rect 11046 19985 11080 20019
rect 11114 19985 11148 20019
rect 11182 19985 11216 20019
rect 11250 19985 11284 20019
rect 11318 19985 11352 20019
rect 11386 19985 11420 20019
rect 11454 19985 11488 20019
rect 11522 19985 11556 20019
rect 11590 19985 11624 20019
rect 11658 19985 11692 20019
rect 11726 19985 11760 20019
rect 11794 19985 11828 20019
rect 11862 19985 11896 20019
rect 11930 19985 11964 20019
rect 11998 19985 12032 20019
rect 12066 19985 12100 20019
rect 12134 19985 12168 20019
rect 12202 19985 12236 20019
rect 12270 19985 12304 20019
rect 12338 19985 12372 20019
rect 12406 19985 12440 20019
rect 12474 19985 12508 20019
rect 12542 19985 12576 20019
rect 12610 19985 12644 20019
rect 12678 19985 12712 20019
rect 12746 19985 12780 20019
rect 12814 19985 12848 20019
rect 12882 19985 12916 20019
rect 12950 19985 12984 20019
rect 13018 19985 13052 20019
rect 13086 19985 13120 20019
rect 13154 19985 13188 20019
rect 13222 19985 13256 20019
rect 13290 19985 13324 20019
rect 13358 19985 13392 20019
rect 13426 19985 13460 20019
rect 13494 19985 13528 20019
rect 13562 19985 13596 20019
rect 13630 19985 13664 20019
rect 4314 19860 4348 19894
rect 4314 19792 4348 19826
rect 4314 19724 4348 19758
rect 4314 19656 4348 19690
rect 4314 19588 4348 19622
rect 4314 19520 4348 19554
rect 4314 19452 4348 19486
rect 4314 19384 4348 19418
rect 4314 19316 4348 19350
rect 4314 19248 4348 19282
rect 4314 19180 4348 19214
rect 4314 19112 4348 19146
rect 4314 19044 4348 19078
rect 4314 18976 4348 19010
rect 4314 18908 4348 18942
rect 4314 18840 4348 18874
rect 4314 18772 4348 18806
rect 4314 18704 4348 18738
rect 4314 18636 4348 18670
rect 4314 18568 4348 18602
rect 4314 18500 4348 18534
rect 4314 18432 4348 18466
rect 4314 18364 4348 18398
rect 4314 18296 4348 18330
rect 4314 18228 4348 18262
rect 4314 18160 4348 18194
rect 4314 18092 4348 18126
rect 4314 18024 4348 18058
rect 4314 17956 4348 17990
rect 4314 17888 4348 17922
rect 4314 17820 4348 17854
rect 4314 17752 4348 17786
rect 4314 17684 4348 17718
rect 4314 17616 4348 17650
rect 4314 17548 4348 17582
rect 4314 17480 4348 17514
rect 4314 17412 4348 17446
rect 4314 17344 4348 17378
rect 4314 17276 4348 17310
rect 4314 17208 4348 17242
rect 4314 17140 4348 17174
rect 4314 17072 4348 17106
rect 4314 17004 4348 17038
rect 4314 16936 4348 16970
rect 4314 16868 4348 16902
rect 4314 16800 4348 16834
rect 4314 16732 4348 16766
rect 4314 16664 4348 16698
rect 2208 16596 2242 16630
rect 2276 16596 2310 16630
rect 2344 16596 2378 16630
rect 2412 16596 2446 16630
rect 2480 16596 2514 16630
rect 2548 16596 2582 16630
rect 2616 16596 2650 16630
rect 2684 16596 2718 16630
rect 2752 16596 2786 16630
rect 2820 16596 2854 16630
rect 2888 16596 2922 16630
rect 2956 16596 2990 16630
rect 3024 16596 3058 16630
rect 3092 16596 3126 16630
rect 3160 16596 3194 16630
rect 3228 16596 3262 16630
rect 3296 16596 3330 16630
rect 3364 16596 3398 16630
rect 3432 16596 3466 16630
rect 3500 16596 3534 16630
rect 3568 16596 3602 16630
rect 3636 16596 3670 16630
rect 3704 16596 3738 16630
rect 3772 16596 3806 16630
rect 3840 16596 3874 16630
rect 3908 16596 3942 16630
rect 3976 16596 4010 16630
rect 4044 16596 4078 16630
rect 4112 16596 4146 16630
rect 4180 16596 4214 16630
rect 1946 4835 2048 5345
rect 13840 5593 13942 39287
rect 2020 4767 2054 4801
rect 2088 4767 2598 4869
rect 2666 4767 13240 4869
rect 13340 4767 13782 4869
rect 13840 4835 13942 5481
rect 13816 4767 13850 4801
<< poly >>
rect 1668 39272 1734 39288
rect 1668 39238 1684 39272
rect 1718 39238 1734 39272
rect 1668 39204 1734 39238
rect 1668 39170 1684 39204
rect 1718 39170 1734 39204
rect 1668 39154 1734 39170
rect 2872 38854 13118 38870
rect 2872 38820 2888 38854
rect 2922 38820 2957 38854
rect 2991 38820 3026 38854
rect 3060 38820 3095 38854
rect 3129 38820 3164 38854
rect 3198 38820 3233 38854
rect 3267 38820 3302 38854
rect 3336 38820 3371 38854
rect 3405 38820 3440 38854
rect 3474 38820 3509 38854
rect 3543 38820 3578 38854
rect 3612 38820 3647 38854
rect 3681 38820 3716 38854
rect 3750 38820 3785 38854
rect 3819 38820 3854 38854
rect 3888 38820 3923 38854
rect 3957 38820 3992 38854
rect 4026 38820 4061 38854
rect 4095 38820 4130 38854
rect 4164 38820 4199 38854
rect 4233 38820 4268 38854
rect 4302 38820 4337 38854
rect 4371 38820 4406 38854
rect 4440 38820 4475 38854
rect 4509 38820 4544 38854
rect 4578 38820 4613 38854
rect 4647 38820 4682 38854
rect 4716 38820 4751 38854
rect 4785 38820 4820 38854
rect 4854 38820 4889 38854
rect 4923 38820 4958 38854
rect 4992 38820 5027 38854
rect 5061 38820 5096 38854
rect 5130 38820 5165 38854
rect 5199 38820 5234 38854
rect 5268 38820 5303 38854
rect 5337 38820 5372 38854
rect 5406 38820 5441 38854
rect 5475 38820 5510 38854
rect 5544 38820 5579 38854
rect 5613 38820 5648 38854
rect 5682 38820 5717 38854
rect 5751 38820 5786 38854
rect 5820 38820 5855 38854
rect 5889 38820 5924 38854
rect 5958 38820 5993 38854
rect 6027 38820 6062 38854
rect 6096 38820 6131 38854
rect 6165 38820 6200 38854
rect 6234 38820 6268 38854
rect 6302 38820 6336 38854
rect 6370 38820 6404 38854
rect 6438 38820 6472 38854
rect 6506 38820 6540 38854
rect 6574 38820 6608 38854
rect 6642 38820 6676 38854
rect 6710 38820 6744 38854
rect 6778 38820 6812 38854
rect 6846 38820 6880 38854
rect 6914 38820 6948 38854
rect 6982 38820 7016 38854
rect 7050 38820 7084 38854
rect 7118 38820 7152 38854
rect 7186 38820 7220 38854
rect 7254 38820 7288 38854
rect 7322 38820 7356 38854
rect 7390 38820 7424 38854
rect 7458 38820 7492 38854
rect 7526 38820 7560 38854
rect 7594 38820 7628 38854
rect 7662 38820 7696 38854
rect 7730 38820 7764 38854
rect 7798 38820 7832 38854
rect 7866 38820 7900 38854
rect 7934 38820 7968 38854
rect 8002 38820 8036 38854
rect 8070 38820 8104 38854
rect 8138 38820 8172 38854
rect 8206 38820 8240 38854
rect 8274 38820 8308 38854
rect 8342 38820 8376 38854
rect 8410 38820 8444 38854
rect 8478 38820 8512 38854
rect 8546 38820 8580 38854
rect 8614 38820 8648 38854
rect 8682 38820 8716 38854
rect 8750 38820 8784 38854
rect 8818 38820 8852 38854
rect 8886 38820 8920 38854
rect 8954 38820 8988 38854
rect 9022 38820 9056 38854
rect 9090 38820 9124 38854
rect 9158 38820 9192 38854
rect 9226 38820 9260 38854
rect 9294 38820 9328 38854
rect 9362 38820 9396 38854
rect 9430 38820 9464 38854
rect 9498 38820 9532 38854
rect 9566 38820 9600 38854
rect 9634 38820 9668 38854
rect 9702 38820 9736 38854
rect 9770 38820 9804 38854
rect 9838 38820 9872 38854
rect 9906 38820 9940 38854
rect 9974 38820 10008 38854
rect 10042 38820 10076 38854
rect 10110 38820 10144 38854
rect 10178 38820 10212 38854
rect 10246 38820 10280 38854
rect 10314 38820 10348 38854
rect 10382 38820 10416 38854
rect 10450 38820 10484 38854
rect 10518 38820 10552 38854
rect 10586 38820 10620 38854
rect 10654 38820 10688 38854
rect 10722 38820 10756 38854
rect 10790 38820 10824 38854
rect 10858 38820 10892 38854
rect 10926 38820 10960 38854
rect 10994 38820 11028 38854
rect 11062 38820 11096 38854
rect 11130 38820 11164 38854
rect 11198 38820 11232 38854
rect 11266 38820 11300 38854
rect 11334 38820 11368 38854
rect 11402 38820 11436 38854
rect 11470 38820 11504 38854
rect 11538 38820 11572 38854
rect 11606 38820 11640 38854
rect 11674 38820 11708 38854
rect 11742 38820 11776 38854
rect 11810 38820 11844 38854
rect 11878 38820 11912 38854
rect 11946 38820 11980 38854
rect 12014 38820 12048 38854
rect 12082 38820 12116 38854
rect 12150 38820 12184 38854
rect 12218 38820 12252 38854
rect 12286 38820 12320 38854
rect 12354 38820 12388 38854
rect 12422 38820 12456 38854
rect 12490 38820 12524 38854
rect 12558 38820 12592 38854
rect 12626 38820 12660 38854
rect 12694 38820 12728 38854
rect 12762 38820 12796 38854
rect 12830 38820 12864 38854
rect 12898 38820 12932 38854
rect 12966 38820 13000 38854
rect 13034 38820 13068 38854
rect 13102 38820 13118 38854
rect 2872 38804 13118 38820
rect 2872 37324 13118 37340
rect 2872 37290 2888 37324
rect 2922 37290 2957 37324
rect 2991 37290 3026 37324
rect 3060 37290 3095 37324
rect 3129 37290 3164 37324
rect 3198 37290 3233 37324
rect 3267 37290 3302 37324
rect 3336 37290 3371 37324
rect 3405 37290 3440 37324
rect 3474 37290 3509 37324
rect 3543 37290 3578 37324
rect 3612 37290 3647 37324
rect 3681 37290 3716 37324
rect 3750 37290 3785 37324
rect 3819 37290 3854 37324
rect 3888 37290 3923 37324
rect 3957 37290 3992 37324
rect 4026 37290 4061 37324
rect 4095 37290 4130 37324
rect 4164 37290 4199 37324
rect 4233 37290 4268 37324
rect 4302 37290 4337 37324
rect 4371 37290 4406 37324
rect 4440 37290 4475 37324
rect 4509 37290 4544 37324
rect 4578 37290 4613 37324
rect 4647 37290 4682 37324
rect 4716 37290 4751 37324
rect 4785 37290 4820 37324
rect 4854 37290 4889 37324
rect 4923 37290 4958 37324
rect 4992 37290 5027 37324
rect 5061 37290 5096 37324
rect 5130 37290 5165 37324
rect 5199 37290 5234 37324
rect 5268 37290 5303 37324
rect 5337 37290 5372 37324
rect 5406 37290 5441 37324
rect 5475 37290 5510 37324
rect 5544 37290 5579 37324
rect 5613 37290 5648 37324
rect 5682 37290 5717 37324
rect 5751 37290 5786 37324
rect 5820 37290 5855 37324
rect 5889 37290 5924 37324
rect 5958 37290 5993 37324
rect 6027 37290 6062 37324
rect 6096 37290 6131 37324
rect 6165 37290 6200 37324
rect 6234 37290 6268 37324
rect 6302 37290 6336 37324
rect 6370 37290 6404 37324
rect 6438 37290 6472 37324
rect 6506 37290 6540 37324
rect 6574 37290 6608 37324
rect 6642 37290 6676 37324
rect 6710 37290 6744 37324
rect 6778 37290 6812 37324
rect 6846 37290 6880 37324
rect 6914 37290 6948 37324
rect 6982 37290 7016 37324
rect 7050 37290 7084 37324
rect 7118 37290 7152 37324
rect 7186 37290 7220 37324
rect 7254 37290 7288 37324
rect 7322 37290 7356 37324
rect 7390 37290 7424 37324
rect 7458 37290 7492 37324
rect 7526 37290 7560 37324
rect 7594 37290 7628 37324
rect 7662 37290 7696 37324
rect 7730 37290 7764 37324
rect 7798 37290 7832 37324
rect 7866 37290 7900 37324
rect 7934 37290 7968 37324
rect 8002 37290 8036 37324
rect 8070 37290 8104 37324
rect 8138 37290 8172 37324
rect 8206 37290 8240 37324
rect 8274 37290 8308 37324
rect 8342 37290 8376 37324
rect 8410 37290 8444 37324
rect 8478 37290 8512 37324
rect 8546 37290 8580 37324
rect 8614 37290 8648 37324
rect 8682 37290 8716 37324
rect 8750 37290 8784 37324
rect 8818 37290 8852 37324
rect 8886 37290 8920 37324
rect 8954 37290 8988 37324
rect 9022 37290 9056 37324
rect 9090 37290 9124 37324
rect 9158 37290 9192 37324
rect 9226 37290 9260 37324
rect 9294 37290 9328 37324
rect 9362 37290 9396 37324
rect 9430 37290 9464 37324
rect 9498 37290 9532 37324
rect 9566 37290 9600 37324
rect 9634 37290 9668 37324
rect 9702 37290 9736 37324
rect 9770 37290 9804 37324
rect 9838 37290 9872 37324
rect 9906 37290 9940 37324
rect 9974 37290 10008 37324
rect 10042 37290 10076 37324
rect 10110 37290 10144 37324
rect 10178 37290 10212 37324
rect 10246 37290 10280 37324
rect 10314 37290 10348 37324
rect 10382 37290 10416 37324
rect 10450 37290 10484 37324
rect 10518 37290 10552 37324
rect 10586 37290 10620 37324
rect 10654 37290 10688 37324
rect 10722 37290 10756 37324
rect 10790 37290 10824 37324
rect 10858 37290 10892 37324
rect 10926 37290 10960 37324
rect 10994 37290 11028 37324
rect 11062 37290 11096 37324
rect 11130 37290 11164 37324
rect 11198 37290 11232 37324
rect 11266 37290 11300 37324
rect 11334 37290 11368 37324
rect 11402 37290 11436 37324
rect 11470 37290 11504 37324
rect 11538 37290 11572 37324
rect 11606 37290 11640 37324
rect 11674 37290 11708 37324
rect 11742 37290 11776 37324
rect 11810 37290 11844 37324
rect 11878 37290 11912 37324
rect 11946 37290 11980 37324
rect 12014 37290 12048 37324
rect 12082 37290 12116 37324
rect 12150 37290 12184 37324
rect 12218 37290 12252 37324
rect 12286 37290 12320 37324
rect 12354 37290 12388 37324
rect 12422 37290 12456 37324
rect 12490 37290 12524 37324
rect 12558 37290 12592 37324
rect 12626 37290 12660 37324
rect 12694 37290 12728 37324
rect 12762 37290 12796 37324
rect 12830 37290 12864 37324
rect 12898 37290 12932 37324
rect 12966 37290 13000 37324
rect 13034 37290 13068 37324
rect 13102 37290 13118 37324
rect 2872 37274 13118 37290
rect 3426 36870 3462 37274
rect 3664 36870 3700 37274
rect 3980 36870 4016 37274
rect 4218 36870 4254 37274
rect 4534 36870 4570 37274
rect 4772 36870 4808 37274
rect 5088 36870 5124 37274
rect 5326 36870 5362 37274
rect 5642 36870 5678 37274
rect 5880 36870 5916 37274
rect 6196 36870 6232 37274
rect 6434 36870 6470 37274
rect 6750 36870 6786 37274
rect 6988 36870 7024 37274
rect 7304 36870 7340 37274
rect 7542 36870 7578 37274
rect 7858 36870 7894 37274
rect 8096 36870 8132 37274
rect 8412 36870 8448 37274
rect 8650 36870 8686 37274
rect 8966 36870 9002 37274
rect 9204 36870 9240 37274
rect 9520 36870 9556 37274
rect 9758 36870 9794 37274
rect 10074 36870 10110 37274
rect 10312 36870 10348 37274
rect 10628 36870 10664 37274
rect 10866 36870 10902 37274
rect 11182 36870 11218 37274
rect 11420 36870 11456 37274
rect 11736 36870 11772 37274
rect 11974 36870 12010 37274
rect 12290 36870 12326 37274
rect 12528 36870 12564 37274
rect 12844 36870 12880 37274
rect 13082 36870 13118 37274
rect 2872 36854 13118 36870
rect 2872 36820 2888 36854
rect 2922 36820 2957 36854
rect 2991 36820 3026 36854
rect 3060 36820 3095 36854
rect 3129 36820 3164 36854
rect 3198 36820 3233 36854
rect 3267 36820 3302 36854
rect 3336 36820 3371 36854
rect 3405 36820 3440 36854
rect 3474 36820 3509 36854
rect 3543 36820 3578 36854
rect 3612 36820 3647 36854
rect 3681 36820 3716 36854
rect 3750 36820 3785 36854
rect 3819 36820 3854 36854
rect 3888 36820 3923 36854
rect 3957 36820 3992 36854
rect 4026 36820 4061 36854
rect 4095 36820 4130 36854
rect 4164 36820 4199 36854
rect 4233 36820 4268 36854
rect 4302 36820 4337 36854
rect 4371 36820 4406 36854
rect 4440 36820 4475 36854
rect 4509 36820 4544 36854
rect 4578 36820 4613 36854
rect 4647 36820 4682 36854
rect 4716 36820 4751 36854
rect 4785 36820 4820 36854
rect 4854 36820 4889 36854
rect 4923 36820 4958 36854
rect 4992 36820 5027 36854
rect 5061 36820 5096 36854
rect 5130 36820 5165 36854
rect 5199 36820 5234 36854
rect 5268 36820 5303 36854
rect 5337 36820 5372 36854
rect 5406 36820 5441 36854
rect 5475 36820 5510 36854
rect 5544 36820 5579 36854
rect 5613 36820 5648 36854
rect 5682 36820 5717 36854
rect 5751 36820 5786 36854
rect 5820 36820 5855 36854
rect 5889 36820 5924 36854
rect 5958 36820 5993 36854
rect 6027 36820 6062 36854
rect 6096 36820 6131 36854
rect 6165 36820 6200 36854
rect 6234 36820 6268 36854
rect 6302 36820 6336 36854
rect 6370 36820 6404 36854
rect 6438 36820 6472 36854
rect 6506 36820 6540 36854
rect 6574 36820 6608 36854
rect 6642 36820 6676 36854
rect 6710 36820 6744 36854
rect 6778 36820 6812 36854
rect 6846 36820 6880 36854
rect 6914 36820 6948 36854
rect 6982 36820 7016 36854
rect 7050 36820 7084 36854
rect 7118 36820 7152 36854
rect 7186 36820 7220 36854
rect 7254 36820 7288 36854
rect 7322 36820 7356 36854
rect 7390 36820 7424 36854
rect 7458 36820 7492 36854
rect 7526 36820 7560 36854
rect 7594 36820 7628 36854
rect 7662 36820 7696 36854
rect 7730 36820 7764 36854
rect 7798 36820 7832 36854
rect 7866 36820 7900 36854
rect 7934 36820 7968 36854
rect 8002 36820 8036 36854
rect 8070 36820 8104 36854
rect 8138 36820 8172 36854
rect 8206 36820 8240 36854
rect 8274 36820 8308 36854
rect 8342 36820 8376 36854
rect 8410 36820 8444 36854
rect 8478 36820 8512 36854
rect 8546 36820 8580 36854
rect 8614 36820 8648 36854
rect 8682 36820 8716 36854
rect 8750 36820 8784 36854
rect 8818 36820 8852 36854
rect 8886 36820 8920 36854
rect 8954 36820 8988 36854
rect 9022 36820 9056 36854
rect 9090 36820 9124 36854
rect 9158 36820 9192 36854
rect 9226 36820 9260 36854
rect 9294 36820 9328 36854
rect 9362 36820 9396 36854
rect 9430 36820 9464 36854
rect 9498 36820 9532 36854
rect 9566 36820 9600 36854
rect 9634 36820 9668 36854
rect 9702 36820 9736 36854
rect 9770 36820 9804 36854
rect 9838 36820 9872 36854
rect 9906 36820 9940 36854
rect 9974 36820 10008 36854
rect 10042 36820 10076 36854
rect 10110 36820 10144 36854
rect 10178 36820 10212 36854
rect 10246 36820 10280 36854
rect 10314 36820 10348 36854
rect 10382 36820 10416 36854
rect 10450 36820 10484 36854
rect 10518 36820 10552 36854
rect 10586 36820 10620 36854
rect 10654 36820 10688 36854
rect 10722 36820 10756 36854
rect 10790 36820 10824 36854
rect 10858 36820 10892 36854
rect 10926 36820 10960 36854
rect 10994 36820 11028 36854
rect 11062 36820 11096 36854
rect 11130 36820 11164 36854
rect 11198 36820 11232 36854
rect 11266 36820 11300 36854
rect 11334 36820 11368 36854
rect 11402 36820 11436 36854
rect 11470 36820 11504 36854
rect 11538 36820 11572 36854
rect 11606 36820 11640 36854
rect 11674 36820 11708 36854
rect 11742 36820 11776 36854
rect 11810 36820 11844 36854
rect 11878 36820 11912 36854
rect 11946 36820 11980 36854
rect 12014 36820 12048 36854
rect 12082 36820 12116 36854
rect 12150 36820 12184 36854
rect 12218 36820 12252 36854
rect 12286 36820 12320 36854
rect 12354 36820 12388 36854
rect 12422 36820 12456 36854
rect 12490 36820 12524 36854
rect 12558 36820 12592 36854
rect 12626 36820 12660 36854
rect 12694 36820 12728 36854
rect 12762 36820 12796 36854
rect 12830 36820 12864 36854
rect 12898 36820 12932 36854
rect 12966 36820 13000 36854
rect 13034 36820 13068 36854
rect 13102 36820 13118 36854
rect 2872 36804 13118 36820
rect 3426 36783 3462 36804
rect 3664 36783 3700 36804
rect 3980 36783 4016 36804
rect 4218 36783 4254 36804
rect 4534 36783 4570 36804
rect 4772 36783 4808 36804
rect 5088 36783 5124 36804
rect 5326 36783 5362 36804
rect 5642 36783 5678 36804
rect 5880 36783 5916 36804
rect 6196 36783 6232 36804
rect 6434 36783 6470 36804
rect 6750 36783 6786 36804
rect 6988 36783 7024 36804
rect 7304 36783 7340 36804
rect 7542 36783 7578 36804
rect 7858 36783 7894 36804
rect 8096 36783 8132 36804
rect 8412 36783 8448 36804
rect 8650 36783 8686 36804
rect 8966 36783 9002 36804
rect 9204 36783 9240 36804
rect 9520 36783 9556 36804
rect 9758 36783 9794 36804
rect 10074 36783 10110 36804
rect 10312 36783 10348 36804
rect 10628 36783 10664 36804
rect 10866 36783 10902 36804
rect 11182 36783 11218 36804
rect 11420 36783 11456 36804
rect 11736 36783 11772 36804
rect 11974 36783 12010 36804
rect 12290 36783 12326 36804
rect 12528 36783 12564 36804
rect 12844 36783 12880 36804
rect 13082 36783 13118 36804
rect 2872 35324 13118 35340
rect 2872 35290 2888 35324
rect 2922 35290 2957 35324
rect 2991 35290 3026 35324
rect 3060 35290 3095 35324
rect 3129 35290 3164 35324
rect 3198 35290 3233 35324
rect 3267 35290 3302 35324
rect 3336 35290 3371 35324
rect 3405 35290 3440 35324
rect 3474 35290 3509 35324
rect 3543 35290 3578 35324
rect 3612 35290 3647 35324
rect 3681 35290 3716 35324
rect 3750 35290 3785 35324
rect 3819 35290 3854 35324
rect 3888 35290 3923 35324
rect 3957 35290 3992 35324
rect 4026 35290 4061 35324
rect 4095 35290 4130 35324
rect 4164 35290 4199 35324
rect 4233 35290 4268 35324
rect 4302 35290 4337 35324
rect 4371 35290 4406 35324
rect 4440 35290 4475 35324
rect 4509 35290 4544 35324
rect 4578 35290 4613 35324
rect 4647 35290 4682 35324
rect 4716 35290 4751 35324
rect 4785 35290 4820 35324
rect 4854 35290 4889 35324
rect 4923 35290 4958 35324
rect 4992 35290 5027 35324
rect 5061 35290 5096 35324
rect 5130 35290 5165 35324
rect 5199 35290 5234 35324
rect 5268 35290 5303 35324
rect 5337 35290 5372 35324
rect 5406 35290 5441 35324
rect 5475 35290 5510 35324
rect 5544 35290 5579 35324
rect 5613 35290 5648 35324
rect 5682 35290 5717 35324
rect 5751 35290 5786 35324
rect 5820 35290 5855 35324
rect 5889 35290 5924 35324
rect 5958 35290 5993 35324
rect 6027 35290 6062 35324
rect 6096 35290 6131 35324
rect 6165 35290 6200 35324
rect 6234 35290 6268 35324
rect 6302 35290 6336 35324
rect 6370 35290 6404 35324
rect 6438 35290 6472 35324
rect 6506 35290 6540 35324
rect 6574 35290 6608 35324
rect 6642 35290 6676 35324
rect 6710 35290 6744 35324
rect 6778 35290 6812 35324
rect 6846 35290 6880 35324
rect 6914 35290 6948 35324
rect 6982 35290 7016 35324
rect 7050 35290 7084 35324
rect 7118 35290 7152 35324
rect 7186 35290 7220 35324
rect 7254 35290 7288 35324
rect 7322 35290 7356 35324
rect 7390 35290 7424 35324
rect 7458 35290 7492 35324
rect 7526 35290 7560 35324
rect 7594 35290 7628 35324
rect 7662 35290 7696 35324
rect 7730 35290 7764 35324
rect 7798 35290 7832 35324
rect 7866 35290 7900 35324
rect 7934 35290 7968 35324
rect 8002 35290 8036 35324
rect 8070 35290 8104 35324
rect 8138 35290 8172 35324
rect 8206 35290 8240 35324
rect 8274 35290 8308 35324
rect 8342 35290 8376 35324
rect 8410 35290 8444 35324
rect 8478 35290 8512 35324
rect 8546 35290 8580 35324
rect 8614 35290 8648 35324
rect 8682 35290 8716 35324
rect 8750 35290 8784 35324
rect 8818 35290 8852 35324
rect 8886 35290 8920 35324
rect 8954 35290 8988 35324
rect 9022 35290 9056 35324
rect 9090 35290 9124 35324
rect 9158 35290 9192 35324
rect 9226 35290 9260 35324
rect 9294 35290 9328 35324
rect 9362 35290 9396 35324
rect 9430 35290 9464 35324
rect 9498 35290 9532 35324
rect 9566 35290 9600 35324
rect 9634 35290 9668 35324
rect 9702 35290 9736 35324
rect 9770 35290 9804 35324
rect 9838 35290 9872 35324
rect 9906 35290 9940 35324
rect 9974 35290 10008 35324
rect 10042 35290 10076 35324
rect 10110 35290 10144 35324
rect 10178 35290 10212 35324
rect 10246 35290 10280 35324
rect 10314 35290 10348 35324
rect 10382 35290 10416 35324
rect 10450 35290 10484 35324
rect 10518 35290 10552 35324
rect 10586 35290 10620 35324
rect 10654 35290 10688 35324
rect 10722 35290 10756 35324
rect 10790 35290 10824 35324
rect 10858 35290 10892 35324
rect 10926 35290 10960 35324
rect 10994 35290 11028 35324
rect 11062 35290 11096 35324
rect 11130 35290 11164 35324
rect 11198 35290 11232 35324
rect 11266 35290 11300 35324
rect 11334 35290 11368 35324
rect 11402 35290 11436 35324
rect 11470 35290 11504 35324
rect 11538 35290 11572 35324
rect 11606 35290 11640 35324
rect 11674 35290 11708 35324
rect 11742 35290 11776 35324
rect 11810 35290 11844 35324
rect 11878 35290 11912 35324
rect 11946 35290 11980 35324
rect 12014 35290 12048 35324
rect 12082 35290 12116 35324
rect 12150 35290 12184 35324
rect 12218 35290 12252 35324
rect 12286 35290 12320 35324
rect 12354 35290 12388 35324
rect 12422 35290 12456 35324
rect 12490 35290 12524 35324
rect 12558 35290 12592 35324
rect 12626 35290 12660 35324
rect 12694 35290 12728 35324
rect 12762 35290 12796 35324
rect 12830 35290 12864 35324
rect 12898 35290 12932 35324
rect 12966 35290 13000 35324
rect 13034 35290 13068 35324
rect 13102 35290 13118 35324
rect 2872 35274 13118 35290
rect 3491 34870 3527 35274
rect 3761 34870 3797 35274
rect 4327 34870 4363 35274
rect 4597 34870 4633 35274
rect 5163 34870 5199 35274
rect 5433 34870 5469 35274
rect 5999 34870 6035 35274
rect 6269 34870 6305 35274
rect 6835 34870 6871 35274
rect 7105 34870 7141 35274
rect 7671 34870 7707 35274
rect 7941 34870 7977 35274
rect 8507 34870 8543 35274
rect 8777 34870 8813 35274
rect 9343 34870 9379 35274
rect 9613 34870 9649 35274
rect 10179 34870 10215 35274
rect 10449 34870 10485 35274
rect 11015 34870 11051 35274
rect 11285 34870 11321 35274
rect 11851 34870 11887 35274
rect 12121 34870 12157 35274
rect 12687 34870 12723 35274
rect 12957 34870 12993 35274
rect 3491 34854 12993 34870
rect 3491 34820 3507 34854
rect 3541 34820 3576 34854
rect 3610 34820 3645 34854
rect 3679 34820 3714 34854
rect 3748 34820 3783 34854
rect 3817 34820 3852 34854
rect 3886 34820 3921 34854
rect 3955 34820 3990 34854
rect 4024 34820 4059 34854
rect 4093 34820 4128 34854
rect 4162 34820 4197 34854
rect 4231 34820 4266 34854
rect 4300 34820 4335 34854
rect 4369 34820 4404 34854
rect 4438 34820 4473 34854
rect 4507 34820 4542 34854
rect 4576 34820 4611 34854
rect 4645 34820 4680 34854
rect 4714 34820 4749 34854
rect 4783 34820 4818 34854
rect 4852 34820 4887 34854
rect 4921 34820 4956 34854
rect 4990 34820 5025 34854
rect 5059 34820 5094 34854
rect 5128 34820 5163 34854
rect 5197 34820 5232 34854
rect 5266 34820 5301 34854
rect 5335 34820 5370 34854
rect 5404 34820 5439 34854
rect 5473 34820 5508 34854
rect 5542 34820 5577 34854
rect 5611 34820 5646 34854
rect 5680 34820 5715 34854
rect 5749 34820 5784 34854
rect 5818 34820 5853 34854
rect 5887 34820 5922 34854
rect 5956 34820 5991 34854
rect 6025 34820 6060 34854
rect 6094 34820 6129 34854
rect 6163 34820 6198 34854
rect 6232 34820 6267 34854
rect 6301 34820 6336 34854
rect 6370 34820 6405 34854
rect 6439 34820 6474 34854
rect 6508 34820 6543 34854
rect 6577 34820 6612 34854
rect 6646 34820 6681 34854
rect 6715 34820 6750 34854
rect 6784 34820 6819 34854
rect 6853 34820 6888 34854
rect 6922 34820 6957 34854
rect 6991 34820 7026 34854
rect 7060 34820 7095 34854
rect 7129 34820 7163 34854
rect 7197 34820 7231 34854
rect 7265 34820 7299 34854
rect 7333 34820 7367 34854
rect 7401 34820 7435 34854
rect 7469 34820 7503 34854
rect 7537 34820 7571 34854
rect 7605 34820 7639 34854
rect 7673 34820 7707 34854
rect 7741 34820 7775 34854
rect 7809 34820 7843 34854
rect 7877 34820 7911 34854
rect 7945 34820 7979 34854
rect 8013 34820 8047 34854
rect 8081 34820 8115 34854
rect 8149 34820 8183 34854
rect 8217 34820 8251 34854
rect 8285 34820 8319 34854
rect 8353 34820 8387 34854
rect 8421 34820 8455 34854
rect 8489 34820 8523 34854
rect 8557 34820 8591 34854
rect 8625 34820 8659 34854
rect 8693 34820 8727 34854
rect 8761 34820 8795 34854
rect 8829 34820 8863 34854
rect 8897 34820 8931 34854
rect 8965 34820 8999 34854
rect 9033 34820 9067 34854
rect 9101 34820 9135 34854
rect 9169 34820 9203 34854
rect 9237 34820 9271 34854
rect 9305 34820 9339 34854
rect 9373 34820 9407 34854
rect 9441 34820 9475 34854
rect 9509 34820 9543 34854
rect 9577 34820 9611 34854
rect 9645 34820 9679 34854
rect 9713 34820 9747 34854
rect 9781 34820 9815 34854
rect 9849 34820 9883 34854
rect 9917 34820 9951 34854
rect 9985 34820 10019 34854
rect 10053 34820 10087 34854
rect 10121 34820 10155 34854
rect 10189 34820 10223 34854
rect 10257 34820 10291 34854
rect 10325 34820 10359 34854
rect 10393 34820 10427 34854
rect 10461 34820 10495 34854
rect 10529 34820 10563 34854
rect 10597 34820 10631 34854
rect 10665 34820 10699 34854
rect 10733 34820 10767 34854
rect 10801 34820 10835 34854
rect 10869 34820 10903 34854
rect 10937 34820 10971 34854
rect 11005 34820 11039 34854
rect 11073 34820 11107 34854
rect 11141 34820 11175 34854
rect 11209 34820 11243 34854
rect 11277 34820 11311 34854
rect 11345 34820 11379 34854
rect 11413 34820 11447 34854
rect 11481 34820 11515 34854
rect 11549 34820 11583 34854
rect 11617 34820 11651 34854
rect 11685 34820 11719 34854
rect 11753 34820 11787 34854
rect 11821 34820 11855 34854
rect 11889 34820 11923 34854
rect 11957 34820 11991 34854
rect 12025 34820 12059 34854
rect 12093 34820 12127 34854
rect 12161 34820 12195 34854
rect 12229 34820 12263 34854
rect 12297 34820 12331 34854
rect 12365 34820 12399 34854
rect 12433 34820 12467 34854
rect 12501 34820 12535 34854
rect 12569 34820 12603 34854
rect 12637 34820 12671 34854
rect 12705 34820 12739 34854
rect 12773 34820 12807 34854
rect 12841 34820 12875 34854
rect 12909 34820 12943 34854
rect 12977 34820 12993 34854
rect 3491 34804 12993 34820
rect 3491 34797 3527 34804
rect 3761 34797 3797 34804
rect 4327 34797 4363 34804
rect 4597 34797 4633 34804
rect 5163 34797 5199 34804
rect 5433 34797 5469 34804
rect 5999 34797 6035 34804
rect 6269 34797 6305 34804
rect 6835 34797 6871 34804
rect 7105 34797 7141 34804
rect 7671 34797 7707 34804
rect 7941 34797 7977 34804
rect 8507 34797 8543 34804
rect 8777 34797 8813 34804
rect 9343 34797 9379 34804
rect 9613 34797 9649 34804
rect 10179 34797 10215 34804
rect 10449 34797 10485 34804
rect 11015 34797 11051 34804
rect 11285 34797 11321 34804
rect 11851 34797 11887 34804
rect 12121 34797 12157 34804
rect 12687 34797 12723 34804
rect 12957 34797 12993 34804
rect 3491 33340 3527 33363
rect 3761 33340 3797 33363
rect 4327 33340 4363 33363
rect 4597 33340 4633 33363
rect 5163 33340 5199 33363
rect 5433 33340 5469 33363
rect 5999 33340 6035 33363
rect 6269 33340 6305 33363
rect 6835 33340 6871 33363
rect 7105 33340 7141 33363
rect 7671 33340 7707 33363
rect 7941 33340 7977 33363
rect 8507 33340 8543 33363
rect 8777 33340 8813 33363
rect 9343 33340 9379 33363
rect 9613 33340 9649 33363
rect 10179 33340 10215 33363
rect 10449 33340 10485 33363
rect 11015 33340 11051 33363
rect 11285 33340 11321 33363
rect 11851 33340 11887 33363
rect 12121 33340 12157 33363
rect 12687 33340 12723 33363
rect 12957 33340 12993 33363
rect 3491 33324 12993 33340
rect 3491 33290 3507 33324
rect 3541 33290 3576 33324
rect 3610 33290 3645 33324
rect 3679 33290 3714 33324
rect 3748 33290 3783 33324
rect 3817 33290 3852 33324
rect 3886 33290 3921 33324
rect 3955 33290 3990 33324
rect 4024 33290 4059 33324
rect 4093 33290 4128 33324
rect 4162 33290 4197 33324
rect 4231 33290 4266 33324
rect 4300 33290 4335 33324
rect 4369 33290 4404 33324
rect 4438 33290 4473 33324
rect 4507 33290 4542 33324
rect 4576 33290 4611 33324
rect 4645 33290 4680 33324
rect 4714 33290 4749 33324
rect 4783 33290 4818 33324
rect 4852 33290 4887 33324
rect 4921 33290 4956 33324
rect 4990 33290 5025 33324
rect 5059 33290 5094 33324
rect 5128 33290 5163 33324
rect 5197 33290 5232 33324
rect 5266 33290 5301 33324
rect 5335 33290 5370 33324
rect 5404 33290 5439 33324
rect 5473 33290 5508 33324
rect 5542 33290 5577 33324
rect 5611 33290 5646 33324
rect 5680 33290 5715 33324
rect 5749 33290 5784 33324
rect 5818 33290 5853 33324
rect 5887 33290 5922 33324
rect 5956 33290 5991 33324
rect 6025 33290 6060 33324
rect 6094 33290 6129 33324
rect 6163 33290 6198 33324
rect 6232 33290 6267 33324
rect 6301 33290 6336 33324
rect 6370 33290 6405 33324
rect 6439 33290 6474 33324
rect 6508 33290 6543 33324
rect 6577 33290 6612 33324
rect 6646 33290 6681 33324
rect 6715 33290 6750 33324
rect 6784 33290 6819 33324
rect 6853 33290 6888 33324
rect 6922 33290 6957 33324
rect 6991 33290 7026 33324
rect 7060 33290 7095 33324
rect 7129 33290 7163 33324
rect 7197 33290 7231 33324
rect 7265 33290 7299 33324
rect 7333 33290 7367 33324
rect 7401 33290 7435 33324
rect 7469 33290 7503 33324
rect 7537 33290 7571 33324
rect 7605 33290 7639 33324
rect 7673 33290 7707 33324
rect 7741 33290 7775 33324
rect 7809 33290 7843 33324
rect 7877 33290 7911 33324
rect 7945 33290 7979 33324
rect 8013 33290 8047 33324
rect 8081 33290 8115 33324
rect 8149 33290 8183 33324
rect 8217 33290 8251 33324
rect 8285 33290 8319 33324
rect 8353 33290 8387 33324
rect 8421 33290 8455 33324
rect 8489 33290 8523 33324
rect 8557 33290 8591 33324
rect 8625 33290 8659 33324
rect 8693 33290 8727 33324
rect 8761 33290 8795 33324
rect 8829 33290 8863 33324
rect 8897 33290 8931 33324
rect 8965 33290 8999 33324
rect 9033 33290 9067 33324
rect 9101 33290 9135 33324
rect 9169 33290 9203 33324
rect 9237 33290 9271 33324
rect 9305 33290 9339 33324
rect 9373 33290 9407 33324
rect 9441 33290 9475 33324
rect 9509 33290 9543 33324
rect 9577 33290 9611 33324
rect 9645 33290 9679 33324
rect 9713 33290 9747 33324
rect 9781 33290 9815 33324
rect 9849 33290 9883 33324
rect 9917 33290 9951 33324
rect 9985 33290 10019 33324
rect 10053 33290 10087 33324
rect 10121 33290 10155 33324
rect 10189 33290 10223 33324
rect 10257 33290 10291 33324
rect 10325 33290 10359 33324
rect 10393 33290 10427 33324
rect 10461 33290 10495 33324
rect 10529 33290 10563 33324
rect 10597 33290 10631 33324
rect 10665 33290 10699 33324
rect 10733 33290 10767 33324
rect 10801 33290 10835 33324
rect 10869 33290 10903 33324
rect 10937 33290 10971 33324
rect 11005 33290 11039 33324
rect 11073 33290 11107 33324
rect 11141 33290 11175 33324
rect 11209 33290 11243 33324
rect 11277 33290 11311 33324
rect 11345 33290 11379 33324
rect 11413 33290 11447 33324
rect 11481 33290 11515 33324
rect 11549 33290 11583 33324
rect 11617 33290 11651 33324
rect 11685 33290 11719 33324
rect 11753 33290 11787 33324
rect 11821 33290 11855 33324
rect 11889 33290 11923 33324
rect 11957 33290 11991 33324
rect 12025 33290 12059 33324
rect 12093 33290 12127 33324
rect 12161 33290 12195 33324
rect 12229 33290 12263 33324
rect 12297 33290 12331 33324
rect 12365 33290 12399 33324
rect 12433 33290 12467 33324
rect 12501 33290 12535 33324
rect 12569 33290 12603 33324
rect 12637 33290 12671 33324
rect 12705 33290 12739 33324
rect 12773 33290 12807 33324
rect 12841 33290 12875 33324
rect 12909 33290 12943 33324
rect 12977 33290 12993 33324
rect 3491 33274 12993 33290
rect 3491 32870 3527 33274
rect 3761 32870 3797 33274
rect 4327 32870 4363 33274
rect 4597 32870 4633 33274
rect 5163 32870 5199 33274
rect 5433 32870 5469 33274
rect 5999 32870 6035 33274
rect 6269 32870 6305 33274
rect 6835 32870 6871 33274
rect 7105 32870 7141 33274
rect 7671 32870 7707 33274
rect 7941 32870 7977 33274
rect 8507 32870 8543 33274
rect 8777 32870 8813 33274
rect 9343 32870 9379 33274
rect 9613 32870 9649 33274
rect 10179 32870 10215 33274
rect 10449 32870 10485 33274
rect 11015 32870 11051 33274
rect 11285 32870 11321 33274
rect 11851 32870 11887 33274
rect 12121 32870 12157 33274
rect 12687 32870 12723 33274
rect 12957 32870 12993 33274
rect 3491 32854 12993 32870
rect 3491 32820 3507 32854
rect 3541 32820 3576 32854
rect 3610 32820 3645 32854
rect 3679 32820 3714 32854
rect 3748 32820 3783 32854
rect 3817 32820 3852 32854
rect 3886 32820 3921 32854
rect 3955 32820 3990 32854
rect 4024 32820 4059 32854
rect 4093 32820 4128 32854
rect 4162 32820 4197 32854
rect 4231 32820 4266 32854
rect 4300 32820 4335 32854
rect 4369 32820 4404 32854
rect 4438 32820 4473 32854
rect 4507 32820 4542 32854
rect 4576 32820 4611 32854
rect 4645 32820 4680 32854
rect 4714 32820 4749 32854
rect 4783 32820 4818 32854
rect 4852 32820 4887 32854
rect 4921 32820 4956 32854
rect 4990 32820 5025 32854
rect 5059 32820 5094 32854
rect 5128 32820 5163 32854
rect 5197 32820 5232 32854
rect 5266 32820 5301 32854
rect 5335 32820 5370 32854
rect 5404 32820 5439 32854
rect 5473 32820 5508 32854
rect 5542 32820 5577 32854
rect 5611 32820 5646 32854
rect 5680 32820 5715 32854
rect 5749 32820 5784 32854
rect 5818 32820 5853 32854
rect 5887 32820 5922 32854
rect 5956 32820 5991 32854
rect 6025 32820 6060 32854
rect 6094 32820 6129 32854
rect 6163 32820 6198 32854
rect 6232 32820 6267 32854
rect 6301 32820 6336 32854
rect 6370 32820 6405 32854
rect 6439 32820 6474 32854
rect 6508 32820 6543 32854
rect 6577 32820 6612 32854
rect 6646 32820 6681 32854
rect 6715 32820 6750 32854
rect 6784 32820 6819 32854
rect 6853 32820 6888 32854
rect 6922 32820 6957 32854
rect 6991 32820 7026 32854
rect 7060 32820 7095 32854
rect 7129 32820 7163 32854
rect 7197 32820 7231 32854
rect 7265 32820 7299 32854
rect 7333 32820 7367 32854
rect 7401 32820 7435 32854
rect 7469 32820 7503 32854
rect 7537 32820 7571 32854
rect 7605 32820 7639 32854
rect 7673 32820 7707 32854
rect 7741 32820 7775 32854
rect 7809 32820 7843 32854
rect 7877 32820 7911 32854
rect 7945 32820 7979 32854
rect 8013 32820 8047 32854
rect 8081 32820 8115 32854
rect 8149 32820 8183 32854
rect 8217 32820 8251 32854
rect 8285 32820 8319 32854
rect 8353 32820 8387 32854
rect 8421 32820 8455 32854
rect 8489 32820 8523 32854
rect 8557 32820 8591 32854
rect 8625 32820 8659 32854
rect 8693 32820 8727 32854
rect 8761 32820 8795 32854
rect 8829 32820 8863 32854
rect 8897 32820 8931 32854
rect 8965 32820 8999 32854
rect 9033 32820 9067 32854
rect 9101 32820 9135 32854
rect 9169 32820 9203 32854
rect 9237 32820 9271 32854
rect 9305 32820 9339 32854
rect 9373 32820 9407 32854
rect 9441 32820 9475 32854
rect 9509 32820 9543 32854
rect 9577 32820 9611 32854
rect 9645 32820 9679 32854
rect 9713 32820 9747 32854
rect 9781 32820 9815 32854
rect 9849 32820 9883 32854
rect 9917 32820 9951 32854
rect 9985 32820 10019 32854
rect 10053 32820 10087 32854
rect 10121 32820 10155 32854
rect 10189 32820 10223 32854
rect 10257 32820 10291 32854
rect 10325 32820 10359 32854
rect 10393 32820 10427 32854
rect 10461 32820 10495 32854
rect 10529 32820 10563 32854
rect 10597 32820 10631 32854
rect 10665 32820 10699 32854
rect 10733 32820 10767 32854
rect 10801 32820 10835 32854
rect 10869 32820 10903 32854
rect 10937 32820 10971 32854
rect 11005 32820 11039 32854
rect 11073 32820 11107 32854
rect 11141 32820 11175 32854
rect 11209 32820 11243 32854
rect 11277 32820 11311 32854
rect 11345 32820 11379 32854
rect 11413 32820 11447 32854
rect 11481 32820 11515 32854
rect 11549 32820 11583 32854
rect 11617 32820 11651 32854
rect 11685 32820 11719 32854
rect 11753 32820 11787 32854
rect 11821 32820 11855 32854
rect 11889 32820 11923 32854
rect 11957 32820 11991 32854
rect 12025 32820 12059 32854
rect 12093 32820 12127 32854
rect 12161 32820 12195 32854
rect 12229 32820 12263 32854
rect 12297 32820 12331 32854
rect 12365 32820 12399 32854
rect 12433 32820 12467 32854
rect 12501 32820 12535 32854
rect 12569 32820 12603 32854
rect 12637 32820 12671 32854
rect 12705 32820 12739 32854
rect 12773 32820 12807 32854
rect 12841 32820 12875 32854
rect 12909 32820 12943 32854
rect 12977 32820 12993 32854
rect 3491 32804 12993 32820
rect 3491 31324 12993 31340
rect 3491 31290 3507 31324
rect 3541 31290 3576 31324
rect 3610 31290 3645 31324
rect 3679 31290 3714 31324
rect 3748 31290 3783 31324
rect 3817 31290 3852 31324
rect 3886 31290 3921 31324
rect 3955 31290 3990 31324
rect 4024 31290 4059 31324
rect 4093 31290 4128 31324
rect 4162 31290 4197 31324
rect 4231 31290 4266 31324
rect 4300 31290 4335 31324
rect 4369 31290 4404 31324
rect 4438 31290 4473 31324
rect 4507 31290 4542 31324
rect 4576 31290 4611 31324
rect 4645 31290 4680 31324
rect 4714 31290 4749 31324
rect 4783 31290 4818 31324
rect 4852 31290 4887 31324
rect 4921 31290 4956 31324
rect 4990 31290 5025 31324
rect 5059 31290 5094 31324
rect 5128 31290 5163 31324
rect 5197 31290 5232 31324
rect 5266 31290 5301 31324
rect 5335 31290 5370 31324
rect 5404 31290 5439 31324
rect 5473 31290 5508 31324
rect 5542 31290 5577 31324
rect 5611 31290 5646 31324
rect 5680 31290 5715 31324
rect 5749 31290 5784 31324
rect 5818 31290 5853 31324
rect 5887 31290 5922 31324
rect 5956 31290 5991 31324
rect 6025 31290 6060 31324
rect 6094 31290 6129 31324
rect 6163 31290 6198 31324
rect 6232 31290 6267 31324
rect 6301 31290 6336 31324
rect 6370 31290 6405 31324
rect 6439 31290 6474 31324
rect 6508 31290 6543 31324
rect 6577 31290 6612 31324
rect 6646 31290 6681 31324
rect 6715 31290 6750 31324
rect 6784 31290 6819 31324
rect 6853 31290 6888 31324
rect 6922 31290 6957 31324
rect 6991 31290 7026 31324
rect 7060 31290 7095 31324
rect 7129 31290 7163 31324
rect 7197 31290 7231 31324
rect 7265 31290 7299 31324
rect 7333 31290 7367 31324
rect 7401 31290 7435 31324
rect 7469 31290 7503 31324
rect 7537 31290 7571 31324
rect 7605 31290 7639 31324
rect 7673 31290 7707 31324
rect 7741 31290 7775 31324
rect 7809 31290 7843 31324
rect 7877 31290 7911 31324
rect 7945 31290 7979 31324
rect 8013 31290 8047 31324
rect 8081 31290 8115 31324
rect 8149 31290 8183 31324
rect 8217 31290 8251 31324
rect 8285 31290 8319 31324
rect 8353 31290 8387 31324
rect 8421 31290 8455 31324
rect 8489 31290 8523 31324
rect 8557 31290 8591 31324
rect 8625 31290 8659 31324
rect 8693 31290 8727 31324
rect 8761 31290 8795 31324
rect 8829 31290 8863 31324
rect 8897 31290 8931 31324
rect 8965 31290 8999 31324
rect 9033 31290 9067 31324
rect 9101 31290 9135 31324
rect 9169 31290 9203 31324
rect 9237 31290 9271 31324
rect 9305 31290 9339 31324
rect 9373 31290 9407 31324
rect 9441 31290 9475 31324
rect 9509 31290 9543 31324
rect 9577 31290 9611 31324
rect 9645 31290 9679 31324
rect 9713 31290 9747 31324
rect 9781 31290 9815 31324
rect 9849 31290 9883 31324
rect 9917 31290 9951 31324
rect 9985 31290 10019 31324
rect 10053 31290 10087 31324
rect 10121 31290 10155 31324
rect 10189 31290 10223 31324
rect 10257 31290 10291 31324
rect 10325 31290 10359 31324
rect 10393 31290 10427 31324
rect 10461 31290 10495 31324
rect 10529 31290 10563 31324
rect 10597 31290 10631 31324
rect 10665 31290 10699 31324
rect 10733 31290 10767 31324
rect 10801 31290 10835 31324
rect 10869 31290 10903 31324
rect 10937 31290 10971 31324
rect 11005 31290 11039 31324
rect 11073 31290 11107 31324
rect 11141 31290 11175 31324
rect 11209 31290 11243 31324
rect 11277 31290 11311 31324
rect 11345 31290 11379 31324
rect 11413 31290 11447 31324
rect 11481 31290 11515 31324
rect 11549 31290 11583 31324
rect 11617 31290 11651 31324
rect 11685 31290 11719 31324
rect 11753 31290 11787 31324
rect 11821 31290 11855 31324
rect 11889 31290 11923 31324
rect 11957 31290 11991 31324
rect 12025 31290 12059 31324
rect 12093 31290 12127 31324
rect 12161 31290 12195 31324
rect 12229 31290 12263 31324
rect 12297 31290 12331 31324
rect 12365 31290 12399 31324
rect 12433 31290 12467 31324
rect 12501 31290 12535 31324
rect 12569 31290 12603 31324
rect 12637 31290 12671 31324
rect 12705 31290 12739 31324
rect 12773 31290 12807 31324
rect 12841 31290 12875 31324
rect 12909 31290 12943 31324
rect 12977 31290 12993 31324
rect 3491 31274 12993 31290
rect 3491 30870 3527 31274
rect 3761 30870 3797 31274
rect 4327 30870 4363 31274
rect 4597 30870 4633 31274
rect 5163 30870 5199 31274
rect 5433 30870 5469 31274
rect 5999 30870 6035 31274
rect 6269 30870 6305 31274
rect 6835 30870 6871 31274
rect 7105 30870 7141 31274
rect 7671 30870 7707 31274
rect 7941 30870 7977 31274
rect 8507 30870 8543 31274
rect 8777 30870 8813 31274
rect 9343 30870 9379 31274
rect 9613 30870 9649 31274
rect 10179 30870 10215 31274
rect 10449 30870 10485 31274
rect 11015 30870 11051 31274
rect 11285 30870 11321 31274
rect 11851 30870 11887 31274
rect 12121 30870 12157 31274
rect 12687 30870 12723 31274
rect 12957 30870 12993 31274
rect 3491 30854 12993 30870
rect 3491 30820 3507 30854
rect 3541 30820 3576 30854
rect 3610 30820 3645 30854
rect 3679 30820 3714 30854
rect 3748 30820 3783 30854
rect 3817 30820 3852 30854
rect 3886 30820 3921 30854
rect 3955 30820 3990 30854
rect 4024 30820 4059 30854
rect 4093 30820 4128 30854
rect 4162 30820 4197 30854
rect 4231 30820 4266 30854
rect 4300 30820 4335 30854
rect 4369 30820 4404 30854
rect 4438 30820 4473 30854
rect 4507 30820 4542 30854
rect 4576 30820 4611 30854
rect 4645 30820 4680 30854
rect 4714 30820 4749 30854
rect 4783 30820 4818 30854
rect 4852 30820 4887 30854
rect 4921 30820 4956 30854
rect 4990 30820 5025 30854
rect 5059 30820 5094 30854
rect 5128 30820 5163 30854
rect 5197 30820 5232 30854
rect 5266 30820 5301 30854
rect 5335 30820 5370 30854
rect 5404 30820 5439 30854
rect 5473 30820 5508 30854
rect 5542 30820 5577 30854
rect 5611 30820 5646 30854
rect 5680 30820 5715 30854
rect 5749 30820 5784 30854
rect 5818 30820 5853 30854
rect 5887 30820 5922 30854
rect 5956 30820 5991 30854
rect 6025 30820 6060 30854
rect 6094 30820 6129 30854
rect 6163 30820 6198 30854
rect 6232 30820 6267 30854
rect 6301 30820 6336 30854
rect 6370 30820 6405 30854
rect 6439 30820 6474 30854
rect 6508 30820 6543 30854
rect 6577 30820 6612 30854
rect 6646 30820 6681 30854
rect 6715 30820 6750 30854
rect 6784 30820 6819 30854
rect 6853 30820 6888 30854
rect 6922 30820 6957 30854
rect 6991 30820 7026 30854
rect 7060 30820 7095 30854
rect 7129 30820 7163 30854
rect 7197 30820 7231 30854
rect 7265 30820 7299 30854
rect 7333 30820 7367 30854
rect 7401 30820 7435 30854
rect 7469 30820 7503 30854
rect 7537 30820 7571 30854
rect 7605 30820 7639 30854
rect 7673 30820 7707 30854
rect 7741 30820 7775 30854
rect 7809 30820 7843 30854
rect 7877 30820 7911 30854
rect 7945 30820 7979 30854
rect 8013 30820 8047 30854
rect 8081 30820 8115 30854
rect 8149 30820 8183 30854
rect 8217 30820 8251 30854
rect 8285 30820 8319 30854
rect 8353 30820 8387 30854
rect 8421 30820 8455 30854
rect 8489 30820 8523 30854
rect 8557 30820 8591 30854
rect 8625 30820 8659 30854
rect 8693 30820 8727 30854
rect 8761 30820 8795 30854
rect 8829 30820 8863 30854
rect 8897 30820 8931 30854
rect 8965 30820 8999 30854
rect 9033 30820 9067 30854
rect 9101 30820 9135 30854
rect 9169 30820 9203 30854
rect 9237 30820 9271 30854
rect 9305 30820 9339 30854
rect 9373 30820 9407 30854
rect 9441 30820 9475 30854
rect 9509 30820 9543 30854
rect 9577 30820 9611 30854
rect 9645 30820 9679 30854
rect 9713 30820 9747 30854
rect 9781 30820 9815 30854
rect 9849 30820 9883 30854
rect 9917 30820 9951 30854
rect 9985 30820 10019 30854
rect 10053 30820 10087 30854
rect 10121 30820 10155 30854
rect 10189 30820 10223 30854
rect 10257 30820 10291 30854
rect 10325 30820 10359 30854
rect 10393 30820 10427 30854
rect 10461 30820 10495 30854
rect 10529 30820 10563 30854
rect 10597 30820 10631 30854
rect 10665 30820 10699 30854
rect 10733 30820 10767 30854
rect 10801 30820 10835 30854
rect 10869 30820 10903 30854
rect 10937 30820 10971 30854
rect 11005 30820 11039 30854
rect 11073 30820 11107 30854
rect 11141 30820 11175 30854
rect 11209 30820 11243 30854
rect 11277 30820 11311 30854
rect 11345 30820 11379 30854
rect 11413 30820 11447 30854
rect 11481 30820 11515 30854
rect 11549 30820 11583 30854
rect 11617 30820 11651 30854
rect 11685 30820 11719 30854
rect 11753 30820 11787 30854
rect 11821 30820 11855 30854
rect 11889 30820 11923 30854
rect 11957 30820 11991 30854
rect 12025 30820 12059 30854
rect 12093 30820 12127 30854
rect 12161 30820 12195 30854
rect 12229 30820 12263 30854
rect 12297 30820 12331 30854
rect 12365 30820 12399 30854
rect 12433 30820 12467 30854
rect 12501 30820 12535 30854
rect 12569 30820 12603 30854
rect 12637 30820 12671 30854
rect 12705 30820 12739 30854
rect 12773 30820 12807 30854
rect 12841 30820 12875 30854
rect 12909 30820 12943 30854
rect 12977 30820 12993 30854
rect 3491 30804 12993 30820
rect 3491 30775 3527 30804
rect 3761 30775 3797 30804
rect 4327 30775 4363 30804
rect 4597 30775 4633 30804
rect 5163 30775 5199 30804
rect 5433 30775 5469 30804
rect 5999 30775 6035 30804
rect 6269 30775 6305 30804
rect 6835 30775 6871 30804
rect 7105 30775 7141 30804
rect 7671 30775 7707 30804
rect 7941 30775 7977 30804
rect 8507 30775 8543 30804
rect 8777 30775 8813 30804
rect 9343 30775 9379 30804
rect 9613 30775 9649 30804
rect 10179 30775 10215 30804
rect 10449 30775 10485 30804
rect 11015 30775 11051 30804
rect 11285 30775 11321 30804
rect 11851 30775 11887 30804
rect 12121 30775 12157 30804
rect 12687 30775 12723 30804
rect 12957 30775 12993 30804
rect 5163 29340 5199 29387
rect 5433 29340 5469 29387
rect 5999 29340 6035 29387
rect 6269 29340 6305 29387
rect 6835 29340 6871 29387
rect 7105 29340 7141 29387
rect 7671 29340 7707 29387
rect 7941 29340 7977 29387
rect 8507 29340 8543 29387
rect 8777 29340 8813 29387
rect 9343 29340 9379 29387
rect 9613 29340 9649 29387
rect 10179 29340 10215 29387
rect 10449 29340 10485 29387
rect 11015 29340 11051 29387
rect 11285 29340 11321 29387
rect 11851 29340 11887 29387
rect 12121 29340 12157 29387
rect 12687 29340 12723 29387
rect 12957 29340 12993 29387
rect 3491 29324 12993 29340
rect 3491 29290 3507 29324
rect 3541 29290 3576 29324
rect 3610 29290 3645 29324
rect 3679 29290 3714 29324
rect 3748 29290 3783 29324
rect 3817 29290 3852 29324
rect 3886 29290 3921 29324
rect 3955 29290 3990 29324
rect 4024 29290 4059 29324
rect 4093 29290 4128 29324
rect 4162 29290 4197 29324
rect 4231 29290 4266 29324
rect 4300 29290 4335 29324
rect 4369 29290 4404 29324
rect 4438 29290 4473 29324
rect 4507 29290 4542 29324
rect 4576 29290 4611 29324
rect 4645 29290 4680 29324
rect 4714 29290 4749 29324
rect 4783 29290 4818 29324
rect 4852 29290 4887 29324
rect 4921 29290 4956 29324
rect 4990 29290 5025 29324
rect 5059 29290 5094 29324
rect 5128 29290 5163 29324
rect 5197 29290 5232 29324
rect 5266 29290 5301 29324
rect 5335 29290 5370 29324
rect 5404 29290 5439 29324
rect 5473 29290 5508 29324
rect 5542 29290 5577 29324
rect 5611 29290 5646 29324
rect 5680 29290 5715 29324
rect 5749 29290 5784 29324
rect 5818 29290 5853 29324
rect 5887 29290 5922 29324
rect 5956 29290 5991 29324
rect 6025 29290 6060 29324
rect 6094 29290 6129 29324
rect 6163 29290 6198 29324
rect 6232 29290 6267 29324
rect 6301 29290 6336 29324
rect 6370 29290 6405 29324
rect 6439 29290 6474 29324
rect 6508 29290 6543 29324
rect 6577 29290 6612 29324
rect 6646 29290 6681 29324
rect 6715 29290 6750 29324
rect 6784 29290 6819 29324
rect 6853 29290 6888 29324
rect 6922 29290 6957 29324
rect 6991 29290 7026 29324
rect 7060 29290 7095 29324
rect 7129 29290 7163 29324
rect 7197 29290 7231 29324
rect 7265 29290 7299 29324
rect 7333 29290 7367 29324
rect 7401 29290 7435 29324
rect 7469 29290 7503 29324
rect 7537 29290 7571 29324
rect 7605 29290 7639 29324
rect 7673 29290 7707 29324
rect 7741 29290 7775 29324
rect 7809 29290 7843 29324
rect 7877 29290 7911 29324
rect 7945 29290 7979 29324
rect 8013 29290 8047 29324
rect 8081 29290 8115 29324
rect 8149 29290 8183 29324
rect 8217 29290 8251 29324
rect 8285 29290 8319 29324
rect 8353 29290 8387 29324
rect 8421 29290 8455 29324
rect 8489 29290 8523 29324
rect 8557 29290 8591 29324
rect 8625 29290 8659 29324
rect 8693 29290 8727 29324
rect 8761 29290 8795 29324
rect 8829 29290 8863 29324
rect 8897 29290 8931 29324
rect 8965 29290 8999 29324
rect 9033 29290 9067 29324
rect 9101 29290 9135 29324
rect 9169 29290 9203 29324
rect 9237 29290 9271 29324
rect 9305 29290 9339 29324
rect 9373 29290 9407 29324
rect 9441 29290 9475 29324
rect 9509 29290 9543 29324
rect 9577 29290 9611 29324
rect 9645 29290 9679 29324
rect 9713 29290 9747 29324
rect 9781 29290 9815 29324
rect 9849 29290 9883 29324
rect 9917 29290 9951 29324
rect 9985 29290 10019 29324
rect 10053 29290 10087 29324
rect 10121 29290 10155 29324
rect 10189 29290 10223 29324
rect 10257 29290 10291 29324
rect 10325 29290 10359 29324
rect 10393 29290 10427 29324
rect 10461 29290 10495 29324
rect 10529 29290 10563 29324
rect 10597 29290 10631 29324
rect 10665 29290 10699 29324
rect 10733 29290 10767 29324
rect 10801 29290 10835 29324
rect 10869 29290 10903 29324
rect 10937 29290 10971 29324
rect 11005 29290 11039 29324
rect 11073 29290 11107 29324
rect 11141 29290 11175 29324
rect 11209 29290 11243 29324
rect 11277 29290 11311 29324
rect 11345 29290 11379 29324
rect 11413 29290 11447 29324
rect 11481 29290 11515 29324
rect 11549 29290 11583 29324
rect 11617 29290 11651 29324
rect 11685 29290 11719 29324
rect 11753 29290 11787 29324
rect 11821 29290 11855 29324
rect 11889 29290 11923 29324
rect 11957 29290 11991 29324
rect 12025 29290 12059 29324
rect 12093 29290 12127 29324
rect 12161 29290 12195 29324
rect 12229 29290 12263 29324
rect 12297 29290 12331 29324
rect 12365 29290 12399 29324
rect 12433 29290 12467 29324
rect 12501 29290 12535 29324
rect 12569 29290 12603 29324
rect 12637 29290 12671 29324
rect 12705 29290 12739 29324
rect 12773 29290 12807 29324
rect 12841 29290 12875 29324
rect 12909 29290 12943 29324
rect 12977 29290 12993 29324
rect 3491 29274 12993 29290
rect 5163 28870 5199 29274
rect 5433 28870 5469 29274
rect 5999 28870 6035 29274
rect 6269 28870 6305 29274
rect 6835 28870 6871 29274
rect 7105 28870 7141 29274
rect 7671 28870 7707 29274
rect 7941 28870 7977 29274
rect 8507 28870 8543 29274
rect 8777 28870 8813 29274
rect 9343 28870 9379 29274
rect 9613 28870 9649 29274
rect 10179 28870 10215 29274
rect 10449 28870 10485 29274
rect 11015 28870 11051 29274
rect 11285 28870 11321 29274
rect 11851 28870 11887 29274
rect 12121 28870 12157 29274
rect 12687 28870 12723 29274
rect 12957 28870 12993 29274
rect 5163 28854 12993 28870
rect 5163 28820 5179 28854
rect 5213 28820 5248 28854
rect 5282 28820 5317 28854
rect 5351 28820 5386 28854
rect 5420 28820 5455 28854
rect 5489 28820 5524 28854
rect 5558 28820 5593 28854
rect 5627 28820 5662 28854
rect 5696 28820 5731 28854
rect 5765 28820 5800 28854
rect 5834 28820 5869 28854
rect 5903 28820 5938 28854
rect 5972 28820 6007 28854
rect 6041 28820 6075 28854
rect 6109 28820 6143 28854
rect 6177 28820 6211 28854
rect 6245 28820 6279 28854
rect 6313 28820 6347 28854
rect 6381 28820 6415 28854
rect 6449 28820 6483 28854
rect 6517 28820 6551 28854
rect 6585 28820 6619 28854
rect 6653 28820 6687 28854
rect 6721 28820 6755 28854
rect 6789 28820 6823 28854
rect 6857 28820 6891 28854
rect 6925 28820 6959 28854
rect 6993 28820 7027 28854
rect 7061 28820 7095 28854
rect 7129 28820 7163 28854
rect 7197 28820 7231 28854
rect 7265 28820 7299 28854
rect 7333 28820 7367 28854
rect 7401 28820 7435 28854
rect 7469 28820 7503 28854
rect 7537 28820 7571 28854
rect 7605 28820 7639 28854
rect 7673 28820 7707 28854
rect 7741 28820 7775 28854
rect 7809 28820 7843 28854
rect 7877 28820 7911 28854
rect 7945 28820 7979 28854
rect 8013 28820 8047 28854
rect 8081 28820 8115 28854
rect 8149 28820 8183 28854
rect 8217 28820 8251 28854
rect 8285 28820 8319 28854
rect 8353 28820 8387 28854
rect 8421 28820 8455 28854
rect 8489 28820 8523 28854
rect 8557 28820 8591 28854
rect 8625 28820 8659 28854
rect 8693 28820 8727 28854
rect 8761 28820 8795 28854
rect 8829 28820 8863 28854
rect 8897 28820 8931 28854
rect 8965 28820 8999 28854
rect 9033 28820 9067 28854
rect 9101 28820 9135 28854
rect 9169 28820 9203 28854
rect 9237 28820 9271 28854
rect 9305 28820 9339 28854
rect 9373 28820 9407 28854
rect 9441 28820 9475 28854
rect 9509 28820 9543 28854
rect 9577 28820 9611 28854
rect 9645 28820 9679 28854
rect 9713 28820 9747 28854
rect 9781 28820 9815 28854
rect 9849 28820 9883 28854
rect 9917 28820 9951 28854
rect 9985 28820 10019 28854
rect 10053 28820 10087 28854
rect 10121 28820 10155 28854
rect 10189 28820 10223 28854
rect 10257 28820 10291 28854
rect 10325 28820 10359 28854
rect 10393 28820 10427 28854
rect 10461 28820 10495 28854
rect 10529 28820 10563 28854
rect 10597 28820 10631 28854
rect 10665 28820 10699 28854
rect 10733 28820 10767 28854
rect 10801 28820 10835 28854
rect 10869 28820 10903 28854
rect 10937 28820 10971 28854
rect 11005 28820 11039 28854
rect 11073 28820 11107 28854
rect 11141 28820 11175 28854
rect 11209 28820 11243 28854
rect 11277 28820 11311 28854
rect 11345 28820 11379 28854
rect 11413 28820 11447 28854
rect 11481 28820 11515 28854
rect 11549 28820 11583 28854
rect 11617 28820 11651 28854
rect 11685 28820 11719 28854
rect 11753 28820 11787 28854
rect 11821 28820 11855 28854
rect 11889 28820 11923 28854
rect 11957 28820 11991 28854
rect 12025 28820 12059 28854
rect 12093 28820 12127 28854
rect 12161 28820 12195 28854
rect 12229 28820 12263 28854
rect 12297 28820 12331 28854
rect 12365 28820 12399 28854
rect 12433 28820 12467 28854
rect 12501 28820 12535 28854
rect 12569 28820 12603 28854
rect 12637 28820 12671 28854
rect 12705 28820 12739 28854
rect 12773 28820 12807 28854
rect 12841 28820 12875 28854
rect 12909 28820 12943 28854
rect 12977 28820 12993 28854
rect 5163 28804 12993 28820
rect 5163 28799 5199 28804
rect 5433 28799 5469 28804
rect 5999 28799 6035 28804
rect 6269 28799 6305 28804
rect 6835 28799 6871 28804
rect 7105 28799 7141 28804
rect 7671 28799 7707 28804
rect 7941 28799 7977 28804
rect 8507 28799 8543 28804
rect 8777 28799 8813 28804
rect 9343 28799 9379 28804
rect 9613 28799 9649 28804
rect 10179 28799 10215 28804
rect 10449 28799 10485 28804
rect 11015 28799 11051 28804
rect 11285 28799 11321 28804
rect 11851 28799 11887 28804
rect 12121 28799 12157 28804
rect 12687 28799 12723 28804
rect 12957 28799 12993 28804
rect 5163 27340 5199 27371
rect 5433 27340 5469 27371
rect 5999 27340 6035 27371
rect 6269 27340 6305 27371
rect 6835 27340 6871 27371
rect 7105 27340 7141 27371
rect 7671 27340 7707 27371
rect 7941 27340 7977 27371
rect 8507 27340 8543 27371
rect 8777 27340 8813 27371
rect 9343 27340 9379 27371
rect 9613 27340 9649 27371
rect 10179 27340 10215 27371
rect 10449 27340 10485 27371
rect 11015 27340 11051 27371
rect 11285 27340 11321 27371
rect 11851 27340 11887 27371
rect 12121 27340 12157 27371
rect 12687 27340 12723 27371
rect 12957 27340 12993 27371
rect 5163 27324 12993 27340
rect 5163 27290 5179 27324
rect 5213 27290 5248 27324
rect 5282 27290 5317 27324
rect 5351 27290 5386 27324
rect 5420 27290 5455 27324
rect 5489 27290 5524 27324
rect 5558 27290 5593 27324
rect 5627 27290 5662 27324
rect 5696 27290 5731 27324
rect 5765 27290 5800 27324
rect 5834 27290 5869 27324
rect 5903 27290 5938 27324
rect 5972 27290 6007 27324
rect 6041 27290 6075 27324
rect 6109 27290 6143 27324
rect 6177 27290 6211 27324
rect 6245 27290 6279 27324
rect 6313 27290 6347 27324
rect 6381 27290 6415 27324
rect 6449 27290 6483 27324
rect 6517 27290 6551 27324
rect 6585 27290 6619 27324
rect 6653 27290 6687 27324
rect 6721 27290 6755 27324
rect 6789 27290 6823 27324
rect 6857 27290 6891 27324
rect 6925 27290 6959 27324
rect 6993 27290 7027 27324
rect 7061 27290 7095 27324
rect 7129 27290 7163 27324
rect 7197 27290 7231 27324
rect 7265 27290 7299 27324
rect 7333 27290 7367 27324
rect 7401 27290 7435 27324
rect 7469 27290 7503 27324
rect 7537 27290 7571 27324
rect 7605 27290 7639 27324
rect 7673 27290 7707 27324
rect 7741 27290 7775 27324
rect 7809 27290 7843 27324
rect 7877 27290 7911 27324
rect 7945 27290 7979 27324
rect 8013 27290 8047 27324
rect 8081 27290 8115 27324
rect 8149 27290 8183 27324
rect 8217 27290 8251 27324
rect 8285 27290 8319 27324
rect 8353 27290 8387 27324
rect 8421 27290 8455 27324
rect 8489 27290 8523 27324
rect 8557 27290 8591 27324
rect 8625 27290 8659 27324
rect 8693 27290 8727 27324
rect 8761 27290 8795 27324
rect 8829 27290 8863 27324
rect 8897 27290 8931 27324
rect 8965 27290 8999 27324
rect 9033 27290 9067 27324
rect 9101 27290 9135 27324
rect 9169 27290 9203 27324
rect 9237 27290 9271 27324
rect 9305 27290 9339 27324
rect 9373 27290 9407 27324
rect 9441 27290 9475 27324
rect 9509 27290 9543 27324
rect 9577 27290 9611 27324
rect 9645 27290 9679 27324
rect 9713 27290 9747 27324
rect 9781 27290 9815 27324
rect 9849 27290 9883 27324
rect 9917 27290 9951 27324
rect 9985 27290 10019 27324
rect 10053 27290 10087 27324
rect 10121 27290 10155 27324
rect 10189 27290 10223 27324
rect 10257 27290 10291 27324
rect 10325 27290 10359 27324
rect 10393 27290 10427 27324
rect 10461 27290 10495 27324
rect 10529 27290 10563 27324
rect 10597 27290 10631 27324
rect 10665 27290 10699 27324
rect 10733 27290 10767 27324
rect 10801 27290 10835 27324
rect 10869 27290 10903 27324
rect 10937 27290 10971 27324
rect 11005 27290 11039 27324
rect 11073 27290 11107 27324
rect 11141 27290 11175 27324
rect 11209 27290 11243 27324
rect 11277 27290 11311 27324
rect 11345 27290 11379 27324
rect 11413 27290 11447 27324
rect 11481 27290 11515 27324
rect 11549 27290 11583 27324
rect 11617 27290 11651 27324
rect 11685 27290 11719 27324
rect 11753 27290 11787 27324
rect 11821 27290 11855 27324
rect 11889 27290 11923 27324
rect 11957 27290 11991 27324
rect 12025 27290 12059 27324
rect 12093 27290 12127 27324
rect 12161 27290 12195 27324
rect 12229 27290 12263 27324
rect 12297 27290 12331 27324
rect 12365 27290 12399 27324
rect 12433 27290 12467 27324
rect 12501 27290 12535 27324
rect 12569 27290 12603 27324
rect 12637 27290 12671 27324
rect 12705 27290 12739 27324
rect 12773 27290 12807 27324
rect 12841 27290 12875 27324
rect 12909 27290 12943 27324
rect 12977 27290 12993 27324
rect 5163 27274 12993 27290
rect 5163 26870 5199 27274
rect 5433 26870 5469 27274
rect 5999 26870 6035 27274
rect 6269 26870 6305 27274
rect 6835 26870 6871 27274
rect 7105 26870 7141 27274
rect 7671 26870 7707 27274
rect 7941 26870 7977 27274
rect 8507 26870 8543 27274
rect 8777 26870 8813 27274
rect 9343 26870 9379 27274
rect 9613 26870 9649 27274
rect 10179 26870 10215 27274
rect 10449 26870 10485 27274
rect 11015 26870 11051 27274
rect 11285 26870 11321 27274
rect 11851 26870 11887 27274
rect 12121 26870 12157 27274
rect 12687 26870 12723 27274
rect 12957 26870 12993 27274
rect 5163 26854 12993 26870
rect 5163 26820 5179 26854
rect 5213 26820 5248 26854
rect 5282 26820 5317 26854
rect 5351 26820 5386 26854
rect 5420 26820 5455 26854
rect 5489 26820 5524 26854
rect 5558 26820 5593 26854
rect 5627 26820 5662 26854
rect 5696 26820 5731 26854
rect 5765 26820 5800 26854
rect 5834 26820 5869 26854
rect 5903 26820 5938 26854
rect 5972 26820 6007 26854
rect 6041 26820 6075 26854
rect 6109 26820 6143 26854
rect 6177 26820 6211 26854
rect 6245 26820 6279 26854
rect 6313 26820 6347 26854
rect 6381 26820 6415 26854
rect 6449 26820 6483 26854
rect 6517 26820 6551 26854
rect 6585 26820 6619 26854
rect 6653 26820 6687 26854
rect 6721 26820 6755 26854
rect 6789 26820 6823 26854
rect 6857 26820 6891 26854
rect 6925 26820 6959 26854
rect 6993 26820 7027 26854
rect 7061 26820 7095 26854
rect 7129 26820 7163 26854
rect 7197 26820 7231 26854
rect 7265 26820 7299 26854
rect 7333 26820 7367 26854
rect 7401 26820 7435 26854
rect 7469 26820 7503 26854
rect 7537 26820 7571 26854
rect 7605 26820 7639 26854
rect 7673 26820 7707 26854
rect 7741 26820 7775 26854
rect 7809 26820 7843 26854
rect 7877 26820 7911 26854
rect 7945 26820 7979 26854
rect 8013 26820 8047 26854
rect 8081 26820 8115 26854
rect 8149 26820 8183 26854
rect 8217 26820 8251 26854
rect 8285 26820 8319 26854
rect 8353 26820 8387 26854
rect 8421 26820 8455 26854
rect 8489 26820 8523 26854
rect 8557 26820 8591 26854
rect 8625 26820 8659 26854
rect 8693 26820 8727 26854
rect 8761 26820 8795 26854
rect 8829 26820 8863 26854
rect 8897 26820 8931 26854
rect 8965 26820 8999 26854
rect 9033 26820 9067 26854
rect 9101 26820 9135 26854
rect 9169 26820 9203 26854
rect 9237 26820 9271 26854
rect 9305 26820 9339 26854
rect 9373 26820 9407 26854
rect 9441 26820 9475 26854
rect 9509 26820 9543 26854
rect 9577 26820 9611 26854
rect 9645 26820 9679 26854
rect 9713 26820 9747 26854
rect 9781 26820 9815 26854
rect 9849 26820 9883 26854
rect 9917 26820 9951 26854
rect 9985 26820 10019 26854
rect 10053 26820 10087 26854
rect 10121 26820 10155 26854
rect 10189 26820 10223 26854
rect 10257 26820 10291 26854
rect 10325 26820 10359 26854
rect 10393 26820 10427 26854
rect 10461 26820 10495 26854
rect 10529 26820 10563 26854
rect 10597 26820 10631 26854
rect 10665 26820 10699 26854
rect 10733 26820 10767 26854
rect 10801 26820 10835 26854
rect 10869 26820 10903 26854
rect 10937 26820 10971 26854
rect 11005 26820 11039 26854
rect 11073 26820 11107 26854
rect 11141 26820 11175 26854
rect 11209 26820 11243 26854
rect 11277 26820 11311 26854
rect 11345 26820 11379 26854
rect 11413 26820 11447 26854
rect 11481 26820 11515 26854
rect 11549 26820 11583 26854
rect 11617 26820 11651 26854
rect 11685 26820 11719 26854
rect 11753 26820 11787 26854
rect 11821 26820 11855 26854
rect 11889 26820 11923 26854
rect 11957 26820 11991 26854
rect 12025 26820 12059 26854
rect 12093 26820 12127 26854
rect 12161 26820 12195 26854
rect 12229 26820 12263 26854
rect 12297 26820 12331 26854
rect 12365 26820 12399 26854
rect 12433 26820 12467 26854
rect 12501 26820 12535 26854
rect 12569 26820 12603 26854
rect 12637 26820 12671 26854
rect 12705 26820 12739 26854
rect 12773 26820 12807 26854
rect 12841 26820 12875 26854
rect 12909 26820 12943 26854
rect 12977 26820 12993 26854
rect 5163 26804 12993 26820
rect 5163 26783 5199 26804
rect 5433 26783 5469 26804
rect 5999 26783 6035 26804
rect 6269 26783 6305 26804
rect 6835 26783 6871 26804
rect 7105 26783 7141 26804
rect 7671 26783 7707 26804
rect 7941 26783 7977 26804
rect 8507 26783 8543 26804
rect 8777 26783 8813 26804
rect 9343 26783 9379 26804
rect 9613 26783 9649 26804
rect 10179 26783 10215 26804
rect 10449 26783 10485 26804
rect 11015 26783 11051 26804
rect 11285 26783 11321 26804
rect 11851 26783 11887 26804
rect 12121 26783 12157 26804
rect 12687 26783 12723 26804
rect 12957 26783 12993 26804
rect 5163 25703 12993 25719
rect 5163 25669 5179 25703
rect 5213 25669 5248 25703
rect 5282 25669 5317 25703
rect 5351 25669 5386 25703
rect 5420 25669 5455 25703
rect 5489 25669 5524 25703
rect 5558 25669 5593 25703
rect 5627 25669 5662 25703
rect 5696 25669 5731 25703
rect 5765 25669 5800 25703
rect 5834 25669 5869 25703
rect 5903 25669 5938 25703
rect 5972 25669 6007 25703
rect 6041 25669 6075 25703
rect 6109 25669 6143 25703
rect 6177 25669 6211 25703
rect 6245 25669 6279 25703
rect 6313 25669 6347 25703
rect 6381 25669 6415 25703
rect 6449 25669 6483 25703
rect 6517 25669 6551 25703
rect 6585 25669 6619 25703
rect 6653 25669 6687 25703
rect 6721 25669 6755 25703
rect 6789 25669 6823 25703
rect 6857 25669 6891 25703
rect 6925 25669 6959 25703
rect 6993 25669 7027 25703
rect 7061 25669 7095 25703
rect 7129 25669 7163 25703
rect 7197 25669 7231 25703
rect 7265 25669 7299 25703
rect 7333 25669 7367 25703
rect 7401 25669 7435 25703
rect 7469 25669 7503 25703
rect 7537 25669 7571 25703
rect 7605 25669 7639 25703
rect 7673 25669 7707 25703
rect 7741 25669 7775 25703
rect 7809 25669 7843 25703
rect 7877 25669 7911 25703
rect 7945 25669 7979 25703
rect 8013 25669 8047 25703
rect 8081 25669 8115 25703
rect 8149 25669 8183 25703
rect 8217 25669 8251 25703
rect 8285 25669 8319 25703
rect 8353 25669 8387 25703
rect 8421 25669 8455 25703
rect 8489 25669 8523 25703
rect 8557 25669 8591 25703
rect 8625 25669 8659 25703
rect 8693 25669 8727 25703
rect 8761 25669 8795 25703
rect 8829 25669 8863 25703
rect 8897 25669 8931 25703
rect 8965 25669 8999 25703
rect 9033 25669 9067 25703
rect 9101 25669 9135 25703
rect 9169 25669 9203 25703
rect 9237 25669 9271 25703
rect 9305 25669 9339 25703
rect 9373 25669 9407 25703
rect 9441 25669 9475 25703
rect 9509 25669 9543 25703
rect 9577 25669 9611 25703
rect 9645 25669 9679 25703
rect 9713 25669 9747 25703
rect 9781 25669 9815 25703
rect 9849 25669 9883 25703
rect 9917 25669 9951 25703
rect 9985 25669 10019 25703
rect 10053 25669 10087 25703
rect 10121 25669 10155 25703
rect 10189 25669 10223 25703
rect 10257 25669 10291 25703
rect 10325 25669 10359 25703
rect 10393 25669 10427 25703
rect 10461 25669 10495 25703
rect 10529 25669 10563 25703
rect 10597 25669 10631 25703
rect 10665 25669 10699 25703
rect 10733 25669 10767 25703
rect 10801 25669 10835 25703
rect 10869 25669 10903 25703
rect 10937 25669 10971 25703
rect 11005 25669 11039 25703
rect 11073 25669 11107 25703
rect 11141 25669 11175 25703
rect 11209 25669 11243 25703
rect 11277 25669 11311 25703
rect 11345 25669 11379 25703
rect 11413 25669 11447 25703
rect 11481 25669 11515 25703
rect 11549 25669 11583 25703
rect 11617 25669 11651 25703
rect 11685 25669 11719 25703
rect 11753 25669 11787 25703
rect 11821 25669 11855 25703
rect 11889 25669 11923 25703
rect 11957 25669 11991 25703
rect 12025 25669 12059 25703
rect 12093 25669 12127 25703
rect 12161 25669 12195 25703
rect 12229 25669 12263 25703
rect 12297 25669 12331 25703
rect 12365 25669 12399 25703
rect 12433 25669 12467 25703
rect 12501 25669 12535 25703
rect 12569 25669 12603 25703
rect 12637 25669 12671 25703
rect 12705 25669 12739 25703
rect 12773 25669 12807 25703
rect 12841 25669 12875 25703
rect 12909 25669 12943 25703
rect 12977 25669 12993 25703
rect 5163 25653 12993 25669
rect 4934 23697 13331 23713
rect 4934 23663 4954 23697
rect 4988 23663 5022 23697
rect 5056 23663 5090 23697
rect 5124 23663 5158 23697
rect 5192 23663 5226 23697
rect 5260 23663 5294 23697
rect 5328 23663 5362 23697
rect 5396 23663 5430 23697
rect 5464 23663 5498 23697
rect 5532 23663 5566 23697
rect 5600 23663 5634 23697
rect 5668 23663 5702 23697
rect 5736 23663 5770 23697
rect 5804 23663 5838 23697
rect 5872 23663 5906 23697
rect 5940 23663 5974 23697
rect 6008 23663 6042 23697
rect 6076 23663 6110 23697
rect 6144 23663 6178 23697
rect 6212 23663 6246 23697
rect 6280 23663 6314 23697
rect 6348 23663 6382 23697
rect 6416 23663 6450 23697
rect 6484 23663 6518 23697
rect 6552 23663 6586 23697
rect 6620 23663 6654 23697
rect 6688 23663 6722 23697
rect 6756 23663 6790 23697
rect 6824 23663 6858 23697
rect 6892 23663 6926 23697
rect 6960 23663 6994 23697
rect 7028 23663 7062 23697
rect 7096 23663 7130 23697
rect 7164 23663 7198 23697
rect 7232 23663 7266 23697
rect 7300 23663 7334 23697
rect 7368 23663 7402 23697
rect 7436 23663 7470 23697
rect 7504 23663 7538 23697
rect 7572 23663 7606 23697
rect 7640 23663 7674 23697
rect 7708 23663 7742 23697
rect 7776 23663 7810 23697
rect 7844 23663 7878 23697
rect 7912 23663 7946 23697
rect 7980 23663 8014 23697
rect 8048 23663 8082 23697
rect 8116 23663 8150 23697
rect 8184 23663 8218 23697
rect 8252 23663 8286 23697
rect 8320 23663 8354 23697
rect 8388 23663 8422 23697
rect 8456 23663 8490 23697
rect 8524 23663 8558 23697
rect 8592 23663 8626 23697
rect 8660 23663 8694 23697
rect 8728 23663 8762 23697
rect 8796 23663 8830 23697
rect 8864 23663 8898 23697
rect 8932 23663 8966 23697
rect 9000 23663 9034 23697
rect 9068 23663 9102 23697
rect 9136 23663 9170 23697
rect 9204 23663 9238 23697
rect 9272 23663 9306 23697
rect 9340 23663 9374 23697
rect 9408 23663 9442 23697
rect 9476 23663 9510 23697
rect 9544 23663 9578 23697
rect 9612 23663 9646 23697
rect 9680 23663 9714 23697
rect 9748 23663 9782 23697
rect 9816 23663 9850 23697
rect 9884 23663 9918 23697
rect 9952 23663 9986 23697
rect 10020 23663 10054 23697
rect 10088 23663 10122 23697
rect 10156 23663 10190 23697
rect 10224 23663 10258 23697
rect 10292 23663 10326 23697
rect 10360 23663 10394 23697
rect 10428 23663 10462 23697
rect 10496 23663 10530 23697
rect 10564 23663 10598 23697
rect 10632 23663 10666 23697
rect 10700 23663 10734 23697
rect 10768 23663 10802 23697
rect 10836 23663 10870 23697
rect 10904 23663 10938 23697
rect 10972 23663 11006 23697
rect 11040 23663 11074 23697
rect 11108 23663 11142 23697
rect 11176 23663 11210 23697
rect 11244 23663 11278 23697
rect 11312 23663 11346 23697
rect 11380 23663 11414 23697
rect 11448 23663 11482 23697
rect 11516 23663 11550 23697
rect 11584 23663 11618 23697
rect 11652 23663 11686 23697
rect 11720 23663 11754 23697
rect 11788 23663 11822 23697
rect 11856 23663 11890 23697
rect 11924 23663 11958 23697
rect 11992 23663 12026 23697
rect 12060 23663 12094 23697
rect 12128 23663 12162 23697
rect 12196 23663 12230 23697
rect 12264 23663 12298 23697
rect 12332 23663 12366 23697
rect 12400 23663 12434 23697
rect 12468 23663 12502 23697
rect 12536 23663 12570 23697
rect 12604 23663 12638 23697
rect 12672 23663 12706 23697
rect 12740 23663 12774 23697
rect 12808 23663 12842 23697
rect 12876 23663 12910 23697
rect 12944 23663 12978 23697
rect 13012 23663 13046 23697
rect 13080 23663 13114 23697
rect 13148 23663 13182 23697
rect 13216 23663 13250 23697
rect 13284 23663 13331 23697
rect 4934 23647 13331 23663
rect 4934 23462 13331 23478
rect 4934 23428 4954 23462
rect 4988 23428 5022 23462
rect 5056 23428 5090 23462
rect 5124 23428 5158 23462
rect 5192 23428 5226 23462
rect 5260 23428 5294 23462
rect 5328 23428 5362 23462
rect 5396 23428 5430 23462
rect 5464 23428 5498 23462
rect 5532 23428 5566 23462
rect 5600 23428 5634 23462
rect 5668 23428 5702 23462
rect 5736 23428 5770 23462
rect 5804 23428 5838 23462
rect 5872 23428 5906 23462
rect 5940 23428 5974 23462
rect 6008 23428 6042 23462
rect 6076 23428 6110 23462
rect 6144 23428 6178 23462
rect 6212 23428 6246 23462
rect 6280 23428 6314 23462
rect 6348 23428 6382 23462
rect 6416 23428 6450 23462
rect 6484 23428 6518 23462
rect 6552 23428 6586 23462
rect 6620 23428 6654 23462
rect 6688 23428 6722 23462
rect 6756 23428 6790 23462
rect 6824 23428 6858 23462
rect 6892 23428 6926 23462
rect 6960 23428 6994 23462
rect 7028 23428 7062 23462
rect 7096 23428 7130 23462
rect 7164 23428 7198 23462
rect 7232 23428 7266 23462
rect 7300 23428 7334 23462
rect 7368 23428 7402 23462
rect 7436 23428 7470 23462
rect 7504 23428 7538 23462
rect 7572 23428 7606 23462
rect 7640 23428 7674 23462
rect 7708 23428 7742 23462
rect 7776 23428 7810 23462
rect 7844 23428 7878 23462
rect 7912 23428 7946 23462
rect 7980 23428 8014 23462
rect 8048 23428 8082 23462
rect 8116 23428 8150 23462
rect 8184 23428 8218 23462
rect 8252 23428 8286 23462
rect 8320 23428 8354 23462
rect 8388 23428 8422 23462
rect 8456 23428 8490 23462
rect 8524 23428 8558 23462
rect 8592 23428 8626 23462
rect 8660 23428 8694 23462
rect 8728 23428 8762 23462
rect 8796 23428 8830 23462
rect 8864 23428 8898 23462
rect 8932 23428 8966 23462
rect 9000 23428 9034 23462
rect 9068 23428 9102 23462
rect 9136 23428 9170 23462
rect 9204 23428 9238 23462
rect 9272 23428 9306 23462
rect 9340 23428 9374 23462
rect 9408 23428 9442 23462
rect 9476 23428 9510 23462
rect 9544 23428 9578 23462
rect 9612 23428 9646 23462
rect 9680 23428 9714 23462
rect 9748 23428 9782 23462
rect 9816 23428 9850 23462
rect 9884 23428 9918 23462
rect 9952 23428 9986 23462
rect 10020 23428 10054 23462
rect 10088 23428 10122 23462
rect 10156 23428 10190 23462
rect 10224 23428 10258 23462
rect 10292 23428 10326 23462
rect 10360 23428 10394 23462
rect 10428 23428 10462 23462
rect 10496 23428 10530 23462
rect 10564 23428 10598 23462
rect 10632 23428 10666 23462
rect 10700 23428 10734 23462
rect 10768 23428 10802 23462
rect 10836 23428 10870 23462
rect 10904 23428 10938 23462
rect 10972 23428 11006 23462
rect 11040 23428 11074 23462
rect 11108 23428 11142 23462
rect 11176 23428 11210 23462
rect 11244 23428 11278 23462
rect 11312 23428 11346 23462
rect 11380 23428 11414 23462
rect 11448 23428 11482 23462
rect 11516 23428 11550 23462
rect 11584 23428 11618 23462
rect 11652 23428 11686 23462
rect 11720 23428 11754 23462
rect 11788 23428 11822 23462
rect 11856 23428 11890 23462
rect 11924 23428 11958 23462
rect 11992 23428 12026 23462
rect 12060 23428 12094 23462
rect 12128 23428 12162 23462
rect 12196 23428 12230 23462
rect 12264 23428 12298 23462
rect 12332 23428 12366 23462
rect 12400 23428 12434 23462
rect 12468 23428 12502 23462
rect 12536 23428 12570 23462
rect 12604 23428 12638 23462
rect 12672 23428 12706 23462
rect 12740 23428 12774 23462
rect 12808 23428 12842 23462
rect 12876 23428 12910 23462
rect 12944 23428 12978 23462
rect 13012 23428 13046 23462
rect 13080 23428 13114 23462
rect 13148 23428 13182 23462
rect 13216 23428 13250 23462
rect 13284 23428 13331 23462
rect 4934 23412 13331 23428
rect 4934 21763 13331 21779
rect 4934 21729 4954 21763
rect 4988 21729 5022 21763
rect 5056 21729 5090 21763
rect 5124 21729 5158 21763
rect 5192 21729 5226 21763
rect 5260 21729 5294 21763
rect 5328 21729 5362 21763
rect 5396 21729 5430 21763
rect 5464 21729 5498 21763
rect 5532 21729 5566 21763
rect 5600 21729 5634 21763
rect 5668 21729 5702 21763
rect 5736 21729 5770 21763
rect 5804 21729 5838 21763
rect 5872 21729 5906 21763
rect 5940 21729 5974 21763
rect 6008 21729 6042 21763
rect 6076 21729 6110 21763
rect 6144 21729 6178 21763
rect 6212 21729 6246 21763
rect 6280 21729 6314 21763
rect 6348 21729 6382 21763
rect 6416 21729 6450 21763
rect 6484 21729 6518 21763
rect 6552 21729 6586 21763
rect 6620 21729 6654 21763
rect 6688 21729 6722 21763
rect 6756 21729 6790 21763
rect 6824 21729 6858 21763
rect 6892 21729 6926 21763
rect 6960 21729 6994 21763
rect 7028 21729 7062 21763
rect 7096 21729 7130 21763
rect 7164 21729 7198 21763
rect 7232 21729 7266 21763
rect 7300 21729 7334 21763
rect 7368 21729 7402 21763
rect 7436 21729 7470 21763
rect 7504 21729 7538 21763
rect 7572 21729 7606 21763
rect 7640 21729 7674 21763
rect 7708 21729 7742 21763
rect 7776 21729 7810 21763
rect 7844 21729 7878 21763
rect 7912 21729 7946 21763
rect 7980 21729 8014 21763
rect 8048 21729 8082 21763
rect 8116 21729 8150 21763
rect 8184 21729 8218 21763
rect 8252 21729 8286 21763
rect 8320 21729 8354 21763
rect 8388 21729 8422 21763
rect 8456 21729 8490 21763
rect 8524 21729 8558 21763
rect 8592 21729 8626 21763
rect 8660 21729 8694 21763
rect 8728 21729 8762 21763
rect 8796 21729 8830 21763
rect 8864 21729 8898 21763
rect 8932 21729 8966 21763
rect 9000 21729 9034 21763
rect 9068 21729 9102 21763
rect 9136 21729 9170 21763
rect 9204 21729 9238 21763
rect 9272 21729 9306 21763
rect 9340 21729 9374 21763
rect 9408 21729 9442 21763
rect 9476 21729 9510 21763
rect 9544 21729 9578 21763
rect 9612 21729 9646 21763
rect 9680 21729 9714 21763
rect 9748 21729 9782 21763
rect 9816 21729 9850 21763
rect 9884 21729 9918 21763
rect 9952 21729 9986 21763
rect 10020 21729 10054 21763
rect 10088 21729 10122 21763
rect 10156 21729 10190 21763
rect 10224 21729 10258 21763
rect 10292 21729 10326 21763
rect 10360 21729 10394 21763
rect 10428 21729 10462 21763
rect 10496 21729 10530 21763
rect 10564 21729 10598 21763
rect 10632 21729 10666 21763
rect 10700 21729 10734 21763
rect 10768 21729 10802 21763
rect 10836 21729 10870 21763
rect 10904 21729 10938 21763
rect 10972 21729 11006 21763
rect 11040 21729 11074 21763
rect 11108 21729 11142 21763
rect 11176 21729 11210 21763
rect 11244 21729 11278 21763
rect 11312 21729 11346 21763
rect 11380 21729 11414 21763
rect 11448 21729 11482 21763
rect 11516 21729 11550 21763
rect 11584 21729 11618 21763
rect 11652 21729 11686 21763
rect 11720 21729 11754 21763
rect 11788 21729 11822 21763
rect 11856 21729 11890 21763
rect 11924 21729 11958 21763
rect 11992 21729 12026 21763
rect 12060 21729 12094 21763
rect 12128 21729 12162 21763
rect 12196 21729 12230 21763
rect 12264 21729 12298 21763
rect 12332 21729 12366 21763
rect 12400 21729 12434 21763
rect 12468 21729 12502 21763
rect 12536 21729 12570 21763
rect 12604 21729 12638 21763
rect 12672 21729 12706 21763
rect 12740 21729 12774 21763
rect 12808 21729 12842 21763
rect 12876 21729 12910 21763
rect 12944 21729 12978 21763
rect 13012 21729 13046 21763
rect 13080 21729 13114 21763
rect 13148 21729 13182 21763
rect 13216 21729 13250 21763
rect 13284 21729 13331 21763
rect 4934 21713 13331 21729
rect 4923 19742 13331 19758
rect 4923 19708 4943 19742
rect 4977 19708 5011 19742
rect 5045 19708 5079 19742
rect 5113 19708 5147 19742
rect 5181 19708 5215 19742
rect 5249 19708 5283 19742
rect 5317 19708 5351 19742
rect 5385 19708 5419 19742
rect 5453 19708 5487 19742
rect 5521 19708 5555 19742
rect 5589 19708 5623 19742
rect 5657 19708 5691 19742
rect 5725 19708 5759 19742
rect 5793 19708 5827 19742
rect 5861 19708 5895 19742
rect 5929 19708 5963 19742
rect 5997 19708 6031 19742
rect 6065 19708 6099 19742
rect 6133 19708 6167 19742
rect 6201 19708 6235 19742
rect 6269 19708 6303 19742
rect 6337 19708 6371 19742
rect 6405 19708 6439 19742
rect 6473 19708 6507 19742
rect 6541 19708 6575 19742
rect 6609 19708 6643 19742
rect 6677 19708 6711 19742
rect 6745 19708 6779 19742
rect 6813 19708 6847 19742
rect 6881 19708 6915 19742
rect 6949 19708 6983 19742
rect 7017 19708 7051 19742
rect 7085 19708 7119 19742
rect 7153 19708 7187 19742
rect 7221 19708 7255 19742
rect 7289 19708 7323 19742
rect 7357 19708 7391 19742
rect 7425 19708 7459 19742
rect 7493 19708 7527 19742
rect 7561 19708 7595 19742
rect 7629 19708 7663 19742
rect 7697 19708 7731 19742
rect 7765 19708 7799 19742
rect 7833 19708 7867 19742
rect 7901 19708 7935 19742
rect 7969 19708 8003 19742
rect 8037 19708 8071 19742
rect 8105 19708 8139 19742
rect 8173 19708 8207 19742
rect 8241 19708 8275 19742
rect 8309 19708 8343 19742
rect 8377 19708 8411 19742
rect 8445 19708 8479 19742
rect 8513 19708 8547 19742
rect 8581 19708 8615 19742
rect 8649 19708 8683 19742
rect 8717 19708 8751 19742
rect 8785 19708 8819 19742
rect 8853 19708 8887 19742
rect 8921 19708 8955 19742
rect 8989 19708 9023 19742
rect 9057 19708 9091 19742
rect 9125 19708 9159 19742
rect 9193 19708 9227 19742
rect 9261 19708 9295 19742
rect 9329 19708 9363 19742
rect 9397 19708 9431 19742
rect 9465 19708 9499 19742
rect 9533 19708 9567 19742
rect 9601 19708 9635 19742
rect 9669 19708 9703 19742
rect 9737 19708 9771 19742
rect 9805 19708 9839 19742
rect 9873 19708 9907 19742
rect 9941 19708 9975 19742
rect 10009 19708 10043 19742
rect 10077 19708 10111 19742
rect 10145 19708 10179 19742
rect 10213 19708 10247 19742
rect 10281 19708 10315 19742
rect 10349 19708 10383 19742
rect 10417 19708 10451 19742
rect 10485 19708 10519 19742
rect 10553 19708 10587 19742
rect 10621 19708 10655 19742
rect 10689 19708 10723 19742
rect 10757 19708 10791 19742
rect 10825 19708 10859 19742
rect 10893 19708 10927 19742
rect 10961 19708 10995 19742
rect 11029 19708 11063 19742
rect 11097 19708 11131 19742
rect 11165 19708 11199 19742
rect 11233 19708 11267 19742
rect 11301 19708 11335 19742
rect 11369 19708 11403 19742
rect 11437 19708 11471 19742
rect 11505 19708 11539 19742
rect 11573 19708 11607 19742
rect 11641 19708 11675 19742
rect 11709 19708 11743 19742
rect 11777 19708 11811 19742
rect 11845 19708 11879 19742
rect 11913 19708 11947 19742
rect 11981 19708 12015 19742
rect 12049 19708 12083 19742
rect 12117 19708 12151 19742
rect 12185 19708 12219 19742
rect 12253 19708 12287 19742
rect 12321 19708 12355 19742
rect 12389 19708 12423 19742
rect 12457 19708 12491 19742
rect 12525 19708 12559 19742
rect 12593 19708 12627 19742
rect 12661 19708 12695 19742
rect 12729 19708 12763 19742
rect 12797 19708 12831 19742
rect 12865 19708 12899 19742
rect 12933 19708 12967 19742
rect 13001 19708 13035 19742
rect 13069 19708 13103 19742
rect 13137 19708 13171 19742
rect 13205 19708 13239 19742
rect 13273 19708 13331 19742
rect 4923 19692 13331 19708
rect 4923 18043 13331 18059
rect 4923 18009 4943 18043
rect 4977 18009 5011 18043
rect 5045 18009 5079 18043
rect 5113 18009 5147 18043
rect 5181 18009 5215 18043
rect 5249 18009 5283 18043
rect 5317 18009 5351 18043
rect 5385 18009 5419 18043
rect 5453 18009 5487 18043
rect 5521 18009 5555 18043
rect 5589 18009 5623 18043
rect 5657 18009 5691 18043
rect 5725 18009 5759 18043
rect 5793 18009 5827 18043
rect 5861 18009 5895 18043
rect 5929 18009 5963 18043
rect 5997 18009 6031 18043
rect 6065 18009 6099 18043
rect 6133 18009 6167 18043
rect 6201 18009 6235 18043
rect 6269 18009 6303 18043
rect 6337 18009 6371 18043
rect 6405 18009 6439 18043
rect 6473 18009 6507 18043
rect 6541 18009 6575 18043
rect 6609 18009 6643 18043
rect 6677 18009 6711 18043
rect 6745 18009 6779 18043
rect 6813 18009 6847 18043
rect 6881 18009 6915 18043
rect 6949 18009 6983 18043
rect 7017 18009 7051 18043
rect 7085 18009 7119 18043
rect 7153 18009 7187 18043
rect 7221 18009 7255 18043
rect 7289 18009 7323 18043
rect 7357 18009 7391 18043
rect 7425 18009 7459 18043
rect 7493 18009 7527 18043
rect 7561 18009 7595 18043
rect 7629 18009 7663 18043
rect 7697 18009 7731 18043
rect 7765 18009 7799 18043
rect 7833 18009 7867 18043
rect 7901 18009 7935 18043
rect 7969 18009 8003 18043
rect 8037 18009 8071 18043
rect 8105 18009 8139 18043
rect 8173 18009 8207 18043
rect 8241 18009 8275 18043
rect 8309 18009 8343 18043
rect 8377 18009 8411 18043
rect 8445 18009 8479 18043
rect 8513 18009 8547 18043
rect 8581 18009 8615 18043
rect 8649 18009 8683 18043
rect 8717 18009 8751 18043
rect 8785 18009 8819 18043
rect 8853 18009 8887 18043
rect 8921 18009 8955 18043
rect 8989 18009 9023 18043
rect 9057 18009 9091 18043
rect 9125 18009 9159 18043
rect 9193 18009 9227 18043
rect 9261 18009 9295 18043
rect 9329 18009 9363 18043
rect 9397 18009 9431 18043
rect 9465 18009 9499 18043
rect 9533 18009 9567 18043
rect 9601 18009 9635 18043
rect 9669 18009 9703 18043
rect 9737 18009 9771 18043
rect 9805 18009 9839 18043
rect 9873 18009 9907 18043
rect 9941 18009 9975 18043
rect 10009 18009 10043 18043
rect 10077 18009 10111 18043
rect 10145 18009 10179 18043
rect 10213 18009 10247 18043
rect 10281 18009 10315 18043
rect 10349 18009 10383 18043
rect 10417 18009 10451 18043
rect 10485 18009 10519 18043
rect 10553 18009 10587 18043
rect 10621 18009 10655 18043
rect 10689 18009 10723 18043
rect 10757 18009 10791 18043
rect 10825 18009 10859 18043
rect 10893 18009 10927 18043
rect 10961 18009 10995 18043
rect 11029 18009 11063 18043
rect 11097 18009 11131 18043
rect 11165 18009 11199 18043
rect 11233 18009 11267 18043
rect 11301 18009 11335 18043
rect 11369 18009 11403 18043
rect 11437 18009 11471 18043
rect 11505 18009 11539 18043
rect 11573 18009 11607 18043
rect 11641 18009 11675 18043
rect 11709 18009 11743 18043
rect 11777 18009 11811 18043
rect 11845 18009 11879 18043
rect 11913 18009 11947 18043
rect 11981 18009 12015 18043
rect 12049 18009 12083 18043
rect 12117 18009 12151 18043
rect 12185 18009 12219 18043
rect 12253 18009 12287 18043
rect 12321 18009 12355 18043
rect 12389 18009 12423 18043
rect 12457 18009 12491 18043
rect 12525 18009 12559 18043
rect 12593 18009 12627 18043
rect 12661 18009 12695 18043
rect 12729 18009 12763 18043
rect 12797 18009 12831 18043
rect 12865 18009 12899 18043
rect 12933 18009 12967 18043
rect 13001 18009 13035 18043
rect 13069 18009 13103 18043
rect 13137 18009 13171 18043
rect 13205 18009 13239 18043
rect 13273 18009 13331 18043
rect 4923 17993 13331 18009
rect 2595 16243 13331 16259
rect 2595 16209 2615 16243
rect 2649 16209 2683 16243
rect 2717 16209 2751 16243
rect 2785 16209 2819 16243
rect 2853 16209 2887 16243
rect 2921 16209 2955 16243
rect 2989 16209 3023 16243
rect 3057 16209 3091 16243
rect 3125 16209 3159 16243
rect 3193 16209 3227 16243
rect 3261 16209 3295 16243
rect 3329 16209 3363 16243
rect 3397 16209 3431 16243
rect 3465 16209 3499 16243
rect 3533 16209 3567 16243
rect 3601 16209 3635 16243
rect 3669 16209 3703 16243
rect 3737 16209 3771 16243
rect 3805 16209 3839 16243
rect 3873 16209 3907 16243
rect 3941 16209 3975 16243
rect 4009 16209 4043 16243
rect 4077 16209 4111 16243
rect 4145 16209 4179 16243
rect 4213 16209 4247 16243
rect 4281 16209 4315 16243
rect 4349 16209 4383 16243
rect 4417 16209 4451 16243
rect 4485 16209 4519 16243
rect 4553 16209 4587 16243
rect 4621 16209 4655 16243
rect 4689 16209 4723 16243
rect 4757 16209 4791 16243
rect 4825 16209 4859 16243
rect 4893 16209 4927 16243
rect 4961 16209 4995 16243
rect 5029 16209 5063 16243
rect 5097 16209 5131 16243
rect 5165 16209 5199 16243
rect 5233 16209 5267 16243
rect 5301 16209 5335 16243
rect 5369 16209 5403 16243
rect 5437 16209 5471 16243
rect 5505 16209 5539 16243
rect 5573 16209 5607 16243
rect 5641 16209 5675 16243
rect 5709 16209 5743 16243
rect 5777 16209 5811 16243
rect 5845 16209 5879 16243
rect 5913 16209 5947 16243
rect 5981 16209 6015 16243
rect 6049 16209 6083 16243
rect 6117 16209 6151 16243
rect 6185 16209 6219 16243
rect 6253 16209 6287 16243
rect 6321 16209 6355 16243
rect 6389 16209 6423 16243
rect 6457 16209 6491 16243
rect 6525 16209 6559 16243
rect 6593 16209 6627 16243
rect 6661 16209 6695 16243
rect 6729 16209 6763 16243
rect 6797 16209 6831 16243
rect 6865 16209 6899 16243
rect 6933 16209 6967 16243
rect 7001 16209 7035 16243
rect 7069 16209 7103 16243
rect 7137 16209 7171 16243
rect 7205 16209 7239 16243
rect 7273 16209 7307 16243
rect 7341 16209 7375 16243
rect 7409 16209 7443 16243
rect 7477 16209 7511 16243
rect 7545 16209 7579 16243
rect 7613 16209 7647 16243
rect 7681 16209 7715 16243
rect 7749 16209 7783 16243
rect 7817 16209 7851 16243
rect 7885 16209 7919 16243
rect 7953 16209 7987 16243
rect 8021 16209 8055 16243
rect 8089 16209 8123 16243
rect 8157 16209 8191 16243
rect 8225 16209 8259 16243
rect 8293 16209 8327 16243
rect 8361 16209 8395 16243
rect 8429 16209 8463 16243
rect 8497 16209 8531 16243
rect 8565 16209 8599 16243
rect 8633 16209 8667 16243
rect 8701 16209 8735 16243
rect 8769 16209 8803 16243
rect 8837 16209 8871 16243
rect 8905 16209 8939 16243
rect 8973 16209 9007 16243
rect 9041 16209 9075 16243
rect 9109 16209 9143 16243
rect 9177 16209 9211 16243
rect 9245 16209 9279 16243
rect 9313 16209 9347 16243
rect 9381 16209 9415 16243
rect 9449 16209 9483 16243
rect 9517 16209 9551 16243
rect 9585 16209 9619 16243
rect 9653 16209 9687 16243
rect 9721 16209 9755 16243
rect 9789 16209 9823 16243
rect 9857 16209 9891 16243
rect 9925 16209 9959 16243
rect 9993 16209 10027 16243
rect 10061 16209 10095 16243
rect 10129 16209 10163 16243
rect 10197 16209 10231 16243
rect 10265 16209 10299 16243
rect 10333 16209 10367 16243
rect 10401 16209 10435 16243
rect 10469 16209 10503 16243
rect 10537 16209 10571 16243
rect 10605 16209 10639 16243
rect 10673 16209 10707 16243
rect 10741 16209 10775 16243
rect 10809 16209 10843 16243
rect 10877 16209 10911 16243
rect 10945 16209 10979 16243
rect 11013 16209 11047 16243
rect 11081 16209 11115 16243
rect 11149 16209 11183 16243
rect 11217 16209 11251 16243
rect 11285 16209 11319 16243
rect 11353 16209 11387 16243
rect 11421 16209 11455 16243
rect 11489 16209 11523 16243
rect 11557 16209 11591 16243
rect 11625 16209 11659 16243
rect 11693 16209 11727 16243
rect 11761 16209 11795 16243
rect 11829 16209 11863 16243
rect 11897 16209 11931 16243
rect 11965 16209 11999 16243
rect 12033 16209 12067 16243
rect 12101 16209 12135 16243
rect 12169 16209 12203 16243
rect 12237 16209 12271 16243
rect 12305 16209 12339 16243
rect 12373 16209 12407 16243
rect 12441 16209 12475 16243
rect 12509 16209 12543 16243
rect 12577 16209 12611 16243
rect 12645 16209 12679 16243
rect 12713 16209 12747 16243
rect 12781 16209 12815 16243
rect 12849 16209 12883 16243
rect 12917 16209 12951 16243
rect 12985 16209 13019 16243
rect 13053 16209 13087 16243
rect 13121 16209 13155 16243
rect 13189 16209 13223 16243
rect 13257 16209 13331 16243
rect 2595 16193 13331 16209
rect 2872 13324 13118 13340
rect 2872 13290 2888 13324
rect 2922 13290 2957 13324
rect 2991 13290 3026 13324
rect 3060 13290 3095 13324
rect 3129 13290 3164 13324
rect 3198 13290 3233 13324
rect 3267 13290 3302 13324
rect 3336 13290 3371 13324
rect 3405 13290 3440 13324
rect 3474 13290 3509 13324
rect 3543 13290 3578 13324
rect 3612 13290 3647 13324
rect 3681 13290 3716 13324
rect 3750 13290 3785 13324
rect 3819 13290 3854 13324
rect 3888 13290 3923 13324
rect 3957 13290 3992 13324
rect 4026 13290 4061 13324
rect 4095 13290 4130 13324
rect 4164 13290 4199 13324
rect 4233 13290 4268 13324
rect 4302 13290 4337 13324
rect 4371 13290 4406 13324
rect 4440 13290 4475 13324
rect 4509 13290 4544 13324
rect 4578 13290 4613 13324
rect 4647 13290 4682 13324
rect 4716 13290 4751 13324
rect 4785 13290 4820 13324
rect 4854 13290 4889 13324
rect 4923 13290 4958 13324
rect 4992 13290 5027 13324
rect 5061 13290 5096 13324
rect 5130 13290 5165 13324
rect 5199 13290 5234 13324
rect 5268 13290 5303 13324
rect 5337 13290 5372 13324
rect 5406 13290 5441 13324
rect 5475 13290 5510 13324
rect 5544 13290 5579 13324
rect 5613 13290 5648 13324
rect 5682 13290 5717 13324
rect 5751 13290 5786 13324
rect 5820 13290 5855 13324
rect 5889 13290 5924 13324
rect 5958 13290 5993 13324
rect 6027 13290 6062 13324
rect 6096 13290 6131 13324
rect 6165 13290 6200 13324
rect 6234 13290 6268 13324
rect 6302 13290 6336 13324
rect 6370 13290 6404 13324
rect 6438 13290 6472 13324
rect 6506 13290 6540 13324
rect 6574 13290 6608 13324
rect 6642 13290 6676 13324
rect 6710 13290 6744 13324
rect 6778 13290 6812 13324
rect 6846 13290 6880 13324
rect 6914 13290 6948 13324
rect 6982 13290 7016 13324
rect 7050 13290 7084 13324
rect 7118 13290 7152 13324
rect 7186 13290 7220 13324
rect 7254 13290 7288 13324
rect 7322 13290 7356 13324
rect 7390 13290 7424 13324
rect 7458 13290 7492 13324
rect 7526 13290 7560 13324
rect 7594 13290 7628 13324
rect 7662 13290 7696 13324
rect 7730 13290 7764 13324
rect 7798 13290 7832 13324
rect 7866 13290 7900 13324
rect 7934 13290 7968 13324
rect 8002 13290 8036 13324
rect 8070 13290 8104 13324
rect 8138 13290 8172 13324
rect 8206 13290 8240 13324
rect 8274 13290 8308 13324
rect 8342 13290 8376 13324
rect 8410 13290 8444 13324
rect 8478 13290 8512 13324
rect 8546 13290 8580 13324
rect 8614 13290 8648 13324
rect 8682 13290 8716 13324
rect 8750 13290 8784 13324
rect 8818 13290 8852 13324
rect 8886 13290 8920 13324
rect 8954 13290 8988 13324
rect 9022 13290 9056 13324
rect 9090 13290 9124 13324
rect 9158 13290 9192 13324
rect 9226 13290 9260 13324
rect 9294 13290 9328 13324
rect 9362 13290 9396 13324
rect 9430 13290 9464 13324
rect 9498 13290 9532 13324
rect 9566 13290 9600 13324
rect 9634 13290 9668 13324
rect 9702 13290 9736 13324
rect 9770 13290 9804 13324
rect 9838 13290 9872 13324
rect 9906 13290 9940 13324
rect 9974 13290 10008 13324
rect 10042 13290 10076 13324
rect 10110 13290 10144 13324
rect 10178 13290 10212 13324
rect 10246 13290 10280 13324
rect 10314 13290 10348 13324
rect 10382 13290 10416 13324
rect 10450 13290 10484 13324
rect 10518 13290 10552 13324
rect 10586 13290 10620 13324
rect 10654 13290 10688 13324
rect 10722 13290 10756 13324
rect 10790 13290 10824 13324
rect 10858 13290 10892 13324
rect 10926 13290 10960 13324
rect 10994 13290 11028 13324
rect 11062 13290 11096 13324
rect 11130 13290 11164 13324
rect 11198 13290 11232 13324
rect 11266 13290 11300 13324
rect 11334 13290 11368 13324
rect 11402 13290 11436 13324
rect 11470 13290 11504 13324
rect 11538 13290 11572 13324
rect 11606 13290 11640 13324
rect 11674 13290 11708 13324
rect 11742 13290 11776 13324
rect 11810 13290 11844 13324
rect 11878 13290 11912 13324
rect 11946 13290 11980 13324
rect 12014 13290 12048 13324
rect 12082 13290 12116 13324
rect 12150 13290 12184 13324
rect 12218 13290 12252 13324
rect 12286 13290 12320 13324
rect 12354 13290 12388 13324
rect 12422 13290 12456 13324
rect 12490 13290 12524 13324
rect 12558 13290 12592 13324
rect 12626 13290 12660 13324
rect 12694 13290 12728 13324
rect 12762 13290 12796 13324
rect 12830 13290 12864 13324
rect 12898 13290 12932 13324
rect 12966 13290 13000 13324
rect 13034 13290 13068 13324
rect 13102 13290 13118 13324
rect 2872 13274 13118 13290
rect 2872 12870 2908 13274
rect 3110 12870 3146 13274
rect 3426 12870 3462 13274
rect 3666 12870 3702 13274
rect 3980 12870 4016 13274
rect 4218 12870 4254 13274
rect 4534 12870 4570 13274
rect 4772 12870 4808 13274
rect 5088 12870 5124 13274
rect 5326 12870 5362 13274
rect 5642 12870 5678 13274
rect 5880 12870 5916 13274
rect 6196 12870 6232 13274
rect 6434 12870 6470 13274
rect 6750 12870 6786 13274
rect 6988 12870 7024 13274
rect 7304 12870 7340 13274
rect 7542 12870 7578 13274
rect 7858 12870 7894 13274
rect 8096 12870 8132 13274
rect 8412 12870 8448 13274
rect 8650 12870 8686 13274
rect 8966 12870 9002 13274
rect 9204 12870 9240 13274
rect 9520 12870 9556 13274
rect 9758 12870 9794 13274
rect 10074 12870 10110 13274
rect 10312 12870 10348 13274
rect 10628 12870 10664 13274
rect 10866 12870 10902 13274
rect 11182 12870 11218 13274
rect 11420 12870 11456 13274
rect 11736 12870 11772 13274
rect 11974 12870 12010 13274
rect 12290 12870 12326 13274
rect 12528 12870 12564 13274
rect 12844 12870 12880 13274
rect 13082 12870 13118 13274
rect 2872 12854 13118 12870
rect 2872 12820 2888 12854
rect 2922 12820 2957 12854
rect 2991 12820 3026 12854
rect 3060 12820 3095 12854
rect 3129 12820 3164 12854
rect 3198 12820 3233 12854
rect 3267 12820 3302 12854
rect 3336 12820 3371 12854
rect 3405 12820 3440 12854
rect 3474 12820 3509 12854
rect 3543 12820 3578 12854
rect 3612 12820 3647 12854
rect 3681 12820 3716 12854
rect 3750 12820 3785 12854
rect 3819 12820 3854 12854
rect 3888 12820 3923 12854
rect 3957 12820 3992 12854
rect 4026 12820 4061 12854
rect 4095 12820 4130 12854
rect 4164 12820 4199 12854
rect 4233 12820 4268 12854
rect 4302 12820 4337 12854
rect 4371 12820 4406 12854
rect 4440 12820 4475 12854
rect 4509 12820 4544 12854
rect 4578 12820 4613 12854
rect 4647 12820 4682 12854
rect 4716 12820 4751 12854
rect 4785 12820 4820 12854
rect 4854 12820 4889 12854
rect 4923 12820 4958 12854
rect 4992 12820 5027 12854
rect 5061 12820 5096 12854
rect 5130 12820 5165 12854
rect 5199 12820 5234 12854
rect 5268 12820 5303 12854
rect 5337 12820 5372 12854
rect 5406 12820 5441 12854
rect 5475 12820 5510 12854
rect 5544 12820 5579 12854
rect 5613 12820 5648 12854
rect 5682 12820 5717 12854
rect 5751 12820 5786 12854
rect 5820 12820 5855 12854
rect 5889 12820 5924 12854
rect 5958 12820 5993 12854
rect 6027 12820 6062 12854
rect 6096 12820 6131 12854
rect 6165 12820 6200 12854
rect 6234 12820 6268 12854
rect 6302 12820 6336 12854
rect 6370 12820 6404 12854
rect 6438 12820 6472 12854
rect 6506 12820 6540 12854
rect 6574 12820 6608 12854
rect 6642 12820 6676 12854
rect 6710 12820 6744 12854
rect 6778 12820 6812 12854
rect 6846 12820 6880 12854
rect 6914 12820 6948 12854
rect 6982 12820 7016 12854
rect 7050 12820 7084 12854
rect 7118 12820 7152 12854
rect 7186 12820 7220 12854
rect 7254 12820 7288 12854
rect 7322 12820 7356 12854
rect 7390 12820 7424 12854
rect 7458 12820 7492 12854
rect 7526 12820 7560 12854
rect 7594 12820 7628 12854
rect 7662 12820 7696 12854
rect 7730 12820 7764 12854
rect 7798 12820 7832 12854
rect 7866 12820 7900 12854
rect 7934 12820 7968 12854
rect 8002 12820 8036 12854
rect 8070 12820 8104 12854
rect 8138 12820 8172 12854
rect 8206 12820 8240 12854
rect 8274 12820 8308 12854
rect 8342 12820 8376 12854
rect 8410 12820 8444 12854
rect 8478 12820 8512 12854
rect 8546 12820 8580 12854
rect 8614 12820 8648 12854
rect 8682 12820 8716 12854
rect 8750 12820 8784 12854
rect 8818 12820 8852 12854
rect 8886 12820 8920 12854
rect 8954 12820 8988 12854
rect 9022 12820 9056 12854
rect 9090 12820 9124 12854
rect 9158 12820 9192 12854
rect 9226 12820 9260 12854
rect 9294 12820 9328 12854
rect 9362 12820 9396 12854
rect 9430 12820 9464 12854
rect 9498 12820 9532 12854
rect 9566 12820 9600 12854
rect 9634 12820 9668 12854
rect 9702 12820 9736 12854
rect 9770 12820 9804 12854
rect 9838 12820 9872 12854
rect 9906 12820 9940 12854
rect 9974 12820 10008 12854
rect 10042 12820 10076 12854
rect 10110 12820 10144 12854
rect 10178 12820 10212 12854
rect 10246 12820 10280 12854
rect 10314 12820 10348 12854
rect 10382 12820 10416 12854
rect 10450 12820 10484 12854
rect 10518 12820 10552 12854
rect 10586 12820 10620 12854
rect 10654 12820 10688 12854
rect 10722 12820 10756 12854
rect 10790 12820 10824 12854
rect 10858 12820 10892 12854
rect 10926 12820 10960 12854
rect 10994 12820 11028 12854
rect 11062 12820 11096 12854
rect 11130 12820 11164 12854
rect 11198 12820 11232 12854
rect 11266 12820 11300 12854
rect 11334 12820 11368 12854
rect 11402 12820 11436 12854
rect 11470 12820 11504 12854
rect 11538 12820 11572 12854
rect 11606 12820 11640 12854
rect 11674 12820 11708 12854
rect 11742 12820 11776 12854
rect 11810 12820 11844 12854
rect 11878 12820 11912 12854
rect 11946 12820 11980 12854
rect 12014 12820 12048 12854
rect 12082 12820 12116 12854
rect 12150 12820 12184 12854
rect 12218 12820 12252 12854
rect 12286 12820 12320 12854
rect 12354 12820 12388 12854
rect 12422 12820 12456 12854
rect 12490 12820 12524 12854
rect 12558 12820 12592 12854
rect 12626 12820 12660 12854
rect 12694 12820 12728 12854
rect 12762 12820 12796 12854
rect 12830 12820 12864 12854
rect 12898 12820 12932 12854
rect 12966 12820 13000 12854
rect 13034 12820 13068 12854
rect 13102 12820 13118 12854
rect 2872 12804 13118 12820
rect 5088 12800 5124 12804
rect 5326 12800 5362 12804
rect 5642 12800 5678 12804
rect 5880 12800 5916 12804
rect 6196 12800 6232 12804
rect 6434 12800 6470 12804
rect 6750 12800 6786 12804
rect 2872 11340 2908 11347
rect 3110 11340 3146 11347
rect 3426 11340 3462 11347
rect 3664 11340 3700 11347
rect 3980 11340 4016 11347
rect 4218 11340 4254 11347
rect 4534 11340 4570 11347
rect 4772 11340 4808 11347
rect 2872 11324 13118 11340
rect 2872 11290 2888 11324
rect 2922 11290 2957 11324
rect 2991 11290 3026 11324
rect 3060 11290 3095 11324
rect 3129 11290 3164 11324
rect 3198 11290 3233 11324
rect 3267 11290 3302 11324
rect 3336 11290 3371 11324
rect 3405 11290 3440 11324
rect 3474 11290 3509 11324
rect 3543 11290 3578 11324
rect 3612 11290 3647 11324
rect 3681 11290 3716 11324
rect 3750 11290 3785 11324
rect 3819 11290 3854 11324
rect 3888 11290 3923 11324
rect 3957 11290 3992 11324
rect 4026 11290 4061 11324
rect 4095 11290 4130 11324
rect 4164 11290 4199 11324
rect 4233 11290 4268 11324
rect 4302 11290 4337 11324
rect 4371 11290 4406 11324
rect 4440 11290 4475 11324
rect 4509 11290 4544 11324
rect 4578 11290 4613 11324
rect 4647 11290 4682 11324
rect 4716 11290 4751 11324
rect 4785 11290 4820 11324
rect 4854 11290 4889 11324
rect 4923 11290 4958 11324
rect 4992 11290 5027 11324
rect 5061 11290 5096 11324
rect 5130 11290 5165 11324
rect 5199 11290 5234 11324
rect 5268 11290 5303 11324
rect 5337 11290 5372 11324
rect 5406 11290 5441 11324
rect 5475 11290 5510 11324
rect 5544 11290 5579 11324
rect 5613 11290 5648 11324
rect 5682 11290 5717 11324
rect 5751 11290 5786 11324
rect 5820 11290 5855 11324
rect 5889 11290 5924 11324
rect 5958 11290 5993 11324
rect 6027 11290 6062 11324
rect 6096 11290 6131 11324
rect 6165 11290 6200 11324
rect 6234 11290 6268 11324
rect 6302 11290 6336 11324
rect 6370 11290 6404 11324
rect 6438 11290 6472 11324
rect 6506 11290 6540 11324
rect 6574 11290 6608 11324
rect 6642 11290 6676 11324
rect 6710 11290 6744 11324
rect 6778 11290 6812 11324
rect 6846 11290 6880 11324
rect 6914 11290 6948 11324
rect 6982 11290 7016 11324
rect 7050 11290 7084 11324
rect 7118 11290 7152 11324
rect 7186 11290 7220 11324
rect 7254 11290 7288 11324
rect 7322 11290 7356 11324
rect 7390 11290 7424 11324
rect 7458 11290 7492 11324
rect 7526 11290 7560 11324
rect 7594 11290 7628 11324
rect 7662 11290 7696 11324
rect 7730 11290 7764 11324
rect 7798 11290 7832 11324
rect 7866 11290 7900 11324
rect 7934 11290 7968 11324
rect 8002 11290 8036 11324
rect 8070 11290 8104 11324
rect 8138 11290 8172 11324
rect 8206 11290 8240 11324
rect 8274 11290 8308 11324
rect 8342 11290 8376 11324
rect 8410 11290 8444 11324
rect 8478 11290 8512 11324
rect 8546 11290 8580 11324
rect 8614 11290 8648 11324
rect 8682 11290 8716 11324
rect 8750 11290 8784 11324
rect 8818 11290 8852 11324
rect 8886 11290 8920 11324
rect 8954 11290 8988 11324
rect 9022 11290 9056 11324
rect 9090 11290 9124 11324
rect 9158 11290 9192 11324
rect 9226 11290 9260 11324
rect 9294 11290 9328 11324
rect 9362 11290 9396 11324
rect 9430 11290 9464 11324
rect 9498 11290 9532 11324
rect 9566 11290 9600 11324
rect 9634 11290 9668 11324
rect 9702 11290 9736 11324
rect 9770 11290 9804 11324
rect 9838 11290 9872 11324
rect 9906 11290 9940 11324
rect 9974 11290 10008 11324
rect 10042 11290 10076 11324
rect 10110 11290 10144 11324
rect 10178 11290 10212 11324
rect 10246 11290 10280 11324
rect 10314 11290 10348 11324
rect 10382 11290 10416 11324
rect 10450 11290 10484 11324
rect 10518 11290 10552 11324
rect 10586 11290 10620 11324
rect 10654 11290 10688 11324
rect 10722 11290 10756 11324
rect 10790 11290 10824 11324
rect 10858 11290 10892 11324
rect 10926 11290 10960 11324
rect 10994 11290 11028 11324
rect 11062 11290 11096 11324
rect 11130 11290 11164 11324
rect 11198 11290 11232 11324
rect 11266 11290 11300 11324
rect 11334 11290 11368 11324
rect 11402 11290 11436 11324
rect 11470 11290 11504 11324
rect 11538 11290 11572 11324
rect 11606 11290 11640 11324
rect 11674 11290 11708 11324
rect 11742 11290 11776 11324
rect 11810 11290 11844 11324
rect 11878 11290 11912 11324
rect 11946 11290 11980 11324
rect 12014 11290 12048 11324
rect 12082 11290 12116 11324
rect 12150 11290 12184 11324
rect 12218 11290 12252 11324
rect 12286 11290 12320 11324
rect 12354 11290 12388 11324
rect 12422 11290 12456 11324
rect 12490 11290 12524 11324
rect 12558 11290 12592 11324
rect 12626 11290 12660 11324
rect 12694 11290 12728 11324
rect 12762 11290 12796 11324
rect 12830 11290 12864 11324
rect 12898 11290 12932 11324
rect 12966 11290 13000 11324
rect 13034 11290 13068 11324
rect 13102 11290 13118 11324
rect 2872 11274 13118 11290
rect 2872 10870 2908 11274
rect 3110 10870 3146 11274
rect 3426 10870 3462 11274
rect 3664 10870 3700 11274
rect 3980 10870 4016 11274
rect 4218 10870 4254 11274
rect 4534 10870 4570 11274
rect 4772 10870 4808 11274
rect 5088 10870 5124 11274
rect 5326 10870 5362 11274
rect 5642 10870 5678 11274
rect 5880 10870 5916 11274
rect 6196 10870 6232 11274
rect 6434 10870 6470 11274
rect 6750 10870 6786 11274
rect 6988 10870 7024 11274
rect 7304 10870 7340 11274
rect 7542 10870 7578 11274
rect 7858 10870 7894 11274
rect 8096 10870 8132 11274
rect 8412 10870 8448 11274
rect 8650 10870 8686 11274
rect 8966 10870 9002 11274
rect 9204 10870 9240 11274
rect 9520 10870 9556 11274
rect 9758 10870 9794 11274
rect 10074 10870 10110 11274
rect 10312 10870 10348 11274
rect 10628 10870 10664 11274
rect 10866 10870 10902 11274
rect 11182 10870 11218 11274
rect 11420 10870 11456 11274
rect 11736 10870 11772 11274
rect 11974 10870 12010 11274
rect 12290 10870 12326 11274
rect 12528 10870 12564 11274
rect 12844 10870 12880 11274
rect 13082 10870 13118 11274
rect 2872 10854 13118 10870
rect 2872 10820 2888 10854
rect 2922 10820 2957 10854
rect 2991 10820 3026 10854
rect 3060 10820 3095 10854
rect 3129 10820 3164 10854
rect 3198 10820 3233 10854
rect 3267 10820 3302 10854
rect 3336 10820 3371 10854
rect 3405 10820 3440 10854
rect 3474 10820 3509 10854
rect 3543 10820 3578 10854
rect 3612 10820 3647 10854
rect 3681 10820 3716 10854
rect 3750 10820 3785 10854
rect 3819 10820 3854 10854
rect 3888 10820 3923 10854
rect 3957 10820 3992 10854
rect 4026 10820 4061 10854
rect 4095 10820 4130 10854
rect 4164 10820 4199 10854
rect 4233 10820 4268 10854
rect 4302 10820 4337 10854
rect 4371 10820 4406 10854
rect 4440 10820 4475 10854
rect 4509 10820 4544 10854
rect 4578 10820 4613 10854
rect 4647 10820 4682 10854
rect 4716 10820 4751 10854
rect 4785 10820 4820 10854
rect 4854 10820 4889 10854
rect 4923 10820 4958 10854
rect 4992 10820 5027 10854
rect 5061 10820 5096 10854
rect 5130 10820 5165 10854
rect 5199 10820 5234 10854
rect 5268 10820 5303 10854
rect 5337 10820 5372 10854
rect 5406 10820 5441 10854
rect 5475 10820 5510 10854
rect 5544 10820 5579 10854
rect 5613 10820 5648 10854
rect 5682 10820 5717 10854
rect 5751 10820 5786 10854
rect 5820 10820 5855 10854
rect 5889 10820 5924 10854
rect 5958 10820 5993 10854
rect 6027 10820 6062 10854
rect 6096 10820 6131 10854
rect 6165 10820 6200 10854
rect 6234 10820 6268 10854
rect 6302 10820 6336 10854
rect 6370 10820 6404 10854
rect 6438 10820 6472 10854
rect 6506 10820 6540 10854
rect 6574 10820 6608 10854
rect 6642 10820 6676 10854
rect 6710 10820 6744 10854
rect 6778 10820 6812 10854
rect 6846 10820 6880 10854
rect 6914 10820 6948 10854
rect 6982 10820 7016 10854
rect 7050 10820 7084 10854
rect 7118 10820 7152 10854
rect 7186 10820 7220 10854
rect 7254 10820 7288 10854
rect 7322 10820 7356 10854
rect 7390 10820 7424 10854
rect 7458 10820 7492 10854
rect 7526 10820 7560 10854
rect 7594 10820 7628 10854
rect 7662 10820 7696 10854
rect 7730 10820 7764 10854
rect 7798 10820 7832 10854
rect 7866 10820 7900 10854
rect 7934 10820 7968 10854
rect 8002 10820 8036 10854
rect 8070 10820 8104 10854
rect 8138 10820 8172 10854
rect 8206 10820 8240 10854
rect 8274 10820 8308 10854
rect 8342 10820 8376 10854
rect 8410 10820 8444 10854
rect 8478 10820 8512 10854
rect 8546 10820 8580 10854
rect 8614 10820 8648 10854
rect 8682 10820 8716 10854
rect 8750 10820 8784 10854
rect 8818 10820 8852 10854
rect 8886 10820 8920 10854
rect 8954 10820 8988 10854
rect 9022 10820 9056 10854
rect 9090 10820 9124 10854
rect 9158 10820 9192 10854
rect 9226 10820 9260 10854
rect 9294 10820 9328 10854
rect 9362 10820 9396 10854
rect 9430 10820 9464 10854
rect 9498 10820 9532 10854
rect 9566 10820 9600 10854
rect 9634 10820 9668 10854
rect 9702 10820 9736 10854
rect 9770 10820 9804 10854
rect 9838 10820 9872 10854
rect 9906 10820 9940 10854
rect 9974 10820 10008 10854
rect 10042 10820 10076 10854
rect 10110 10820 10144 10854
rect 10178 10820 10212 10854
rect 10246 10820 10280 10854
rect 10314 10820 10348 10854
rect 10382 10820 10416 10854
rect 10450 10820 10484 10854
rect 10518 10820 10552 10854
rect 10586 10820 10620 10854
rect 10654 10820 10688 10854
rect 10722 10820 10756 10854
rect 10790 10820 10824 10854
rect 10858 10820 10892 10854
rect 10926 10820 10960 10854
rect 10994 10820 11028 10854
rect 11062 10820 11096 10854
rect 11130 10820 11164 10854
rect 11198 10820 11232 10854
rect 11266 10820 11300 10854
rect 11334 10820 11368 10854
rect 11402 10820 11436 10854
rect 11470 10820 11504 10854
rect 11538 10820 11572 10854
rect 11606 10820 11640 10854
rect 11674 10820 11708 10854
rect 11742 10820 11776 10854
rect 11810 10820 11844 10854
rect 11878 10820 11912 10854
rect 11946 10820 11980 10854
rect 12014 10820 12048 10854
rect 12082 10820 12116 10854
rect 12150 10820 12184 10854
rect 12218 10820 12252 10854
rect 12286 10820 12320 10854
rect 12354 10820 12388 10854
rect 12422 10820 12456 10854
rect 12490 10820 12524 10854
rect 12558 10820 12592 10854
rect 12626 10820 12660 10854
rect 12694 10820 12728 10854
rect 12762 10820 12796 10854
rect 12830 10820 12864 10854
rect 12898 10820 12932 10854
rect 12966 10820 13000 10854
rect 13034 10820 13068 10854
rect 13102 10820 13118 10854
rect 2872 10804 13118 10820
rect 2872 9324 13118 9340
rect 2872 9290 2888 9324
rect 2922 9290 2957 9324
rect 2991 9290 3026 9324
rect 3060 9290 3095 9324
rect 3129 9290 3164 9324
rect 3198 9290 3233 9324
rect 3267 9290 3302 9324
rect 3336 9290 3371 9324
rect 3405 9290 3440 9324
rect 3474 9290 3509 9324
rect 3543 9290 3578 9324
rect 3612 9290 3647 9324
rect 3681 9290 3716 9324
rect 3750 9290 3785 9324
rect 3819 9290 3854 9324
rect 3888 9290 3923 9324
rect 3957 9290 3992 9324
rect 4026 9290 4061 9324
rect 4095 9290 4130 9324
rect 4164 9290 4199 9324
rect 4233 9290 4268 9324
rect 4302 9290 4337 9324
rect 4371 9290 4406 9324
rect 4440 9290 4475 9324
rect 4509 9290 4544 9324
rect 4578 9290 4613 9324
rect 4647 9290 4682 9324
rect 4716 9290 4751 9324
rect 4785 9290 4820 9324
rect 4854 9290 4889 9324
rect 4923 9290 4958 9324
rect 4992 9290 5027 9324
rect 5061 9290 5096 9324
rect 5130 9290 5165 9324
rect 5199 9290 5234 9324
rect 5268 9290 5303 9324
rect 5337 9290 5372 9324
rect 5406 9290 5441 9324
rect 5475 9290 5510 9324
rect 5544 9290 5579 9324
rect 5613 9290 5648 9324
rect 5682 9290 5717 9324
rect 5751 9290 5786 9324
rect 5820 9290 5855 9324
rect 5889 9290 5924 9324
rect 5958 9290 5993 9324
rect 6027 9290 6062 9324
rect 6096 9290 6131 9324
rect 6165 9290 6200 9324
rect 6234 9290 6268 9324
rect 6302 9290 6336 9324
rect 6370 9290 6404 9324
rect 6438 9290 6472 9324
rect 6506 9290 6540 9324
rect 6574 9290 6608 9324
rect 6642 9290 6676 9324
rect 6710 9290 6744 9324
rect 6778 9290 6812 9324
rect 6846 9290 6880 9324
rect 6914 9290 6948 9324
rect 6982 9290 7016 9324
rect 7050 9290 7084 9324
rect 7118 9290 7152 9324
rect 7186 9290 7220 9324
rect 7254 9290 7288 9324
rect 7322 9290 7356 9324
rect 7390 9290 7424 9324
rect 7458 9290 7492 9324
rect 7526 9290 7560 9324
rect 7594 9290 7628 9324
rect 7662 9290 7696 9324
rect 7730 9290 7764 9324
rect 7798 9290 7832 9324
rect 7866 9290 7900 9324
rect 7934 9290 7968 9324
rect 8002 9290 8036 9324
rect 8070 9290 8104 9324
rect 8138 9290 8172 9324
rect 8206 9290 8240 9324
rect 8274 9290 8308 9324
rect 8342 9290 8376 9324
rect 8410 9290 8444 9324
rect 8478 9290 8512 9324
rect 8546 9290 8580 9324
rect 8614 9290 8648 9324
rect 8682 9290 8716 9324
rect 8750 9290 8784 9324
rect 8818 9290 8852 9324
rect 8886 9290 8920 9324
rect 8954 9290 8988 9324
rect 9022 9290 9056 9324
rect 9090 9290 9124 9324
rect 9158 9290 9192 9324
rect 9226 9290 9260 9324
rect 9294 9290 9328 9324
rect 9362 9290 9396 9324
rect 9430 9290 9464 9324
rect 9498 9290 9532 9324
rect 9566 9290 9600 9324
rect 9634 9290 9668 9324
rect 9702 9290 9736 9324
rect 9770 9290 9804 9324
rect 9838 9290 9872 9324
rect 9906 9290 9940 9324
rect 9974 9290 10008 9324
rect 10042 9290 10076 9324
rect 10110 9290 10144 9324
rect 10178 9290 10212 9324
rect 10246 9290 10280 9324
rect 10314 9290 10348 9324
rect 10382 9290 10416 9324
rect 10450 9290 10484 9324
rect 10518 9290 10552 9324
rect 10586 9290 10620 9324
rect 10654 9290 10688 9324
rect 10722 9290 10756 9324
rect 10790 9290 10824 9324
rect 10858 9290 10892 9324
rect 10926 9290 10960 9324
rect 10994 9290 11028 9324
rect 11062 9290 11096 9324
rect 11130 9290 11164 9324
rect 11198 9290 11232 9324
rect 11266 9290 11300 9324
rect 11334 9290 11368 9324
rect 11402 9290 11436 9324
rect 11470 9290 11504 9324
rect 11538 9290 11572 9324
rect 11606 9290 11640 9324
rect 11674 9290 11708 9324
rect 11742 9290 11776 9324
rect 11810 9290 11844 9324
rect 11878 9290 11912 9324
rect 11946 9290 11980 9324
rect 12014 9290 12048 9324
rect 12082 9290 12116 9324
rect 12150 9290 12184 9324
rect 12218 9290 12252 9324
rect 12286 9290 12320 9324
rect 12354 9290 12388 9324
rect 12422 9290 12456 9324
rect 12490 9290 12524 9324
rect 12558 9290 12592 9324
rect 12626 9290 12660 9324
rect 12694 9290 12728 9324
rect 12762 9290 12796 9324
rect 12830 9290 12864 9324
rect 12898 9290 12932 9324
rect 12966 9290 13000 9324
rect 13034 9290 13068 9324
rect 13102 9290 13118 9324
rect 2872 9274 13118 9290
rect 2872 8870 2908 9274
rect 3110 8870 3146 9274
rect 3426 8870 3462 9274
rect 3666 8870 3702 9274
rect 3980 8870 4016 9274
rect 4218 8870 4254 9274
rect 4534 8870 4570 9274
rect 4772 8870 4808 9274
rect 5088 8870 5124 9274
rect 5326 8870 5362 9274
rect 5642 8870 5678 9274
rect 5880 8870 5916 9274
rect 6196 8870 6232 9274
rect 6434 8870 6470 9274
rect 6750 8870 6786 9274
rect 6988 8870 7024 9274
rect 7304 8870 7340 9274
rect 7542 8870 7578 9274
rect 7858 8870 7894 9274
rect 8096 8870 8132 9274
rect 8412 8870 8448 9274
rect 8650 8870 8686 9274
rect 8966 8870 9002 9274
rect 9204 8870 9240 9274
rect 9520 8870 9556 9274
rect 9758 8870 9794 9274
rect 10074 8870 10110 9274
rect 10312 8870 10348 9274
rect 10628 8870 10664 9274
rect 10866 8870 10902 9274
rect 11182 8870 11218 9274
rect 11420 8870 11456 9274
rect 11736 8870 11772 9274
rect 11974 8870 12010 9274
rect 12290 8870 12326 9274
rect 12528 8870 12564 9274
rect 12844 8870 12880 9274
rect 13082 8870 13118 9274
rect 2872 8854 13118 8870
rect 2872 8820 2888 8854
rect 2922 8820 2957 8854
rect 2991 8820 3026 8854
rect 3060 8820 3095 8854
rect 3129 8820 3164 8854
rect 3198 8820 3233 8854
rect 3267 8820 3302 8854
rect 3336 8820 3371 8854
rect 3405 8820 3440 8854
rect 3474 8820 3509 8854
rect 3543 8820 3578 8854
rect 3612 8820 3647 8854
rect 3681 8820 3716 8854
rect 3750 8820 3785 8854
rect 3819 8820 3854 8854
rect 3888 8820 3923 8854
rect 3957 8820 3992 8854
rect 4026 8820 4061 8854
rect 4095 8820 4130 8854
rect 4164 8820 4199 8854
rect 4233 8820 4268 8854
rect 4302 8820 4337 8854
rect 4371 8820 4406 8854
rect 4440 8820 4475 8854
rect 4509 8820 4544 8854
rect 4578 8820 4613 8854
rect 4647 8820 4682 8854
rect 4716 8820 4751 8854
rect 4785 8820 4820 8854
rect 4854 8820 4889 8854
rect 4923 8820 4958 8854
rect 4992 8820 5027 8854
rect 5061 8820 5096 8854
rect 5130 8820 5165 8854
rect 5199 8820 5234 8854
rect 5268 8820 5303 8854
rect 5337 8820 5372 8854
rect 5406 8820 5441 8854
rect 5475 8820 5510 8854
rect 5544 8820 5579 8854
rect 5613 8820 5648 8854
rect 5682 8820 5717 8854
rect 5751 8820 5786 8854
rect 5820 8820 5855 8854
rect 5889 8820 5924 8854
rect 5958 8820 5993 8854
rect 6027 8820 6062 8854
rect 6096 8820 6131 8854
rect 6165 8820 6200 8854
rect 6234 8820 6268 8854
rect 6302 8820 6336 8854
rect 6370 8820 6404 8854
rect 6438 8820 6472 8854
rect 6506 8820 6540 8854
rect 6574 8820 6608 8854
rect 6642 8820 6676 8854
rect 6710 8820 6744 8854
rect 6778 8820 6812 8854
rect 6846 8820 6880 8854
rect 6914 8820 6948 8854
rect 6982 8820 7016 8854
rect 7050 8820 7084 8854
rect 7118 8820 7152 8854
rect 7186 8820 7220 8854
rect 7254 8820 7288 8854
rect 7322 8820 7356 8854
rect 7390 8820 7424 8854
rect 7458 8820 7492 8854
rect 7526 8820 7560 8854
rect 7594 8820 7628 8854
rect 7662 8820 7696 8854
rect 7730 8820 7764 8854
rect 7798 8820 7832 8854
rect 7866 8820 7900 8854
rect 7934 8820 7968 8854
rect 8002 8820 8036 8854
rect 8070 8820 8104 8854
rect 8138 8820 8172 8854
rect 8206 8820 8240 8854
rect 8274 8820 8308 8854
rect 8342 8820 8376 8854
rect 8410 8820 8444 8854
rect 8478 8820 8512 8854
rect 8546 8820 8580 8854
rect 8614 8820 8648 8854
rect 8682 8820 8716 8854
rect 8750 8820 8784 8854
rect 8818 8820 8852 8854
rect 8886 8820 8920 8854
rect 8954 8820 8988 8854
rect 9022 8820 9056 8854
rect 9090 8820 9124 8854
rect 9158 8820 9192 8854
rect 9226 8820 9260 8854
rect 9294 8820 9328 8854
rect 9362 8820 9396 8854
rect 9430 8820 9464 8854
rect 9498 8820 9532 8854
rect 9566 8820 9600 8854
rect 9634 8820 9668 8854
rect 9702 8820 9736 8854
rect 9770 8820 9804 8854
rect 9838 8820 9872 8854
rect 9906 8820 9940 8854
rect 9974 8820 10008 8854
rect 10042 8820 10076 8854
rect 10110 8820 10144 8854
rect 10178 8820 10212 8854
rect 10246 8820 10280 8854
rect 10314 8820 10348 8854
rect 10382 8820 10416 8854
rect 10450 8820 10484 8854
rect 10518 8820 10552 8854
rect 10586 8820 10620 8854
rect 10654 8820 10688 8854
rect 10722 8820 10756 8854
rect 10790 8820 10824 8854
rect 10858 8820 10892 8854
rect 10926 8820 10960 8854
rect 10994 8820 11028 8854
rect 11062 8820 11096 8854
rect 11130 8820 11164 8854
rect 11198 8820 11232 8854
rect 11266 8820 11300 8854
rect 11334 8820 11368 8854
rect 11402 8820 11436 8854
rect 11470 8820 11504 8854
rect 11538 8820 11572 8854
rect 11606 8820 11640 8854
rect 11674 8820 11708 8854
rect 11742 8820 11776 8854
rect 11810 8820 11844 8854
rect 11878 8820 11912 8854
rect 11946 8820 11980 8854
rect 12014 8820 12048 8854
rect 12082 8820 12116 8854
rect 12150 8820 12184 8854
rect 12218 8820 12252 8854
rect 12286 8820 12320 8854
rect 12354 8820 12388 8854
rect 12422 8820 12456 8854
rect 12490 8820 12524 8854
rect 12558 8820 12592 8854
rect 12626 8820 12660 8854
rect 12694 8820 12728 8854
rect 12762 8820 12796 8854
rect 12830 8820 12864 8854
rect 12898 8820 12932 8854
rect 12966 8820 13000 8854
rect 13034 8820 13068 8854
rect 13102 8820 13118 8854
rect 2872 8804 13118 8820
rect 5088 8800 5124 8804
rect 5326 8800 5362 8804
rect 5642 8800 5678 8804
rect 5880 8800 5916 8804
rect 6196 8800 6232 8804
rect 6434 8800 6470 8804
rect 6750 8800 6786 8804
rect 2872 7340 2908 7347
rect 3110 7340 3146 7347
rect 3426 7340 3462 7347
rect 3664 7340 3700 7347
rect 3980 7340 4016 7347
rect 4218 7340 4254 7347
rect 4534 7340 4570 7347
rect 4772 7340 4808 7347
rect 2872 7324 13118 7340
rect 2872 7290 2888 7324
rect 2922 7290 2957 7324
rect 2991 7290 3026 7324
rect 3060 7290 3095 7324
rect 3129 7290 3164 7324
rect 3198 7290 3233 7324
rect 3267 7290 3302 7324
rect 3336 7290 3371 7324
rect 3405 7290 3440 7324
rect 3474 7290 3509 7324
rect 3543 7290 3578 7324
rect 3612 7290 3647 7324
rect 3681 7290 3716 7324
rect 3750 7290 3785 7324
rect 3819 7290 3854 7324
rect 3888 7290 3923 7324
rect 3957 7290 3992 7324
rect 4026 7290 4061 7324
rect 4095 7290 4130 7324
rect 4164 7290 4199 7324
rect 4233 7290 4268 7324
rect 4302 7290 4337 7324
rect 4371 7290 4406 7324
rect 4440 7290 4475 7324
rect 4509 7290 4544 7324
rect 4578 7290 4613 7324
rect 4647 7290 4682 7324
rect 4716 7290 4751 7324
rect 4785 7290 4820 7324
rect 4854 7290 4889 7324
rect 4923 7290 4958 7324
rect 4992 7290 5027 7324
rect 5061 7290 5096 7324
rect 5130 7290 5165 7324
rect 5199 7290 5234 7324
rect 5268 7290 5303 7324
rect 5337 7290 5372 7324
rect 5406 7290 5441 7324
rect 5475 7290 5510 7324
rect 5544 7290 5579 7324
rect 5613 7290 5648 7324
rect 5682 7290 5717 7324
rect 5751 7290 5786 7324
rect 5820 7290 5855 7324
rect 5889 7290 5924 7324
rect 5958 7290 5993 7324
rect 6027 7290 6062 7324
rect 6096 7290 6131 7324
rect 6165 7290 6200 7324
rect 6234 7290 6268 7324
rect 6302 7290 6336 7324
rect 6370 7290 6404 7324
rect 6438 7290 6472 7324
rect 6506 7290 6540 7324
rect 6574 7290 6608 7324
rect 6642 7290 6676 7324
rect 6710 7290 6744 7324
rect 6778 7290 6812 7324
rect 6846 7290 6880 7324
rect 6914 7290 6948 7324
rect 6982 7290 7016 7324
rect 7050 7290 7084 7324
rect 7118 7290 7152 7324
rect 7186 7290 7220 7324
rect 7254 7290 7288 7324
rect 7322 7290 7356 7324
rect 7390 7290 7424 7324
rect 7458 7290 7492 7324
rect 7526 7290 7560 7324
rect 7594 7290 7628 7324
rect 7662 7290 7696 7324
rect 7730 7290 7764 7324
rect 7798 7290 7832 7324
rect 7866 7290 7900 7324
rect 7934 7290 7968 7324
rect 8002 7290 8036 7324
rect 8070 7290 8104 7324
rect 8138 7290 8172 7324
rect 8206 7290 8240 7324
rect 8274 7290 8308 7324
rect 8342 7290 8376 7324
rect 8410 7290 8444 7324
rect 8478 7290 8512 7324
rect 8546 7290 8580 7324
rect 8614 7290 8648 7324
rect 8682 7290 8716 7324
rect 8750 7290 8784 7324
rect 8818 7290 8852 7324
rect 8886 7290 8920 7324
rect 8954 7290 8988 7324
rect 9022 7290 9056 7324
rect 9090 7290 9124 7324
rect 9158 7290 9192 7324
rect 9226 7290 9260 7324
rect 9294 7290 9328 7324
rect 9362 7290 9396 7324
rect 9430 7290 9464 7324
rect 9498 7290 9532 7324
rect 9566 7290 9600 7324
rect 9634 7290 9668 7324
rect 9702 7290 9736 7324
rect 9770 7290 9804 7324
rect 9838 7290 9872 7324
rect 9906 7290 9940 7324
rect 9974 7290 10008 7324
rect 10042 7290 10076 7324
rect 10110 7290 10144 7324
rect 10178 7290 10212 7324
rect 10246 7290 10280 7324
rect 10314 7290 10348 7324
rect 10382 7290 10416 7324
rect 10450 7290 10484 7324
rect 10518 7290 10552 7324
rect 10586 7290 10620 7324
rect 10654 7290 10688 7324
rect 10722 7290 10756 7324
rect 10790 7290 10824 7324
rect 10858 7290 10892 7324
rect 10926 7290 10960 7324
rect 10994 7290 11028 7324
rect 11062 7290 11096 7324
rect 11130 7290 11164 7324
rect 11198 7290 11232 7324
rect 11266 7290 11300 7324
rect 11334 7290 11368 7324
rect 11402 7290 11436 7324
rect 11470 7290 11504 7324
rect 11538 7290 11572 7324
rect 11606 7290 11640 7324
rect 11674 7290 11708 7324
rect 11742 7290 11776 7324
rect 11810 7290 11844 7324
rect 11878 7290 11912 7324
rect 11946 7290 11980 7324
rect 12014 7290 12048 7324
rect 12082 7290 12116 7324
rect 12150 7290 12184 7324
rect 12218 7290 12252 7324
rect 12286 7290 12320 7324
rect 12354 7290 12388 7324
rect 12422 7290 12456 7324
rect 12490 7290 12524 7324
rect 12558 7290 12592 7324
rect 12626 7290 12660 7324
rect 12694 7290 12728 7324
rect 12762 7290 12796 7324
rect 12830 7290 12864 7324
rect 12898 7290 12932 7324
rect 12966 7290 13000 7324
rect 13034 7290 13068 7324
rect 13102 7290 13118 7324
rect 2872 7274 13118 7290
rect 2872 6870 2908 7274
rect 3110 6870 3146 7274
rect 3426 6870 3462 7274
rect 3664 6870 3700 7274
rect 3980 6870 4016 7274
rect 4218 6870 4254 7274
rect 4534 6870 4570 7274
rect 4772 6870 4808 7274
rect 5088 6870 5124 7274
rect 5326 6870 5362 7274
rect 5642 6870 5678 7274
rect 5880 6870 5916 7274
rect 6196 6870 6232 7274
rect 6434 6870 6470 7274
rect 6750 6870 6786 7274
rect 6988 6870 7024 7274
rect 7304 6870 7340 7274
rect 7542 6870 7578 7274
rect 7858 6870 7894 7274
rect 8096 6870 8132 7274
rect 8412 6870 8448 7274
rect 8650 6870 8686 7274
rect 8966 6870 9002 7274
rect 9204 6870 9240 7274
rect 9520 6870 9556 7274
rect 9758 6870 9794 7274
rect 10074 6870 10110 7274
rect 10312 6870 10348 7274
rect 10628 6870 10664 7274
rect 10866 6870 10902 7274
rect 11182 6870 11218 7274
rect 11420 6870 11456 7274
rect 11736 6870 11772 7274
rect 11974 6870 12010 7274
rect 12290 6870 12326 7274
rect 12528 6870 12564 7274
rect 12844 6870 12880 7274
rect 13082 6870 13118 7274
rect 2872 6854 13118 6870
rect 2872 6820 2888 6854
rect 2922 6820 2957 6854
rect 2991 6820 3026 6854
rect 3060 6820 3095 6854
rect 3129 6820 3164 6854
rect 3198 6820 3233 6854
rect 3267 6820 3302 6854
rect 3336 6820 3371 6854
rect 3405 6820 3440 6854
rect 3474 6820 3509 6854
rect 3543 6820 3578 6854
rect 3612 6820 3647 6854
rect 3681 6820 3716 6854
rect 3750 6820 3785 6854
rect 3819 6820 3854 6854
rect 3888 6820 3923 6854
rect 3957 6820 3992 6854
rect 4026 6820 4061 6854
rect 4095 6820 4130 6854
rect 4164 6820 4199 6854
rect 4233 6820 4268 6854
rect 4302 6820 4337 6854
rect 4371 6820 4406 6854
rect 4440 6820 4475 6854
rect 4509 6820 4544 6854
rect 4578 6820 4613 6854
rect 4647 6820 4682 6854
rect 4716 6820 4751 6854
rect 4785 6820 4820 6854
rect 4854 6820 4889 6854
rect 4923 6820 4958 6854
rect 4992 6820 5027 6854
rect 5061 6820 5096 6854
rect 5130 6820 5165 6854
rect 5199 6820 5234 6854
rect 5268 6820 5303 6854
rect 5337 6820 5372 6854
rect 5406 6820 5441 6854
rect 5475 6820 5510 6854
rect 5544 6820 5579 6854
rect 5613 6820 5648 6854
rect 5682 6820 5717 6854
rect 5751 6820 5786 6854
rect 5820 6820 5855 6854
rect 5889 6820 5924 6854
rect 5958 6820 5993 6854
rect 6027 6820 6062 6854
rect 6096 6820 6131 6854
rect 6165 6820 6200 6854
rect 6234 6820 6268 6854
rect 6302 6820 6336 6854
rect 6370 6820 6404 6854
rect 6438 6820 6472 6854
rect 6506 6820 6540 6854
rect 6574 6820 6608 6854
rect 6642 6820 6676 6854
rect 6710 6820 6744 6854
rect 6778 6820 6812 6854
rect 6846 6820 6880 6854
rect 6914 6820 6948 6854
rect 6982 6820 7016 6854
rect 7050 6820 7084 6854
rect 7118 6820 7152 6854
rect 7186 6820 7220 6854
rect 7254 6820 7288 6854
rect 7322 6820 7356 6854
rect 7390 6820 7424 6854
rect 7458 6820 7492 6854
rect 7526 6820 7560 6854
rect 7594 6820 7628 6854
rect 7662 6820 7696 6854
rect 7730 6820 7764 6854
rect 7798 6820 7832 6854
rect 7866 6820 7900 6854
rect 7934 6820 7968 6854
rect 8002 6820 8036 6854
rect 8070 6820 8104 6854
rect 8138 6820 8172 6854
rect 8206 6820 8240 6854
rect 8274 6820 8308 6854
rect 8342 6820 8376 6854
rect 8410 6820 8444 6854
rect 8478 6820 8512 6854
rect 8546 6820 8580 6854
rect 8614 6820 8648 6854
rect 8682 6820 8716 6854
rect 8750 6820 8784 6854
rect 8818 6820 8852 6854
rect 8886 6820 8920 6854
rect 8954 6820 8988 6854
rect 9022 6820 9056 6854
rect 9090 6820 9124 6854
rect 9158 6820 9192 6854
rect 9226 6820 9260 6854
rect 9294 6820 9328 6854
rect 9362 6820 9396 6854
rect 9430 6820 9464 6854
rect 9498 6820 9532 6854
rect 9566 6820 9600 6854
rect 9634 6820 9668 6854
rect 9702 6820 9736 6854
rect 9770 6820 9804 6854
rect 9838 6820 9872 6854
rect 9906 6820 9940 6854
rect 9974 6820 10008 6854
rect 10042 6820 10076 6854
rect 10110 6820 10144 6854
rect 10178 6820 10212 6854
rect 10246 6820 10280 6854
rect 10314 6820 10348 6854
rect 10382 6820 10416 6854
rect 10450 6820 10484 6854
rect 10518 6820 10552 6854
rect 10586 6820 10620 6854
rect 10654 6820 10688 6854
rect 10722 6820 10756 6854
rect 10790 6820 10824 6854
rect 10858 6820 10892 6854
rect 10926 6820 10960 6854
rect 10994 6820 11028 6854
rect 11062 6820 11096 6854
rect 11130 6820 11164 6854
rect 11198 6820 11232 6854
rect 11266 6820 11300 6854
rect 11334 6820 11368 6854
rect 11402 6820 11436 6854
rect 11470 6820 11504 6854
rect 11538 6820 11572 6854
rect 11606 6820 11640 6854
rect 11674 6820 11708 6854
rect 11742 6820 11776 6854
rect 11810 6820 11844 6854
rect 11878 6820 11912 6854
rect 11946 6820 11980 6854
rect 12014 6820 12048 6854
rect 12082 6820 12116 6854
rect 12150 6820 12184 6854
rect 12218 6820 12252 6854
rect 12286 6820 12320 6854
rect 12354 6820 12388 6854
rect 12422 6820 12456 6854
rect 12490 6820 12524 6854
rect 12558 6820 12592 6854
rect 12626 6820 12660 6854
rect 12694 6820 12728 6854
rect 12762 6820 12796 6854
rect 12830 6820 12864 6854
rect 12898 6820 12932 6854
rect 12966 6820 13000 6854
rect 13034 6820 13068 6854
rect 13102 6820 13118 6854
rect 2872 6804 13118 6820
rect 1871 4534 2022 4550
rect 1871 4500 1887 4534
rect 1921 4500 1955 4534
rect 1989 4500 2022 4534
rect 1871 4484 2022 4500
rect 48 3840 114 3856
rect 48 3806 64 3840
rect 98 3806 114 3840
rect 48 3772 114 3806
rect 48 3738 64 3772
rect 98 3738 114 3772
rect 48 3722 114 3738
rect 414 1886 1278 1902
rect 414 1852 430 1886
rect 464 1852 503 1886
rect 537 1852 576 1886
rect 610 1852 649 1886
rect 683 1852 722 1886
rect 756 1852 795 1886
rect 829 1852 868 1886
rect 902 1852 940 1886
rect 974 1852 1012 1886
rect 1046 1852 1084 1886
rect 1118 1852 1156 1886
rect 1190 1852 1228 1886
rect 1262 1852 1278 1886
rect 414 1836 1278 1852
rect 414 356 1278 372
rect 414 322 430 356
rect 464 322 503 356
rect 537 322 576 356
rect 610 322 649 356
rect 683 322 722 356
rect 756 322 795 356
rect 829 322 868 356
rect 902 322 940 356
rect 974 322 1012 356
rect 1046 322 1084 356
rect 1118 322 1156 356
rect 1190 322 1228 356
rect 1262 322 1278 356
rect 414 306 1278 322
rect 13667 1898 14531 1914
rect 13667 1864 13683 1898
rect 13717 1864 13756 1898
rect 13790 1864 13829 1898
rect 13863 1864 13902 1898
rect 13936 1864 13975 1898
rect 14009 1864 14048 1898
rect 14082 1864 14121 1898
rect 14155 1864 14193 1898
rect 14227 1864 14265 1898
rect 14299 1864 14337 1898
rect 14371 1864 14409 1898
rect 14443 1864 14481 1898
rect 14515 1864 14531 1898
rect 13667 1848 14531 1864
rect 13667 368 14531 384
rect 13667 334 13683 368
rect 13717 334 13756 368
rect 13790 334 13829 368
rect 13863 334 13902 368
rect 13936 334 13975 368
rect 14009 334 14048 368
rect 14082 334 14121 368
rect 14155 334 14193 368
rect 14227 334 14265 368
rect 14299 334 14337 368
rect 14371 334 14409 368
rect 14443 334 14481 368
rect 14515 334 14531 368
rect 13667 318 14531 334
<< polycont >>
rect 1684 39238 1718 39272
rect 1684 39170 1718 39204
rect 2888 38820 2922 38854
rect 2957 38820 2991 38854
rect 3026 38820 3060 38854
rect 3095 38820 3129 38854
rect 3164 38820 3198 38854
rect 3233 38820 3267 38854
rect 3302 38820 3336 38854
rect 3371 38820 3405 38854
rect 3440 38820 3474 38854
rect 3509 38820 3543 38854
rect 3578 38820 3612 38854
rect 3647 38820 3681 38854
rect 3716 38820 3750 38854
rect 3785 38820 3819 38854
rect 3854 38820 3888 38854
rect 3923 38820 3957 38854
rect 3992 38820 4026 38854
rect 4061 38820 4095 38854
rect 4130 38820 4164 38854
rect 4199 38820 4233 38854
rect 4268 38820 4302 38854
rect 4337 38820 4371 38854
rect 4406 38820 4440 38854
rect 4475 38820 4509 38854
rect 4544 38820 4578 38854
rect 4613 38820 4647 38854
rect 4682 38820 4716 38854
rect 4751 38820 4785 38854
rect 4820 38820 4854 38854
rect 4889 38820 4923 38854
rect 4958 38820 4992 38854
rect 5027 38820 5061 38854
rect 5096 38820 5130 38854
rect 5165 38820 5199 38854
rect 5234 38820 5268 38854
rect 5303 38820 5337 38854
rect 5372 38820 5406 38854
rect 5441 38820 5475 38854
rect 5510 38820 5544 38854
rect 5579 38820 5613 38854
rect 5648 38820 5682 38854
rect 5717 38820 5751 38854
rect 5786 38820 5820 38854
rect 5855 38820 5889 38854
rect 5924 38820 5958 38854
rect 5993 38820 6027 38854
rect 6062 38820 6096 38854
rect 6131 38820 6165 38854
rect 6200 38820 6234 38854
rect 6268 38820 6302 38854
rect 6336 38820 6370 38854
rect 6404 38820 6438 38854
rect 6472 38820 6506 38854
rect 6540 38820 6574 38854
rect 6608 38820 6642 38854
rect 6676 38820 6710 38854
rect 6744 38820 6778 38854
rect 6812 38820 6846 38854
rect 6880 38820 6914 38854
rect 6948 38820 6982 38854
rect 7016 38820 7050 38854
rect 7084 38820 7118 38854
rect 7152 38820 7186 38854
rect 7220 38820 7254 38854
rect 7288 38820 7322 38854
rect 7356 38820 7390 38854
rect 7424 38820 7458 38854
rect 7492 38820 7526 38854
rect 7560 38820 7594 38854
rect 7628 38820 7662 38854
rect 7696 38820 7730 38854
rect 7764 38820 7798 38854
rect 7832 38820 7866 38854
rect 7900 38820 7934 38854
rect 7968 38820 8002 38854
rect 8036 38820 8070 38854
rect 8104 38820 8138 38854
rect 8172 38820 8206 38854
rect 8240 38820 8274 38854
rect 8308 38820 8342 38854
rect 8376 38820 8410 38854
rect 8444 38820 8478 38854
rect 8512 38820 8546 38854
rect 8580 38820 8614 38854
rect 8648 38820 8682 38854
rect 8716 38820 8750 38854
rect 8784 38820 8818 38854
rect 8852 38820 8886 38854
rect 8920 38820 8954 38854
rect 8988 38820 9022 38854
rect 9056 38820 9090 38854
rect 9124 38820 9158 38854
rect 9192 38820 9226 38854
rect 9260 38820 9294 38854
rect 9328 38820 9362 38854
rect 9396 38820 9430 38854
rect 9464 38820 9498 38854
rect 9532 38820 9566 38854
rect 9600 38820 9634 38854
rect 9668 38820 9702 38854
rect 9736 38820 9770 38854
rect 9804 38820 9838 38854
rect 9872 38820 9906 38854
rect 9940 38820 9974 38854
rect 10008 38820 10042 38854
rect 10076 38820 10110 38854
rect 10144 38820 10178 38854
rect 10212 38820 10246 38854
rect 10280 38820 10314 38854
rect 10348 38820 10382 38854
rect 10416 38820 10450 38854
rect 10484 38820 10518 38854
rect 10552 38820 10586 38854
rect 10620 38820 10654 38854
rect 10688 38820 10722 38854
rect 10756 38820 10790 38854
rect 10824 38820 10858 38854
rect 10892 38820 10926 38854
rect 10960 38820 10994 38854
rect 11028 38820 11062 38854
rect 11096 38820 11130 38854
rect 11164 38820 11198 38854
rect 11232 38820 11266 38854
rect 11300 38820 11334 38854
rect 11368 38820 11402 38854
rect 11436 38820 11470 38854
rect 11504 38820 11538 38854
rect 11572 38820 11606 38854
rect 11640 38820 11674 38854
rect 11708 38820 11742 38854
rect 11776 38820 11810 38854
rect 11844 38820 11878 38854
rect 11912 38820 11946 38854
rect 11980 38820 12014 38854
rect 12048 38820 12082 38854
rect 12116 38820 12150 38854
rect 12184 38820 12218 38854
rect 12252 38820 12286 38854
rect 12320 38820 12354 38854
rect 12388 38820 12422 38854
rect 12456 38820 12490 38854
rect 12524 38820 12558 38854
rect 12592 38820 12626 38854
rect 12660 38820 12694 38854
rect 12728 38820 12762 38854
rect 12796 38820 12830 38854
rect 12864 38820 12898 38854
rect 12932 38820 12966 38854
rect 13000 38820 13034 38854
rect 13068 38820 13102 38854
rect 2888 37290 2922 37324
rect 2957 37290 2991 37324
rect 3026 37290 3060 37324
rect 3095 37290 3129 37324
rect 3164 37290 3198 37324
rect 3233 37290 3267 37324
rect 3302 37290 3336 37324
rect 3371 37290 3405 37324
rect 3440 37290 3474 37324
rect 3509 37290 3543 37324
rect 3578 37290 3612 37324
rect 3647 37290 3681 37324
rect 3716 37290 3750 37324
rect 3785 37290 3819 37324
rect 3854 37290 3888 37324
rect 3923 37290 3957 37324
rect 3992 37290 4026 37324
rect 4061 37290 4095 37324
rect 4130 37290 4164 37324
rect 4199 37290 4233 37324
rect 4268 37290 4302 37324
rect 4337 37290 4371 37324
rect 4406 37290 4440 37324
rect 4475 37290 4509 37324
rect 4544 37290 4578 37324
rect 4613 37290 4647 37324
rect 4682 37290 4716 37324
rect 4751 37290 4785 37324
rect 4820 37290 4854 37324
rect 4889 37290 4923 37324
rect 4958 37290 4992 37324
rect 5027 37290 5061 37324
rect 5096 37290 5130 37324
rect 5165 37290 5199 37324
rect 5234 37290 5268 37324
rect 5303 37290 5337 37324
rect 5372 37290 5406 37324
rect 5441 37290 5475 37324
rect 5510 37290 5544 37324
rect 5579 37290 5613 37324
rect 5648 37290 5682 37324
rect 5717 37290 5751 37324
rect 5786 37290 5820 37324
rect 5855 37290 5889 37324
rect 5924 37290 5958 37324
rect 5993 37290 6027 37324
rect 6062 37290 6096 37324
rect 6131 37290 6165 37324
rect 6200 37290 6234 37324
rect 6268 37290 6302 37324
rect 6336 37290 6370 37324
rect 6404 37290 6438 37324
rect 6472 37290 6506 37324
rect 6540 37290 6574 37324
rect 6608 37290 6642 37324
rect 6676 37290 6710 37324
rect 6744 37290 6778 37324
rect 6812 37290 6846 37324
rect 6880 37290 6914 37324
rect 6948 37290 6982 37324
rect 7016 37290 7050 37324
rect 7084 37290 7118 37324
rect 7152 37290 7186 37324
rect 7220 37290 7254 37324
rect 7288 37290 7322 37324
rect 7356 37290 7390 37324
rect 7424 37290 7458 37324
rect 7492 37290 7526 37324
rect 7560 37290 7594 37324
rect 7628 37290 7662 37324
rect 7696 37290 7730 37324
rect 7764 37290 7798 37324
rect 7832 37290 7866 37324
rect 7900 37290 7934 37324
rect 7968 37290 8002 37324
rect 8036 37290 8070 37324
rect 8104 37290 8138 37324
rect 8172 37290 8206 37324
rect 8240 37290 8274 37324
rect 8308 37290 8342 37324
rect 8376 37290 8410 37324
rect 8444 37290 8478 37324
rect 8512 37290 8546 37324
rect 8580 37290 8614 37324
rect 8648 37290 8682 37324
rect 8716 37290 8750 37324
rect 8784 37290 8818 37324
rect 8852 37290 8886 37324
rect 8920 37290 8954 37324
rect 8988 37290 9022 37324
rect 9056 37290 9090 37324
rect 9124 37290 9158 37324
rect 9192 37290 9226 37324
rect 9260 37290 9294 37324
rect 9328 37290 9362 37324
rect 9396 37290 9430 37324
rect 9464 37290 9498 37324
rect 9532 37290 9566 37324
rect 9600 37290 9634 37324
rect 9668 37290 9702 37324
rect 9736 37290 9770 37324
rect 9804 37290 9838 37324
rect 9872 37290 9906 37324
rect 9940 37290 9974 37324
rect 10008 37290 10042 37324
rect 10076 37290 10110 37324
rect 10144 37290 10178 37324
rect 10212 37290 10246 37324
rect 10280 37290 10314 37324
rect 10348 37290 10382 37324
rect 10416 37290 10450 37324
rect 10484 37290 10518 37324
rect 10552 37290 10586 37324
rect 10620 37290 10654 37324
rect 10688 37290 10722 37324
rect 10756 37290 10790 37324
rect 10824 37290 10858 37324
rect 10892 37290 10926 37324
rect 10960 37290 10994 37324
rect 11028 37290 11062 37324
rect 11096 37290 11130 37324
rect 11164 37290 11198 37324
rect 11232 37290 11266 37324
rect 11300 37290 11334 37324
rect 11368 37290 11402 37324
rect 11436 37290 11470 37324
rect 11504 37290 11538 37324
rect 11572 37290 11606 37324
rect 11640 37290 11674 37324
rect 11708 37290 11742 37324
rect 11776 37290 11810 37324
rect 11844 37290 11878 37324
rect 11912 37290 11946 37324
rect 11980 37290 12014 37324
rect 12048 37290 12082 37324
rect 12116 37290 12150 37324
rect 12184 37290 12218 37324
rect 12252 37290 12286 37324
rect 12320 37290 12354 37324
rect 12388 37290 12422 37324
rect 12456 37290 12490 37324
rect 12524 37290 12558 37324
rect 12592 37290 12626 37324
rect 12660 37290 12694 37324
rect 12728 37290 12762 37324
rect 12796 37290 12830 37324
rect 12864 37290 12898 37324
rect 12932 37290 12966 37324
rect 13000 37290 13034 37324
rect 13068 37290 13102 37324
rect 2888 36820 2922 36854
rect 2957 36820 2991 36854
rect 3026 36820 3060 36854
rect 3095 36820 3129 36854
rect 3164 36820 3198 36854
rect 3233 36820 3267 36854
rect 3302 36820 3336 36854
rect 3371 36820 3405 36854
rect 3440 36820 3474 36854
rect 3509 36820 3543 36854
rect 3578 36820 3612 36854
rect 3647 36820 3681 36854
rect 3716 36820 3750 36854
rect 3785 36820 3819 36854
rect 3854 36820 3888 36854
rect 3923 36820 3957 36854
rect 3992 36820 4026 36854
rect 4061 36820 4095 36854
rect 4130 36820 4164 36854
rect 4199 36820 4233 36854
rect 4268 36820 4302 36854
rect 4337 36820 4371 36854
rect 4406 36820 4440 36854
rect 4475 36820 4509 36854
rect 4544 36820 4578 36854
rect 4613 36820 4647 36854
rect 4682 36820 4716 36854
rect 4751 36820 4785 36854
rect 4820 36820 4854 36854
rect 4889 36820 4923 36854
rect 4958 36820 4992 36854
rect 5027 36820 5061 36854
rect 5096 36820 5130 36854
rect 5165 36820 5199 36854
rect 5234 36820 5268 36854
rect 5303 36820 5337 36854
rect 5372 36820 5406 36854
rect 5441 36820 5475 36854
rect 5510 36820 5544 36854
rect 5579 36820 5613 36854
rect 5648 36820 5682 36854
rect 5717 36820 5751 36854
rect 5786 36820 5820 36854
rect 5855 36820 5889 36854
rect 5924 36820 5958 36854
rect 5993 36820 6027 36854
rect 6062 36820 6096 36854
rect 6131 36820 6165 36854
rect 6200 36820 6234 36854
rect 6268 36820 6302 36854
rect 6336 36820 6370 36854
rect 6404 36820 6438 36854
rect 6472 36820 6506 36854
rect 6540 36820 6574 36854
rect 6608 36820 6642 36854
rect 6676 36820 6710 36854
rect 6744 36820 6778 36854
rect 6812 36820 6846 36854
rect 6880 36820 6914 36854
rect 6948 36820 6982 36854
rect 7016 36820 7050 36854
rect 7084 36820 7118 36854
rect 7152 36820 7186 36854
rect 7220 36820 7254 36854
rect 7288 36820 7322 36854
rect 7356 36820 7390 36854
rect 7424 36820 7458 36854
rect 7492 36820 7526 36854
rect 7560 36820 7594 36854
rect 7628 36820 7662 36854
rect 7696 36820 7730 36854
rect 7764 36820 7798 36854
rect 7832 36820 7866 36854
rect 7900 36820 7934 36854
rect 7968 36820 8002 36854
rect 8036 36820 8070 36854
rect 8104 36820 8138 36854
rect 8172 36820 8206 36854
rect 8240 36820 8274 36854
rect 8308 36820 8342 36854
rect 8376 36820 8410 36854
rect 8444 36820 8478 36854
rect 8512 36820 8546 36854
rect 8580 36820 8614 36854
rect 8648 36820 8682 36854
rect 8716 36820 8750 36854
rect 8784 36820 8818 36854
rect 8852 36820 8886 36854
rect 8920 36820 8954 36854
rect 8988 36820 9022 36854
rect 9056 36820 9090 36854
rect 9124 36820 9158 36854
rect 9192 36820 9226 36854
rect 9260 36820 9294 36854
rect 9328 36820 9362 36854
rect 9396 36820 9430 36854
rect 9464 36820 9498 36854
rect 9532 36820 9566 36854
rect 9600 36820 9634 36854
rect 9668 36820 9702 36854
rect 9736 36820 9770 36854
rect 9804 36820 9838 36854
rect 9872 36820 9906 36854
rect 9940 36820 9974 36854
rect 10008 36820 10042 36854
rect 10076 36820 10110 36854
rect 10144 36820 10178 36854
rect 10212 36820 10246 36854
rect 10280 36820 10314 36854
rect 10348 36820 10382 36854
rect 10416 36820 10450 36854
rect 10484 36820 10518 36854
rect 10552 36820 10586 36854
rect 10620 36820 10654 36854
rect 10688 36820 10722 36854
rect 10756 36820 10790 36854
rect 10824 36820 10858 36854
rect 10892 36820 10926 36854
rect 10960 36820 10994 36854
rect 11028 36820 11062 36854
rect 11096 36820 11130 36854
rect 11164 36820 11198 36854
rect 11232 36820 11266 36854
rect 11300 36820 11334 36854
rect 11368 36820 11402 36854
rect 11436 36820 11470 36854
rect 11504 36820 11538 36854
rect 11572 36820 11606 36854
rect 11640 36820 11674 36854
rect 11708 36820 11742 36854
rect 11776 36820 11810 36854
rect 11844 36820 11878 36854
rect 11912 36820 11946 36854
rect 11980 36820 12014 36854
rect 12048 36820 12082 36854
rect 12116 36820 12150 36854
rect 12184 36820 12218 36854
rect 12252 36820 12286 36854
rect 12320 36820 12354 36854
rect 12388 36820 12422 36854
rect 12456 36820 12490 36854
rect 12524 36820 12558 36854
rect 12592 36820 12626 36854
rect 12660 36820 12694 36854
rect 12728 36820 12762 36854
rect 12796 36820 12830 36854
rect 12864 36820 12898 36854
rect 12932 36820 12966 36854
rect 13000 36820 13034 36854
rect 13068 36820 13102 36854
rect 2888 35290 2922 35324
rect 2957 35290 2991 35324
rect 3026 35290 3060 35324
rect 3095 35290 3129 35324
rect 3164 35290 3198 35324
rect 3233 35290 3267 35324
rect 3302 35290 3336 35324
rect 3371 35290 3405 35324
rect 3440 35290 3474 35324
rect 3509 35290 3543 35324
rect 3578 35290 3612 35324
rect 3647 35290 3681 35324
rect 3716 35290 3750 35324
rect 3785 35290 3819 35324
rect 3854 35290 3888 35324
rect 3923 35290 3957 35324
rect 3992 35290 4026 35324
rect 4061 35290 4095 35324
rect 4130 35290 4164 35324
rect 4199 35290 4233 35324
rect 4268 35290 4302 35324
rect 4337 35290 4371 35324
rect 4406 35290 4440 35324
rect 4475 35290 4509 35324
rect 4544 35290 4578 35324
rect 4613 35290 4647 35324
rect 4682 35290 4716 35324
rect 4751 35290 4785 35324
rect 4820 35290 4854 35324
rect 4889 35290 4923 35324
rect 4958 35290 4992 35324
rect 5027 35290 5061 35324
rect 5096 35290 5130 35324
rect 5165 35290 5199 35324
rect 5234 35290 5268 35324
rect 5303 35290 5337 35324
rect 5372 35290 5406 35324
rect 5441 35290 5475 35324
rect 5510 35290 5544 35324
rect 5579 35290 5613 35324
rect 5648 35290 5682 35324
rect 5717 35290 5751 35324
rect 5786 35290 5820 35324
rect 5855 35290 5889 35324
rect 5924 35290 5958 35324
rect 5993 35290 6027 35324
rect 6062 35290 6096 35324
rect 6131 35290 6165 35324
rect 6200 35290 6234 35324
rect 6268 35290 6302 35324
rect 6336 35290 6370 35324
rect 6404 35290 6438 35324
rect 6472 35290 6506 35324
rect 6540 35290 6574 35324
rect 6608 35290 6642 35324
rect 6676 35290 6710 35324
rect 6744 35290 6778 35324
rect 6812 35290 6846 35324
rect 6880 35290 6914 35324
rect 6948 35290 6982 35324
rect 7016 35290 7050 35324
rect 7084 35290 7118 35324
rect 7152 35290 7186 35324
rect 7220 35290 7254 35324
rect 7288 35290 7322 35324
rect 7356 35290 7390 35324
rect 7424 35290 7458 35324
rect 7492 35290 7526 35324
rect 7560 35290 7594 35324
rect 7628 35290 7662 35324
rect 7696 35290 7730 35324
rect 7764 35290 7798 35324
rect 7832 35290 7866 35324
rect 7900 35290 7934 35324
rect 7968 35290 8002 35324
rect 8036 35290 8070 35324
rect 8104 35290 8138 35324
rect 8172 35290 8206 35324
rect 8240 35290 8274 35324
rect 8308 35290 8342 35324
rect 8376 35290 8410 35324
rect 8444 35290 8478 35324
rect 8512 35290 8546 35324
rect 8580 35290 8614 35324
rect 8648 35290 8682 35324
rect 8716 35290 8750 35324
rect 8784 35290 8818 35324
rect 8852 35290 8886 35324
rect 8920 35290 8954 35324
rect 8988 35290 9022 35324
rect 9056 35290 9090 35324
rect 9124 35290 9158 35324
rect 9192 35290 9226 35324
rect 9260 35290 9294 35324
rect 9328 35290 9362 35324
rect 9396 35290 9430 35324
rect 9464 35290 9498 35324
rect 9532 35290 9566 35324
rect 9600 35290 9634 35324
rect 9668 35290 9702 35324
rect 9736 35290 9770 35324
rect 9804 35290 9838 35324
rect 9872 35290 9906 35324
rect 9940 35290 9974 35324
rect 10008 35290 10042 35324
rect 10076 35290 10110 35324
rect 10144 35290 10178 35324
rect 10212 35290 10246 35324
rect 10280 35290 10314 35324
rect 10348 35290 10382 35324
rect 10416 35290 10450 35324
rect 10484 35290 10518 35324
rect 10552 35290 10586 35324
rect 10620 35290 10654 35324
rect 10688 35290 10722 35324
rect 10756 35290 10790 35324
rect 10824 35290 10858 35324
rect 10892 35290 10926 35324
rect 10960 35290 10994 35324
rect 11028 35290 11062 35324
rect 11096 35290 11130 35324
rect 11164 35290 11198 35324
rect 11232 35290 11266 35324
rect 11300 35290 11334 35324
rect 11368 35290 11402 35324
rect 11436 35290 11470 35324
rect 11504 35290 11538 35324
rect 11572 35290 11606 35324
rect 11640 35290 11674 35324
rect 11708 35290 11742 35324
rect 11776 35290 11810 35324
rect 11844 35290 11878 35324
rect 11912 35290 11946 35324
rect 11980 35290 12014 35324
rect 12048 35290 12082 35324
rect 12116 35290 12150 35324
rect 12184 35290 12218 35324
rect 12252 35290 12286 35324
rect 12320 35290 12354 35324
rect 12388 35290 12422 35324
rect 12456 35290 12490 35324
rect 12524 35290 12558 35324
rect 12592 35290 12626 35324
rect 12660 35290 12694 35324
rect 12728 35290 12762 35324
rect 12796 35290 12830 35324
rect 12864 35290 12898 35324
rect 12932 35290 12966 35324
rect 13000 35290 13034 35324
rect 13068 35290 13102 35324
rect 3507 34820 3541 34854
rect 3576 34820 3610 34854
rect 3645 34820 3679 34854
rect 3714 34820 3748 34854
rect 3783 34820 3817 34854
rect 3852 34820 3886 34854
rect 3921 34820 3955 34854
rect 3990 34820 4024 34854
rect 4059 34820 4093 34854
rect 4128 34820 4162 34854
rect 4197 34820 4231 34854
rect 4266 34820 4300 34854
rect 4335 34820 4369 34854
rect 4404 34820 4438 34854
rect 4473 34820 4507 34854
rect 4542 34820 4576 34854
rect 4611 34820 4645 34854
rect 4680 34820 4714 34854
rect 4749 34820 4783 34854
rect 4818 34820 4852 34854
rect 4887 34820 4921 34854
rect 4956 34820 4990 34854
rect 5025 34820 5059 34854
rect 5094 34820 5128 34854
rect 5163 34820 5197 34854
rect 5232 34820 5266 34854
rect 5301 34820 5335 34854
rect 5370 34820 5404 34854
rect 5439 34820 5473 34854
rect 5508 34820 5542 34854
rect 5577 34820 5611 34854
rect 5646 34820 5680 34854
rect 5715 34820 5749 34854
rect 5784 34820 5818 34854
rect 5853 34820 5887 34854
rect 5922 34820 5956 34854
rect 5991 34820 6025 34854
rect 6060 34820 6094 34854
rect 6129 34820 6163 34854
rect 6198 34820 6232 34854
rect 6267 34820 6301 34854
rect 6336 34820 6370 34854
rect 6405 34820 6439 34854
rect 6474 34820 6508 34854
rect 6543 34820 6577 34854
rect 6612 34820 6646 34854
rect 6681 34820 6715 34854
rect 6750 34820 6784 34854
rect 6819 34820 6853 34854
rect 6888 34820 6922 34854
rect 6957 34820 6991 34854
rect 7026 34820 7060 34854
rect 7095 34820 7129 34854
rect 7163 34820 7197 34854
rect 7231 34820 7265 34854
rect 7299 34820 7333 34854
rect 7367 34820 7401 34854
rect 7435 34820 7469 34854
rect 7503 34820 7537 34854
rect 7571 34820 7605 34854
rect 7639 34820 7673 34854
rect 7707 34820 7741 34854
rect 7775 34820 7809 34854
rect 7843 34820 7877 34854
rect 7911 34820 7945 34854
rect 7979 34820 8013 34854
rect 8047 34820 8081 34854
rect 8115 34820 8149 34854
rect 8183 34820 8217 34854
rect 8251 34820 8285 34854
rect 8319 34820 8353 34854
rect 8387 34820 8421 34854
rect 8455 34820 8489 34854
rect 8523 34820 8557 34854
rect 8591 34820 8625 34854
rect 8659 34820 8693 34854
rect 8727 34820 8761 34854
rect 8795 34820 8829 34854
rect 8863 34820 8897 34854
rect 8931 34820 8965 34854
rect 8999 34820 9033 34854
rect 9067 34820 9101 34854
rect 9135 34820 9169 34854
rect 9203 34820 9237 34854
rect 9271 34820 9305 34854
rect 9339 34820 9373 34854
rect 9407 34820 9441 34854
rect 9475 34820 9509 34854
rect 9543 34820 9577 34854
rect 9611 34820 9645 34854
rect 9679 34820 9713 34854
rect 9747 34820 9781 34854
rect 9815 34820 9849 34854
rect 9883 34820 9917 34854
rect 9951 34820 9985 34854
rect 10019 34820 10053 34854
rect 10087 34820 10121 34854
rect 10155 34820 10189 34854
rect 10223 34820 10257 34854
rect 10291 34820 10325 34854
rect 10359 34820 10393 34854
rect 10427 34820 10461 34854
rect 10495 34820 10529 34854
rect 10563 34820 10597 34854
rect 10631 34820 10665 34854
rect 10699 34820 10733 34854
rect 10767 34820 10801 34854
rect 10835 34820 10869 34854
rect 10903 34820 10937 34854
rect 10971 34820 11005 34854
rect 11039 34820 11073 34854
rect 11107 34820 11141 34854
rect 11175 34820 11209 34854
rect 11243 34820 11277 34854
rect 11311 34820 11345 34854
rect 11379 34820 11413 34854
rect 11447 34820 11481 34854
rect 11515 34820 11549 34854
rect 11583 34820 11617 34854
rect 11651 34820 11685 34854
rect 11719 34820 11753 34854
rect 11787 34820 11821 34854
rect 11855 34820 11889 34854
rect 11923 34820 11957 34854
rect 11991 34820 12025 34854
rect 12059 34820 12093 34854
rect 12127 34820 12161 34854
rect 12195 34820 12229 34854
rect 12263 34820 12297 34854
rect 12331 34820 12365 34854
rect 12399 34820 12433 34854
rect 12467 34820 12501 34854
rect 12535 34820 12569 34854
rect 12603 34820 12637 34854
rect 12671 34820 12705 34854
rect 12739 34820 12773 34854
rect 12807 34820 12841 34854
rect 12875 34820 12909 34854
rect 12943 34820 12977 34854
rect 3507 33290 3541 33324
rect 3576 33290 3610 33324
rect 3645 33290 3679 33324
rect 3714 33290 3748 33324
rect 3783 33290 3817 33324
rect 3852 33290 3886 33324
rect 3921 33290 3955 33324
rect 3990 33290 4024 33324
rect 4059 33290 4093 33324
rect 4128 33290 4162 33324
rect 4197 33290 4231 33324
rect 4266 33290 4300 33324
rect 4335 33290 4369 33324
rect 4404 33290 4438 33324
rect 4473 33290 4507 33324
rect 4542 33290 4576 33324
rect 4611 33290 4645 33324
rect 4680 33290 4714 33324
rect 4749 33290 4783 33324
rect 4818 33290 4852 33324
rect 4887 33290 4921 33324
rect 4956 33290 4990 33324
rect 5025 33290 5059 33324
rect 5094 33290 5128 33324
rect 5163 33290 5197 33324
rect 5232 33290 5266 33324
rect 5301 33290 5335 33324
rect 5370 33290 5404 33324
rect 5439 33290 5473 33324
rect 5508 33290 5542 33324
rect 5577 33290 5611 33324
rect 5646 33290 5680 33324
rect 5715 33290 5749 33324
rect 5784 33290 5818 33324
rect 5853 33290 5887 33324
rect 5922 33290 5956 33324
rect 5991 33290 6025 33324
rect 6060 33290 6094 33324
rect 6129 33290 6163 33324
rect 6198 33290 6232 33324
rect 6267 33290 6301 33324
rect 6336 33290 6370 33324
rect 6405 33290 6439 33324
rect 6474 33290 6508 33324
rect 6543 33290 6577 33324
rect 6612 33290 6646 33324
rect 6681 33290 6715 33324
rect 6750 33290 6784 33324
rect 6819 33290 6853 33324
rect 6888 33290 6922 33324
rect 6957 33290 6991 33324
rect 7026 33290 7060 33324
rect 7095 33290 7129 33324
rect 7163 33290 7197 33324
rect 7231 33290 7265 33324
rect 7299 33290 7333 33324
rect 7367 33290 7401 33324
rect 7435 33290 7469 33324
rect 7503 33290 7537 33324
rect 7571 33290 7605 33324
rect 7639 33290 7673 33324
rect 7707 33290 7741 33324
rect 7775 33290 7809 33324
rect 7843 33290 7877 33324
rect 7911 33290 7945 33324
rect 7979 33290 8013 33324
rect 8047 33290 8081 33324
rect 8115 33290 8149 33324
rect 8183 33290 8217 33324
rect 8251 33290 8285 33324
rect 8319 33290 8353 33324
rect 8387 33290 8421 33324
rect 8455 33290 8489 33324
rect 8523 33290 8557 33324
rect 8591 33290 8625 33324
rect 8659 33290 8693 33324
rect 8727 33290 8761 33324
rect 8795 33290 8829 33324
rect 8863 33290 8897 33324
rect 8931 33290 8965 33324
rect 8999 33290 9033 33324
rect 9067 33290 9101 33324
rect 9135 33290 9169 33324
rect 9203 33290 9237 33324
rect 9271 33290 9305 33324
rect 9339 33290 9373 33324
rect 9407 33290 9441 33324
rect 9475 33290 9509 33324
rect 9543 33290 9577 33324
rect 9611 33290 9645 33324
rect 9679 33290 9713 33324
rect 9747 33290 9781 33324
rect 9815 33290 9849 33324
rect 9883 33290 9917 33324
rect 9951 33290 9985 33324
rect 10019 33290 10053 33324
rect 10087 33290 10121 33324
rect 10155 33290 10189 33324
rect 10223 33290 10257 33324
rect 10291 33290 10325 33324
rect 10359 33290 10393 33324
rect 10427 33290 10461 33324
rect 10495 33290 10529 33324
rect 10563 33290 10597 33324
rect 10631 33290 10665 33324
rect 10699 33290 10733 33324
rect 10767 33290 10801 33324
rect 10835 33290 10869 33324
rect 10903 33290 10937 33324
rect 10971 33290 11005 33324
rect 11039 33290 11073 33324
rect 11107 33290 11141 33324
rect 11175 33290 11209 33324
rect 11243 33290 11277 33324
rect 11311 33290 11345 33324
rect 11379 33290 11413 33324
rect 11447 33290 11481 33324
rect 11515 33290 11549 33324
rect 11583 33290 11617 33324
rect 11651 33290 11685 33324
rect 11719 33290 11753 33324
rect 11787 33290 11821 33324
rect 11855 33290 11889 33324
rect 11923 33290 11957 33324
rect 11991 33290 12025 33324
rect 12059 33290 12093 33324
rect 12127 33290 12161 33324
rect 12195 33290 12229 33324
rect 12263 33290 12297 33324
rect 12331 33290 12365 33324
rect 12399 33290 12433 33324
rect 12467 33290 12501 33324
rect 12535 33290 12569 33324
rect 12603 33290 12637 33324
rect 12671 33290 12705 33324
rect 12739 33290 12773 33324
rect 12807 33290 12841 33324
rect 12875 33290 12909 33324
rect 12943 33290 12977 33324
rect 3507 32820 3541 32854
rect 3576 32820 3610 32854
rect 3645 32820 3679 32854
rect 3714 32820 3748 32854
rect 3783 32820 3817 32854
rect 3852 32820 3886 32854
rect 3921 32820 3955 32854
rect 3990 32820 4024 32854
rect 4059 32820 4093 32854
rect 4128 32820 4162 32854
rect 4197 32820 4231 32854
rect 4266 32820 4300 32854
rect 4335 32820 4369 32854
rect 4404 32820 4438 32854
rect 4473 32820 4507 32854
rect 4542 32820 4576 32854
rect 4611 32820 4645 32854
rect 4680 32820 4714 32854
rect 4749 32820 4783 32854
rect 4818 32820 4852 32854
rect 4887 32820 4921 32854
rect 4956 32820 4990 32854
rect 5025 32820 5059 32854
rect 5094 32820 5128 32854
rect 5163 32820 5197 32854
rect 5232 32820 5266 32854
rect 5301 32820 5335 32854
rect 5370 32820 5404 32854
rect 5439 32820 5473 32854
rect 5508 32820 5542 32854
rect 5577 32820 5611 32854
rect 5646 32820 5680 32854
rect 5715 32820 5749 32854
rect 5784 32820 5818 32854
rect 5853 32820 5887 32854
rect 5922 32820 5956 32854
rect 5991 32820 6025 32854
rect 6060 32820 6094 32854
rect 6129 32820 6163 32854
rect 6198 32820 6232 32854
rect 6267 32820 6301 32854
rect 6336 32820 6370 32854
rect 6405 32820 6439 32854
rect 6474 32820 6508 32854
rect 6543 32820 6577 32854
rect 6612 32820 6646 32854
rect 6681 32820 6715 32854
rect 6750 32820 6784 32854
rect 6819 32820 6853 32854
rect 6888 32820 6922 32854
rect 6957 32820 6991 32854
rect 7026 32820 7060 32854
rect 7095 32820 7129 32854
rect 7163 32820 7197 32854
rect 7231 32820 7265 32854
rect 7299 32820 7333 32854
rect 7367 32820 7401 32854
rect 7435 32820 7469 32854
rect 7503 32820 7537 32854
rect 7571 32820 7605 32854
rect 7639 32820 7673 32854
rect 7707 32820 7741 32854
rect 7775 32820 7809 32854
rect 7843 32820 7877 32854
rect 7911 32820 7945 32854
rect 7979 32820 8013 32854
rect 8047 32820 8081 32854
rect 8115 32820 8149 32854
rect 8183 32820 8217 32854
rect 8251 32820 8285 32854
rect 8319 32820 8353 32854
rect 8387 32820 8421 32854
rect 8455 32820 8489 32854
rect 8523 32820 8557 32854
rect 8591 32820 8625 32854
rect 8659 32820 8693 32854
rect 8727 32820 8761 32854
rect 8795 32820 8829 32854
rect 8863 32820 8897 32854
rect 8931 32820 8965 32854
rect 8999 32820 9033 32854
rect 9067 32820 9101 32854
rect 9135 32820 9169 32854
rect 9203 32820 9237 32854
rect 9271 32820 9305 32854
rect 9339 32820 9373 32854
rect 9407 32820 9441 32854
rect 9475 32820 9509 32854
rect 9543 32820 9577 32854
rect 9611 32820 9645 32854
rect 9679 32820 9713 32854
rect 9747 32820 9781 32854
rect 9815 32820 9849 32854
rect 9883 32820 9917 32854
rect 9951 32820 9985 32854
rect 10019 32820 10053 32854
rect 10087 32820 10121 32854
rect 10155 32820 10189 32854
rect 10223 32820 10257 32854
rect 10291 32820 10325 32854
rect 10359 32820 10393 32854
rect 10427 32820 10461 32854
rect 10495 32820 10529 32854
rect 10563 32820 10597 32854
rect 10631 32820 10665 32854
rect 10699 32820 10733 32854
rect 10767 32820 10801 32854
rect 10835 32820 10869 32854
rect 10903 32820 10937 32854
rect 10971 32820 11005 32854
rect 11039 32820 11073 32854
rect 11107 32820 11141 32854
rect 11175 32820 11209 32854
rect 11243 32820 11277 32854
rect 11311 32820 11345 32854
rect 11379 32820 11413 32854
rect 11447 32820 11481 32854
rect 11515 32820 11549 32854
rect 11583 32820 11617 32854
rect 11651 32820 11685 32854
rect 11719 32820 11753 32854
rect 11787 32820 11821 32854
rect 11855 32820 11889 32854
rect 11923 32820 11957 32854
rect 11991 32820 12025 32854
rect 12059 32820 12093 32854
rect 12127 32820 12161 32854
rect 12195 32820 12229 32854
rect 12263 32820 12297 32854
rect 12331 32820 12365 32854
rect 12399 32820 12433 32854
rect 12467 32820 12501 32854
rect 12535 32820 12569 32854
rect 12603 32820 12637 32854
rect 12671 32820 12705 32854
rect 12739 32820 12773 32854
rect 12807 32820 12841 32854
rect 12875 32820 12909 32854
rect 12943 32820 12977 32854
rect 3507 31290 3541 31324
rect 3576 31290 3610 31324
rect 3645 31290 3679 31324
rect 3714 31290 3748 31324
rect 3783 31290 3817 31324
rect 3852 31290 3886 31324
rect 3921 31290 3955 31324
rect 3990 31290 4024 31324
rect 4059 31290 4093 31324
rect 4128 31290 4162 31324
rect 4197 31290 4231 31324
rect 4266 31290 4300 31324
rect 4335 31290 4369 31324
rect 4404 31290 4438 31324
rect 4473 31290 4507 31324
rect 4542 31290 4576 31324
rect 4611 31290 4645 31324
rect 4680 31290 4714 31324
rect 4749 31290 4783 31324
rect 4818 31290 4852 31324
rect 4887 31290 4921 31324
rect 4956 31290 4990 31324
rect 5025 31290 5059 31324
rect 5094 31290 5128 31324
rect 5163 31290 5197 31324
rect 5232 31290 5266 31324
rect 5301 31290 5335 31324
rect 5370 31290 5404 31324
rect 5439 31290 5473 31324
rect 5508 31290 5542 31324
rect 5577 31290 5611 31324
rect 5646 31290 5680 31324
rect 5715 31290 5749 31324
rect 5784 31290 5818 31324
rect 5853 31290 5887 31324
rect 5922 31290 5956 31324
rect 5991 31290 6025 31324
rect 6060 31290 6094 31324
rect 6129 31290 6163 31324
rect 6198 31290 6232 31324
rect 6267 31290 6301 31324
rect 6336 31290 6370 31324
rect 6405 31290 6439 31324
rect 6474 31290 6508 31324
rect 6543 31290 6577 31324
rect 6612 31290 6646 31324
rect 6681 31290 6715 31324
rect 6750 31290 6784 31324
rect 6819 31290 6853 31324
rect 6888 31290 6922 31324
rect 6957 31290 6991 31324
rect 7026 31290 7060 31324
rect 7095 31290 7129 31324
rect 7163 31290 7197 31324
rect 7231 31290 7265 31324
rect 7299 31290 7333 31324
rect 7367 31290 7401 31324
rect 7435 31290 7469 31324
rect 7503 31290 7537 31324
rect 7571 31290 7605 31324
rect 7639 31290 7673 31324
rect 7707 31290 7741 31324
rect 7775 31290 7809 31324
rect 7843 31290 7877 31324
rect 7911 31290 7945 31324
rect 7979 31290 8013 31324
rect 8047 31290 8081 31324
rect 8115 31290 8149 31324
rect 8183 31290 8217 31324
rect 8251 31290 8285 31324
rect 8319 31290 8353 31324
rect 8387 31290 8421 31324
rect 8455 31290 8489 31324
rect 8523 31290 8557 31324
rect 8591 31290 8625 31324
rect 8659 31290 8693 31324
rect 8727 31290 8761 31324
rect 8795 31290 8829 31324
rect 8863 31290 8897 31324
rect 8931 31290 8965 31324
rect 8999 31290 9033 31324
rect 9067 31290 9101 31324
rect 9135 31290 9169 31324
rect 9203 31290 9237 31324
rect 9271 31290 9305 31324
rect 9339 31290 9373 31324
rect 9407 31290 9441 31324
rect 9475 31290 9509 31324
rect 9543 31290 9577 31324
rect 9611 31290 9645 31324
rect 9679 31290 9713 31324
rect 9747 31290 9781 31324
rect 9815 31290 9849 31324
rect 9883 31290 9917 31324
rect 9951 31290 9985 31324
rect 10019 31290 10053 31324
rect 10087 31290 10121 31324
rect 10155 31290 10189 31324
rect 10223 31290 10257 31324
rect 10291 31290 10325 31324
rect 10359 31290 10393 31324
rect 10427 31290 10461 31324
rect 10495 31290 10529 31324
rect 10563 31290 10597 31324
rect 10631 31290 10665 31324
rect 10699 31290 10733 31324
rect 10767 31290 10801 31324
rect 10835 31290 10869 31324
rect 10903 31290 10937 31324
rect 10971 31290 11005 31324
rect 11039 31290 11073 31324
rect 11107 31290 11141 31324
rect 11175 31290 11209 31324
rect 11243 31290 11277 31324
rect 11311 31290 11345 31324
rect 11379 31290 11413 31324
rect 11447 31290 11481 31324
rect 11515 31290 11549 31324
rect 11583 31290 11617 31324
rect 11651 31290 11685 31324
rect 11719 31290 11753 31324
rect 11787 31290 11821 31324
rect 11855 31290 11889 31324
rect 11923 31290 11957 31324
rect 11991 31290 12025 31324
rect 12059 31290 12093 31324
rect 12127 31290 12161 31324
rect 12195 31290 12229 31324
rect 12263 31290 12297 31324
rect 12331 31290 12365 31324
rect 12399 31290 12433 31324
rect 12467 31290 12501 31324
rect 12535 31290 12569 31324
rect 12603 31290 12637 31324
rect 12671 31290 12705 31324
rect 12739 31290 12773 31324
rect 12807 31290 12841 31324
rect 12875 31290 12909 31324
rect 12943 31290 12977 31324
rect 3507 30820 3541 30854
rect 3576 30820 3610 30854
rect 3645 30820 3679 30854
rect 3714 30820 3748 30854
rect 3783 30820 3817 30854
rect 3852 30820 3886 30854
rect 3921 30820 3955 30854
rect 3990 30820 4024 30854
rect 4059 30820 4093 30854
rect 4128 30820 4162 30854
rect 4197 30820 4231 30854
rect 4266 30820 4300 30854
rect 4335 30820 4369 30854
rect 4404 30820 4438 30854
rect 4473 30820 4507 30854
rect 4542 30820 4576 30854
rect 4611 30820 4645 30854
rect 4680 30820 4714 30854
rect 4749 30820 4783 30854
rect 4818 30820 4852 30854
rect 4887 30820 4921 30854
rect 4956 30820 4990 30854
rect 5025 30820 5059 30854
rect 5094 30820 5128 30854
rect 5163 30820 5197 30854
rect 5232 30820 5266 30854
rect 5301 30820 5335 30854
rect 5370 30820 5404 30854
rect 5439 30820 5473 30854
rect 5508 30820 5542 30854
rect 5577 30820 5611 30854
rect 5646 30820 5680 30854
rect 5715 30820 5749 30854
rect 5784 30820 5818 30854
rect 5853 30820 5887 30854
rect 5922 30820 5956 30854
rect 5991 30820 6025 30854
rect 6060 30820 6094 30854
rect 6129 30820 6163 30854
rect 6198 30820 6232 30854
rect 6267 30820 6301 30854
rect 6336 30820 6370 30854
rect 6405 30820 6439 30854
rect 6474 30820 6508 30854
rect 6543 30820 6577 30854
rect 6612 30820 6646 30854
rect 6681 30820 6715 30854
rect 6750 30820 6784 30854
rect 6819 30820 6853 30854
rect 6888 30820 6922 30854
rect 6957 30820 6991 30854
rect 7026 30820 7060 30854
rect 7095 30820 7129 30854
rect 7163 30820 7197 30854
rect 7231 30820 7265 30854
rect 7299 30820 7333 30854
rect 7367 30820 7401 30854
rect 7435 30820 7469 30854
rect 7503 30820 7537 30854
rect 7571 30820 7605 30854
rect 7639 30820 7673 30854
rect 7707 30820 7741 30854
rect 7775 30820 7809 30854
rect 7843 30820 7877 30854
rect 7911 30820 7945 30854
rect 7979 30820 8013 30854
rect 8047 30820 8081 30854
rect 8115 30820 8149 30854
rect 8183 30820 8217 30854
rect 8251 30820 8285 30854
rect 8319 30820 8353 30854
rect 8387 30820 8421 30854
rect 8455 30820 8489 30854
rect 8523 30820 8557 30854
rect 8591 30820 8625 30854
rect 8659 30820 8693 30854
rect 8727 30820 8761 30854
rect 8795 30820 8829 30854
rect 8863 30820 8897 30854
rect 8931 30820 8965 30854
rect 8999 30820 9033 30854
rect 9067 30820 9101 30854
rect 9135 30820 9169 30854
rect 9203 30820 9237 30854
rect 9271 30820 9305 30854
rect 9339 30820 9373 30854
rect 9407 30820 9441 30854
rect 9475 30820 9509 30854
rect 9543 30820 9577 30854
rect 9611 30820 9645 30854
rect 9679 30820 9713 30854
rect 9747 30820 9781 30854
rect 9815 30820 9849 30854
rect 9883 30820 9917 30854
rect 9951 30820 9985 30854
rect 10019 30820 10053 30854
rect 10087 30820 10121 30854
rect 10155 30820 10189 30854
rect 10223 30820 10257 30854
rect 10291 30820 10325 30854
rect 10359 30820 10393 30854
rect 10427 30820 10461 30854
rect 10495 30820 10529 30854
rect 10563 30820 10597 30854
rect 10631 30820 10665 30854
rect 10699 30820 10733 30854
rect 10767 30820 10801 30854
rect 10835 30820 10869 30854
rect 10903 30820 10937 30854
rect 10971 30820 11005 30854
rect 11039 30820 11073 30854
rect 11107 30820 11141 30854
rect 11175 30820 11209 30854
rect 11243 30820 11277 30854
rect 11311 30820 11345 30854
rect 11379 30820 11413 30854
rect 11447 30820 11481 30854
rect 11515 30820 11549 30854
rect 11583 30820 11617 30854
rect 11651 30820 11685 30854
rect 11719 30820 11753 30854
rect 11787 30820 11821 30854
rect 11855 30820 11889 30854
rect 11923 30820 11957 30854
rect 11991 30820 12025 30854
rect 12059 30820 12093 30854
rect 12127 30820 12161 30854
rect 12195 30820 12229 30854
rect 12263 30820 12297 30854
rect 12331 30820 12365 30854
rect 12399 30820 12433 30854
rect 12467 30820 12501 30854
rect 12535 30820 12569 30854
rect 12603 30820 12637 30854
rect 12671 30820 12705 30854
rect 12739 30820 12773 30854
rect 12807 30820 12841 30854
rect 12875 30820 12909 30854
rect 12943 30820 12977 30854
rect 3507 29290 3541 29324
rect 3576 29290 3610 29324
rect 3645 29290 3679 29324
rect 3714 29290 3748 29324
rect 3783 29290 3817 29324
rect 3852 29290 3886 29324
rect 3921 29290 3955 29324
rect 3990 29290 4024 29324
rect 4059 29290 4093 29324
rect 4128 29290 4162 29324
rect 4197 29290 4231 29324
rect 4266 29290 4300 29324
rect 4335 29290 4369 29324
rect 4404 29290 4438 29324
rect 4473 29290 4507 29324
rect 4542 29290 4576 29324
rect 4611 29290 4645 29324
rect 4680 29290 4714 29324
rect 4749 29290 4783 29324
rect 4818 29290 4852 29324
rect 4887 29290 4921 29324
rect 4956 29290 4990 29324
rect 5025 29290 5059 29324
rect 5094 29290 5128 29324
rect 5163 29290 5197 29324
rect 5232 29290 5266 29324
rect 5301 29290 5335 29324
rect 5370 29290 5404 29324
rect 5439 29290 5473 29324
rect 5508 29290 5542 29324
rect 5577 29290 5611 29324
rect 5646 29290 5680 29324
rect 5715 29290 5749 29324
rect 5784 29290 5818 29324
rect 5853 29290 5887 29324
rect 5922 29290 5956 29324
rect 5991 29290 6025 29324
rect 6060 29290 6094 29324
rect 6129 29290 6163 29324
rect 6198 29290 6232 29324
rect 6267 29290 6301 29324
rect 6336 29290 6370 29324
rect 6405 29290 6439 29324
rect 6474 29290 6508 29324
rect 6543 29290 6577 29324
rect 6612 29290 6646 29324
rect 6681 29290 6715 29324
rect 6750 29290 6784 29324
rect 6819 29290 6853 29324
rect 6888 29290 6922 29324
rect 6957 29290 6991 29324
rect 7026 29290 7060 29324
rect 7095 29290 7129 29324
rect 7163 29290 7197 29324
rect 7231 29290 7265 29324
rect 7299 29290 7333 29324
rect 7367 29290 7401 29324
rect 7435 29290 7469 29324
rect 7503 29290 7537 29324
rect 7571 29290 7605 29324
rect 7639 29290 7673 29324
rect 7707 29290 7741 29324
rect 7775 29290 7809 29324
rect 7843 29290 7877 29324
rect 7911 29290 7945 29324
rect 7979 29290 8013 29324
rect 8047 29290 8081 29324
rect 8115 29290 8149 29324
rect 8183 29290 8217 29324
rect 8251 29290 8285 29324
rect 8319 29290 8353 29324
rect 8387 29290 8421 29324
rect 8455 29290 8489 29324
rect 8523 29290 8557 29324
rect 8591 29290 8625 29324
rect 8659 29290 8693 29324
rect 8727 29290 8761 29324
rect 8795 29290 8829 29324
rect 8863 29290 8897 29324
rect 8931 29290 8965 29324
rect 8999 29290 9033 29324
rect 9067 29290 9101 29324
rect 9135 29290 9169 29324
rect 9203 29290 9237 29324
rect 9271 29290 9305 29324
rect 9339 29290 9373 29324
rect 9407 29290 9441 29324
rect 9475 29290 9509 29324
rect 9543 29290 9577 29324
rect 9611 29290 9645 29324
rect 9679 29290 9713 29324
rect 9747 29290 9781 29324
rect 9815 29290 9849 29324
rect 9883 29290 9917 29324
rect 9951 29290 9985 29324
rect 10019 29290 10053 29324
rect 10087 29290 10121 29324
rect 10155 29290 10189 29324
rect 10223 29290 10257 29324
rect 10291 29290 10325 29324
rect 10359 29290 10393 29324
rect 10427 29290 10461 29324
rect 10495 29290 10529 29324
rect 10563 29290 10597 29324
rect 10631 29290 10665 29324
rect 10699 29290 10733 29324
rect 10767 29290 10801 29324
rect 10835 29290 10869 29324
rect 10903 29290 10937 29324
rect 10971 29290 11005 29324
rect 11039 29290 11073 29324
rect 11107 29290 11141 29324
rect 11175 29290 11209 29324
rect 11243 29290 11277 29324
rect 11311 29290 11345 29324
rect 11379 29290 11413 29324
rect 11447 29290 11481 29324
rect 11515 29290 11549 29324
rect 11583 29290 11617 29324
rect 11651 29290 11685 29324
rect 11719 29290 11753 29324
rect 11787 29290 11821 29324
rect 11855 29290 11889 29324
rect 11923 29290 11957 29324
rect 11991 29290 12025 29324
rect 12059 29290 12093 29324
rect 12127 29290 12161 29324
rect 12195 29290 12229 29324
rect 12263 29290 12297 29324
rect 12331 29290 12365 29324
rect 12399 29290 12433 29324
rect 12467 29290 12501 29324
rect 12535 29290 12569 29324
rect 12603 29290 12637 29324
rect 12671 29290 12705 29324
rect 12739 29290 12773 29324
rect 12807 29290 12841 29324
rect 12875 29290 12909 29324
rect 12943 29290 12977 29324
rect 5179 28820 5213 28854
rect 5248 28820 5282 28854
rect 5317 28820 5351 28854
rect 5386 28820 5420 28854
rect 5455 28820 5489 28854
rect 5524 28820 5558 28854
rect 5593 28820 5627 28854
rect 5662 28820 5696 28854
rect 5731 28820 5765 28854
rect 5800 28820 5834 28854
rect 5869 28820 5903 28854
rect 5938 28820 5972 28854
rect 6007 28820 6041 28854
rect 6075 28820 6109 28854
rect 6143 28820 6177 28854
rect 6211 28820 6245 28854
rect 6279 28820 6313 28854
rect 6347 28820 6381 28854
rect 6415 28820 6449 28854
rect 6483 28820 6517 28854
rect 6551 28820 6585 28854
rect 6619 28820 6653 28854
rect 6687 28820 6721 28854
rect 6755 28820 6789 28854
rect 6823 28820 6857 28854
rect 6891 28820 6925 28854
rect 6959 28820 6993 28854
rect 7027 28820 7061 28854
rect 7095 28820 7129 28854
rect 7163 28820 7197 28854
rect 7231 28820 7265 28854
rect 7299 28820 7333 28854
rect 7367 28820 7401 28854
rect 7435 28820 7469 28854
rect 7503 28820 7537 28854
rect 7571 28820 7605 28854
rect 7639 28820 7673 28854
rect 7707 28820 7741 28854
rect 7775 28820 7809 28854
rect 7843 28820 7877 28854
rect 7911 28820 7945 28854
rect 7979 28820 8013 28854
rect 8047 28820 8081 28854
rect 8115 28820 8149 28854
rect 8183 28820 8217 28854
rect 8251 28820 8285 28854
rect 8319 28820 8353 28854
rect 8387 28820 8421 28854
rect 8455 28820 8489 28854
rect 8523 28820 8557 28854
rect 8591 28820 8625 28854
rect 8659 28820 8693 28854
rect 8727 28820 8761 28854
rect 8795 28820 8829 28854
rect 8863 28820 8897 28854
rect 8931 28820 8965 28854
rect 8999 28820 9033 28854
rect 9067 28820 9101 28854
rect 9135 28820 9169 28854
rect 9203 28820 9237 28854
rect 9271 28820 9305 28854
rect 9339 28820 9373 28854
rect 9407 28820 9441 28854
rect 9475 28820 9509 28854
rect 9543 28820 9577 28854
rect 9611 28820 9645 28854
rect 9679 28820 9713 28854
rect 9747 28820 9781 28854
rect 9815 28820 9849 28854
rect 9883 28820 9917 28854
rect 9951 28820 9985 28854
rect 10019 28820 10053 28854
rect 10087 28820 10121 28854
rect 10155 28820 10189 28854
rect 10223 28820 10257 28854
rect 10291 28820 10325 28854
rect 10359 28820 10393 28854
rect 10427 28820 10461 28854
rect 10495 28820 10529 28854
rect 10563 28820 10597 28854
rect 10631 28820 10665 28854
rect 10699 28820 10733 28854
rect 10767 28820 10801 28854
rect 10835 28820 10869 28854
rect 10903 28820 10937 28854
rect 10971 28820 11005 28854
rect 11039 28820 11073 28854
rect 11107 28820 11141 28854
rect 11175 28820 11209 28854
rect 11243 28820 11277 28854
rect 11311 28820 11345 28854
rect 11379 28820 11413 28854
rect 11447 28820 11481 28854
rect 11515 28820 11549 28854
rect 11583 28820 11617 28854
rect 11651 28820 11685 28854
rect 11719 28820 11753 28854
rect 11787 28820 11821 28854
rect 11855 28820 11889 28854
rect 11923 28820 11957 28854
rect 11991 28820 12025 28854
rect 12059 28820 12093 28854
rect 12127 28820 12161 28854
rect 12195 28820 12229 28854
rect 12263 28820 12297 28854
rect 12331 28820 12365 28854
rect 12399 28820 12433 28854
rect 12467 28820 12501 28854
rect 12535 28820 12569 28854
rect 12603 28820 12637 28854
rect 12671 28820 12705 28854
rect 12739 28820 12773 28854
rect 12807 28820 12841 28854
rect 12875 28820 12909 28854
rect 12943 28820 12977 28854
rect 5179 27290 5213 27324
rect 5248 27290 5282 27324
rect 5317 27290 5351 27324
rect 5386 27290 5420 27324
rect 5455 27290 5489 27324
rect 5524 27290 5558 27324
rect 5593 27290 5627 27324
rect 5662 27290 5696 27324
rect 5731 27290 5765 27324
rect 5800 27290 5834 27324
rect 5869 27290 5903 27324
rect 5938 27290 5972 27324
rect 6007 27290 6041 27324
rect 6075 27290 6109 27324
rect 6143 27290 6177 27324
rect 6211 27290 6245 27324
rect 6279 27290 6313 27324
rect 6347 27290 6381 27324
rect 6415 27290 6449 27324
rect 6483 27290 6517 27324
rect 6551 27290 6585 27324
rect 6619 27290 6653 27324
rect 6687 27290 6721 27324
rect 6755 27290 6789 27324
rect 6823 27290 6857 27324
rect 6891 27290 6925 27324
rect 6959 27290 6993 27324
rect 7027 27290 7061 27324
rect 7095 27290 7129 27324
rect 7163 27290 7197 27324
rect 7231 27290 7265 27324
rect 7299 27290 7333 27324
rect 7367 27290 7401 27324
rect 7435 27290 7469 27324
rect 7503 27290 7537 27324
rect 7571 27290 7605 27324
rect 7639 27290 7673 27324
rect 7707 27290 7741 27324
rect 7775 27290 7809 27324
rect 7843 27290 7877 27324
rect 7911 27290 7945 27324
rect 7979 27290 8013 27324
rect 8047 27290 8081 27324
rect 8115 27290 8149 27324
rect 8183 27290 8217 27324
rect 8251 27290 8285 27324
rect 8319 27290 8353 27324
rect 8387 27290 8421 27324
rect 8455 27290 8489 27324
rect 8523 27290 8557 27324
rect 8591 27290 8625 27324
rect 8659 27290 8693 27324
rect 8727 27290 8761 27324
rect 8795 27290 8829 27324
rect 8863 27290 8897 27324
rect 8931 27290 8965 27324
rect 8999 27290 9033 27324
rect 9067 27290 9101 27324
rect 9135 27290 9169 27324
rect 9203 27290 9237 27324
rect 9271 27290 9305 27324
rect 9339 27290 9373 27324
rect 9407 27290 9441 27324
rect 9475 27290 9509 27324
rect 9543 27290 9577 27324
rect 9611 27290 9645 27324
rect 9679 27290 9713 27324
rect 9747 27290 9781 27324
rect 9815 27290 9849 27324
rect 9883 27290 9917 27324
rect 9951 27290 9985 27324
rect 10019 27290 10053 27324
rect 10087 27290 10121 27324
rect 10155 27290 10189 27324
rect 10223 27290 10257 27324
rect 10291 27290 10325 27324
rect 10359 27290 10393 27324
rect 10427 27290 10461 27324
rect 10495 27290 10529 27324
rect 10563 27290 10597 27324
rect 10631 27290 10665 27324
rect 10699 27290 10733 27324
rect 10767 27290 10801 27324
rect 10835 27290 10869 27324
rect 10903 27290 10937 27324
rect 10971 27290 11005 27324
rect 11039 27290 11073 27324
rect 11107 27290 11141 27324
rect 11175 27290 11209 27324
rect 11243 27290 11277 27324
rect 11311 27290 11345 27324
rect 11379 27290 11413 27324
rect 11447 27290 11481 27324
rect 11515 27290 11549 27324
rect 11583 27290 11617 27324
rect 11651 27290 11685 27324
rect 11719 27290 11753 27324
rect 11787 27290 11821 27324
rect 11855 27290 11889 27324
rect 11923 27290 11957 27324
rect 11991 27290 12025 27324
rect 12059 27290 12093 27324
rect 12127 27290 12161 27324
rect 12195 27290 12229 27324
rect 12263 27290 12297 27324
rect 12331 27290 12365 27324
rect 12399 27290 12433 27324
rect 12467 27290 12501 27324
rect 12535 27290 12569 27324
rect 12603 27290 12637 27324
rect 12671 27290 12705 27324
rect 12739 27290 12773 27324
rect 12807 27290 12841 27324
rect 12875 27290 12909 27324
rect 12943 27290 12977 27324
rect 5179 26820 5213 26854
rect 5248 26820 5282 26854
rect 5317 26820 5351 26854
rect 5386 26820 5420 26854
rect 5455 26820 5489 26854
rect 5524 26820 5558 26854
rect 5593 26820 5627 26854
rect 5662 26820 5696 26854
rect 5731 26820 5765 26854
rect 5800 26820 5834 26854
rect 5869 26820 5903 26854
rect 5938 26820 5972 26854
rect 6007 26820 6041 26854
rect 6075 26820 6109 26854
rect 6143 26820 6177 26854
rect 6211 26820 6245 26854
rect 6279 26820 6313 26854
rect 6347 26820 6381 26854
rect 6415 26820 6449 26854
rect 6483 26820 6517 26854
rect 6551 26820 6585 26854
rect 6619 26820 6653 26854
rect 6687 26820 6721 26854
rect 6755 26820 6789 26854
rect 6823 26820 6857 26854
rect 6891 26820 6925 26854
rect 6959 26820 6993 26854
rect 7027 26820 7061 26854
rect 7095 26820 7129 26854
rect 7163 26820 7197 26854
rect 7231 26820 7265 26854
rect 7299 26820 7333 26854
rect 7367 26820 7401 26854
rect 7435 26820 7469 26854
rect 7503 26820 7537 26854
rect 7571 26820 7605 26854
rect 7639 26820 7673 26854
rect 7707 26820 7741 26854
rect 7775 26820 7809 26854
rect 7843 26820 7877 26854
rect 7911 26820 7945 26854
rect 7979 26820 8013 26854
rect 8047 26820 8081 26854
rect 8115 26820 8149 26854
rect 8183 26820 8217 26854
rect 8251 26820 8285 26854
rect 8319 26820 8353 26854
rect 8387 26820 8421 26854
rect 8455 26820 8489 26854
rect 8523 26820 8557 26854
rect 8591 26820 8625 26854
rect 8659 26820 8693 26854
rect 8727 26820 8761 26854
rect 8795 26820 8829 26854
rect 8863 26820 8897 26854
rect 8931 26820 8965 26854
rect 8999 26820 9033 26854
rect 9067 26820 9101 26854
rect 9135 26820 9169 26854
rect 9203 26820 9237 26854
rect 9271 26820 9305 26854
rect 9339 26820 9373 26854
rect 9407 26820 9441 26854
rect 9475 26820 9509 26854
rect 9543 26820 9577 26854
rect 9611 26820 9645 26854
rect 9679 26820 9713 26854
rect 9747 26820 9781 26854
rect 9815 26820 9849 26854
rect 9883 26820 9917 26854
rect 9951 26820 9985 26854
rect 10019 26820 10053 26854
rect 10087 26820 10121 26854
rect 10155 26820 10189 26854
rect 10223 26820 10257 26854
rect 10291 26820 10325 26854
rect 10359 26820 10393 26854
rect 10427 26820 10461 26854
rect 10495 26820 10529 26854
rect 10563 26820 10597 26854
rect 10631 26820 10665 26854
rect 10699 26820 10733 26854
rect 10767 26820 10801 26854
rect 10835 26820 10869 26854
rect 10903 26820 10937 26854
rect 10971 26820 11005 26854
rect 11039 26820 11073 26854
rect 11107 26820 11141 26854
rect 11175 26820 11209 26854
rect 11243 26820 11277 26854
rect 11311 26820 11345 26854
rect 11379 26820 11413 26854
rect 11447 26820 11481 26854
rect 11515 26820 11549 26854
rect 11583 26820 11617 26854
rect 11651 26820 11685 26854
rect 11719 26820 11753 26854
rect 11787 26820 11821 26854
rect 11855 26820 11889 26854
rect 11923 26820 11957 26854
rect 11991 26820 12025 26854
rect 12059 26820 12093 26854
rect 12127 26820 12161 26854
rect 12195 26820 12229 26854
rect 12263 26820 12297 26854
rect 12331 26820 12365 26854
rect 12399 26820 12433 26854
rect 12467 26820 12501 26854
rect 12535 26820 12569 26854
rect 12603 26820 12637 26854
rect 12671 26820 12705 26854
rect 12739 26820 12773 26854
rect 12807 26820 12841 26854
rect 12875 26820 12909 26854
rect 12943 26820 12977 26854
rect 5179 25669 5213 25703
rect 5248 25669 5282 25703
rect 5317 25669 5351 25703
rect 5386 25669 5420 25703
rect 5455 25669 5489 25703
rect 5524 25669 5558 25703
rect 5593 25669 5627 25703
rect 5662 25669 5696 25703
rect 5731 25669 5765 25703
rect 5800 25669 5834 25703
rect 5869 25669 5903 25703
rect 5938 25669 5972 25703
rect 6007 25669 6041 25703
rect 6075 25669 6109 25703
rect 6143 25669 6177 25703
rect 6211 25669 6245 25703
rect 6279 25669 6313 25703
rect 6347 25669 6381 25703
rect 6415 25669 6449 25703
rect 6483 25669 6517 25703
rect 6551 25669 6585 25703
rect 6619 25669 6653 25703
rect 6687 25669 6721 25703
rect 6755 25669 6789 25703
rect 6823 25669 6857 25703
rect 6891 25669 6925 25703
rect 6959 25669 6993 25703
rect 7027 25669 7061 25703
rect 7095 25669 7129 25703
rect 7163 25669 7197 25703
rect 7231 25669 7265 25703
rect 7299 25669 7333 25703
rect 7367 25669 7401 25703
rect 7435 25669 7469 25703
rect 7503 25669 7537 25703
rect 7571 25669 7605 25703
rect 7639 25669 7673 25703
rect 7707 25669 7741 25703
rect 7775 25669 7809 25703
rect 7843 25669 7877 25703
rect 7911 25669 7945 25703
rect 7979 25669 8013 25703
rect 8047 25669 8081 25703
rect 8115 25669 8149 25703
rect 8183 25669 8217 25703
rect 8251 25669 8285 25703
rect 8319 25669 8353 25703
rect 8387 25669 8421 25703
rect 8455 25669 8489 25703
rect 8523 25669 8557 25703
rect 8591 25669 8625 25703
rect 8659 25669 8693 25703
rect 8727 25669 8761 25703
rect 8795 25669 8829 25703
rect 8863 25669 8897 25703
rect 8931 25669 8965 25703
rect 8999 25669 9033 25703
rect 9067 25669 9101 25703
rect 9135 25669 9169 25703
rect 9203 25669 9237 25703
rect 9271 25669 9305 25703
rect 9339 25669 9373 25703
rect 9407 25669 9441 25703
rect 9475 25669 9509 25703
rect 9543 25669 9577 25703
rect 9611 25669 9645 25703
rect 9679 25669 9713 25703
rect 9747 25669 9781 25703
rect 9815 25669 9849 25703
rect 9883 25669 9917 25703
rect 9951 25669 9985 25703
rect 10019 25669 10053 25703
rect 10087 25669 10121 25703
rect 10155 25669 10189 25703
rect 10223 25669 10257 25703
rect 10291 25669 10325 25703
rect 10359 25669 10393 25703
rect 10427 25669 10461 25703
rect 10495 25669 10529 25703
rect 10563 25669 10597 25703
rect 10631 25669 10665 25703
rect 10699 25669 10733 25703
rect 10767 25669 10801 25703
rect 10835 25669 10869 25703
rect 10903 25669 10937 25703
rect 10971 25669 11005 25703
rect 11039 25669 11073 25703
rect 11107 25669 11141 25703
rect 11175 25669 11209 25703
rect 11243 25669 11277 25703
rect 11311 25669 11345 25703
rect 11379 25669 11413 25703
rect 11447 25669 11481 25703
rect 11515 25669 11549 25703
rect 11583 25669 11617 25703
rect 11651 25669 11685 25703
rect 11719 25669 11753 25703
rect 11787 25669 11821 25703
rect 11855 25669 11889 25703
rect 11923 25669 11957 25703
rect 11991 25669 12025 25703
rect 12059 25669 12093 25703
rect 12127 25669 12161 25703
rect 12195 25669 12229 25703
rect 12263 25669 12297 25703
rect 12331 25669 12365 25703
rect 12399 25669 12433 25703
rect 12467 25669 12501 25703
rect 12535 25669 12569 25703
rect 12603 25669 12637 25703
rect 12671 25669 12705 25703
rect 12739 25669 12773 25703
rect 12807 25669 12841 25703
rect 12875 25669 12909 25703
rect 12943 25669 12977 25703
rect 4954 23663 4988 23697
rect 5022 23663 5056 23697
rect 5090 23663 5124 23697
rect 5158 23663 5192 23697
rect 5226 23663 5260 23697
rect 5294 23663 5328 23697
rect 5362 23663 5396 23697
rect 5430 23663 5464 23697
rect 5498 23663 5532 23697
rect 5566 23663 5600 23697
rect 5634 23663 5668 23697
rect 5702 23663 5736 23697
rect 5770 23663 5804 23697
rect 5838 23663 5872 23697
rect 5906 23663 5940 23697
rect 5974 23663 6008 23697
rect 6042 23663 6076 23697
rect 6110 23663 6144 23697
rect 6178 23663 6212 23697
rect 6246 23663 6280 23697
rect 6314 23663 6348 23697
rect 6382 23663 6416 23697
rect 6450 23663 6484 23697
rect 6518 23663 6552 23697
rect 6586 23663 6620 23697
rect 6654 23663 6688 23697
rect 6722 23663 6756 23697
rect 6790 23663 6824 23697
rect 6858 23663 6892 23697
rect 6926 23663 6960 23697
rect 6994 23663 7028 23697
rect 7062 23663 7096 23697
rect 7130 23663 7164 23697
rect 7198 23663 7232 23697
rect 7266 23663 7300 23697
rect 7334 23663 7368 23697
rect 7402 23663 7436 23697
rect 7470 23663 7504 23697
rect 7538 23663 7572 23697
rect 7606 23663 7640 23697
rect 7674 23663 7708 23697
rect 7742 23663 7776 23697
rect 7810 23663 7844 23697
rect 7878 23663 7912 23697
rect 7946 23663 7980 23697
rect 8014 23663 8048 23697
rect 8082 23663 8116 23697
rect 8150 23663 8184 23697
rect 8218 23663 8252 23697
rect 8286 23663 8320 23697
rect 8354 23663 8388 23697
rect 8422 23663 8456 23697
rect 8490 23663 8524 23697
rect 8558 23663 8592 23697
rect 8626 23663 8660 23697
rect 8694 23663 8728 23697
rect 8762 23663 8796 23697
rect 8830 23663 8864 23697
rect 8898 23663 8932 23697
rect 8966 23663 9000 23697
rect 9034 23663 9068 23697
rect 9102 23663 9136 23697
rect 9170 23663 9204 23697
rect 9238 23663 9272 23697
rect 9306 23663 9340 23697
rect 9374 23663 9408 23697
rect 9442 23663 9476 23697
rect 9510 23663 9544 23697
rect 9578 23663 9612 23697
rect 9646 23663 9680 23697
rect 9714 23663 9748 23697
rect 9782 23663 9816 23697
rect 9850 23663 9884 23697
rect 9918 23663 9952 23697
rect 9986 23663 10020 23697
rect 10054 23663 10088 23697
rect 10122 23663 10156 23697
rect 10190 23663 10224 23697
rect 10258 23663 10292 23697
rect 10326 23663 10360 23697
rect 10394 23663 10428 23697
rect 10462 23663 10496 23697
rect 10530 23663 10564 23697
rect 10598 23663 10632 23697
rect 10666 23663 10700 23697
rect 10734 23663 10768 23697
rect 10802 23663 10836 23697
rect 10870 23663 10904 23697
rect 10938 23663 10972 23697
rect 11006 23663 11040 23697
rect 11074 23663 11108 23697
rect 11142 23663 11176 23697
rect 11210 23663 11244 23697
rect 11278 23663 11312 23697
rect 11346 23663 11380 23697
rect 11414 23663 11448 23697
rect 11482 23663 11516 23697
rect 11550 23663 11584 23697
rect 11618 23663 11652 23697
rect 11686 23663 11720 23697
rect 11754 23663 11788 23697
rect 11822 23663 11856 23697
rect 11890 23663 11924 23697
rect 11958 23663 11992 23697
rect 12026 23663 12060 23697
rect 12094 23663 12128 23697
rect 12162 23663 12196 23697
rect 12230 23663 12264 23697
rect 12298 23663 12332 23697
rect 12366 23663 12400 23697
rect 12434 23663 12468 23697
rect 12502 23663 12536 23697
rect 12570 23663 12604 23697
rect 12638 23663 12672 23697
rect 12706 23663 12740 23697
rect 12774 23663 12808 23697
rect 12842 23663 12876 23697
rect 12910 23663 12944 23697
rect 12978 23663 13012 23697
rect 13046 23663 13080 23697
rect 13114 23663 13148 23697
rect 13182 23663 13216 23697
rect 13250 23663 13284 23697
rect 4954 23428 4988 23462
rect 5022 23428 5056 23462
rect 5090 23428 5124 23462
rect 5158 23428 5192 23462
rect 5226 23428 5260 23462
rect 5294 23428 5328 23462
rect 5362 23428 5396 23462
rect 5430 23428 5464 23462
rect 5498 23428 5532 23462
rect 5566 23428 5600 23462
rect 5634 23428 5668 23462
rect 5702 23428 5736 23462
rect 5770 23428 5804 23462
rect 5838 23428 5872 23462
rect 5906 23428 5940 23462
rect 5974 23428 6008 23462
rect 6042 23428 6076 23462
rect 6110 23428 6144 23462
rect 6178 23428 6212 23462
rect 6246 23428 6280 23462
rect 6314 23428 6348 23462
rect 6382 23428 6416 23462
rect 6450 23428 6484 23462
rect 6518 23428 6552 23462
rect 6586 23428 6620 23462
rect 6654 23428 6688 23462
rect 6722 23428 6756 23462
rect 6790 23428 6824 23462
rect 6858 23428 6892 23462
rect 6926 23428 6960 23462
rect 6994 23428 7028 23462
rect 7062 23428 7096 23462
rect 7130 23428 7164 23462
rect 7198 23428 7232 23462
rect 7266 23428 7300 23462
rect 7334 23428 7368 23462
rect 7402 23428 7436 23462
rect 7470 23428 7504 23462
rect 7538 23428 7572 23462
rect 7606 23428 7640 23462
rect 7674 23428 7708 23462
rect 7742 23428 7776 23462
rect 7810 23428 7844 23462
rect 7878 23428 7912 23462
rect 7946 23428 7980 23462
rect 8014 23428 8048 23462
rect 8082 23428 8116 23462
rect 8150 23428 8184 23462
rect 8218 23428 8252 23462
rect 8286 23428 8320 23462
rect 8354 23428 8388 23462
rect 8422 23428 8456 23462
rect 8490 23428 8524 23462
rect 8558 23428 8592 23462
rect 8626 23428 8660 23462
rect 8694 23428 8728 23462
rect 8762 23428 8796 23462
rect 8830 23428 8864 23462
rect 8898 23428 8932 23462
rect 8966 23428 9000 23462
rect 9034 23428 9068 23462
rect 9102 23428 9136 23462
rect 9170 23428 9204 23462
rect 9238 23428 9272 23462
rect 9306 23428 9340 23462
rect 9374 23428 9408 23462
rect 9442 23428 9476 23462
rect 9510 23428 9544 23462
rect 9578 23428 9612 23462
rect 9646 23428 9680 23462
rect 9714 23428 9748 23462
rect 9782 23428 9816 23462
rect 9850 23428 9884 23462
rect 9918 23428 9952 23462
rect 9986 23428 10020 23462
rect 10054 23428 10088 23462
rect 10122 23428 10156 23462
rect 10190 23428 10224 23462
rect 10258 23428 10292 23462
rect 10326 23428 10360 23462
rect 10394 23428 10428 23462
rect 10462 23428 10496 23462
rect 10530 23428 10564 23462
rect 10598 23428 10632 23462
rect 10666 23428 10700 23462
rect 10734 23428 10768 23462
rect 10802 23428 10836 23462
rect 10870 23428 10904 23462
rect 10938 23428 10972 23462
rect 11006 23428 11040 23462
rect 11074 23428 11108 23462
rect 11142 23428 11176 23462
rect 11210 23428 11244 23462
rect 11278 23428 11312 23462
rect 11346 23428 11380 23462
rect 11414 23428 11448 23462
rect 11482 23428 11516 23462
rect 11550 23428 11584 23462
rect 11618 23428 11652 23462
rect 11686 23428 11720 23462
rect 11754 23428 11788 23462
rect 11822 23428 11856 23462
rect 11890 23428 11924 23462
rect 11958 23428 11992 23462
rect 12026 23428 12060 23462
rect 12094 23428 12128 23462
rect 12162 23428 12196 23462
rect 12230 23428 12264 23462
rect 12298 23428 12332 23462
rect 12366 23428 12400 23462
rect 12434 23428 12468 23462
rect 12502 23428 12536 23462
rect 12570 23428 12604 23462
rect 12638 23428 12672 23462
rect 12706 23428 12740 23462
rect 12774 23428 12808 23462
rect 12842 23428 12876 23462
rect 12910 23428 12944 23462
rect 12978 23428 13012 23462
rect 13046 23428 13080 23462
rect 13114 23428 13148 23462
rect 13182 23428 13216 23462
rect 13250 23428 13284 23462
rect 4954 21729 4988 21763
rect 5022 21729 5056 21763
rect 5090 21729 5124 21763
rect 5158 21729 5192 21763
rect 5226 21729 5260 21763
rect 5294 21729 5328 21763
rect 5362 21729 5396 21763
rect 5430 21729 5464 21763
rect 5498 21729 5532 21763
rect 5566 21729 5600 21763
rect 5634 21729 5668 21763
rect 5702 21729 5736 21763
rect 5770 21729 5804 21763
rect 5838 21729 5872 21763
rect 5906 21729 5940 21763
rect 5974 21729 6008 21763
rect 6042 21729 6076 21763
rect 6110 21729 6144 21763
rect 6178 21729 6212 21763
rect 6246 21729 6280 21763
rect 6314 21729 6348 21763
rect 6382 21729 6416 21763
rect 6450 21729 6484 21763
rect 6518 21729 6552 21763
rect 6586 21729 6620 21763
rect 6654 21729 6688 21763
rect 6722 21729 6756 21763
rect 6790 21729 6824 21763
rect 6858 21729 6892 21763
rect 6926 21729 6960 21763
rect 6994 21729 7028 21763
rect 7062 21729 7096 21763
rect 7130 21729 7164 21763
rect 7198 21729 7232 21763
rect 7266 21729 7300 21763
rect 7334 21729 7368 21763
rect 7402 21729 7436 21763
rect 7470 21729 7504 21763
rect 7538 21729 7572 21763
rect 7606 21729 7640 21763
rect 7674 21729 7708 21763
rect 7742 21729 7776 21763
rect 7810 21729 7844 21763
rect 7878 21729 7912 21763
rect 7946 21729 7980 21763
rect 8014 21729 8048 21763
rect 8082 21729 8116 21763
rect 8150 21729 8184 21763
rect 8218 21729 8252 21763
rect 8286 21729 8320 21763
rect 8354 21729 8388 21763
rect 8422 21729 8456 21763
rect 8490 21729 8524 21763
rect 8558 21729 8592 21763
rect 8626 21729 8660 21763
rect 8694 21729 8728 21763
rect 8762 21729 8796 21763
rect 8830 21729 8864 21763
rect 8898 21729 8932 21763
rect 8966 21729 9000 21763
rect 9034 21729 9068 21763
rect 9102 21729 9136 21763
rect 9170 21729 9204 21763
rect 9238 21729 9272 21763
rect 9306 21729 9340 21763
rect 9374 21729 9408 21763
rect 9442 21729 9476 21763
rect 9510 21729 9544 21763
rect 9578 21729 9612 21763
rect 9646 21729 9680 21763
rect 9714 21729 9748 21763
rect 9782 21729 9816 21763
rect 9850 21729 9884 21763
rect 9918 21729 9952 21763
rect 9986 21729 10020 21763
rect 10054 21729 10088 21763
rect 10122 21729 10156 21763
rect 10190 21729 10224 21763
rect 10258 21729 10292 21763
rect 10326 21729 10360 21763
rect 10394 21729 10428 21763
rect 10462 21729 10496 21763
rect 10530 21729 10564 21763
rect 10598 21729 10632 21763
rect 10666 21729 10700 21763
rect 10734 21729 10768 21763
rect 10802 21729 10836 21763
rect 10870 21729 10904 21763
rect 10938 21729 10972 21763
rect 11006 21729 11040 21763
rect 11074 21729 11108 21763
rect 11142 21729 11176 21763
rect 11210 21729 11244 21763
rect 11278 21729 11312 21763
rect 11346 21729 11380 21763
rect 11414 21729 11448 21763
rect 11482 21729 11516 21763
rect 11550 21729 11584 21763
rect 11618 21729 11652 21763
rect 11686 21729 11720 21763
rect 11754 21729 11788 21763
rect 11822 21729 11856 21763
rect 11890 21729 11924 21763
rect 11958 21729 11992 21763
rect 12026 21729 12060 21763
rect 12094 21729 12128 21763
rect 12162 21729 12196 21763
rect 12230 21729 12264 21763
rect 12298 21729 12332 21763
rect 12366 21729 12400 21763
rect 12434 21729 12468 21763
rect 12502 21729 12536 21763
rect 12570 21729 12604 21763
rect 12638 21729 12672 21763
rect 12706 21729 12740 21763
rect 12774 21729 12808 21763
rect 12842 21729 12876 21763
rect 12910 21729 12944 21763
rect 12978 21729 13012 21763
rect 13046 21729 13080 21763
rect 13114 21729 13148 21763
rect 13182 21729 13216 21763
rect 13250 21729 13284 21763
rect 4943 19708 4977 19742
rect 5011 19708 5045 19742
rect 5079 19708 5113 19742
rect 5147 19708 5181 19742
rect 5215 19708 5249 19742
rect 5283 19708 5317 19742
rect 5351 19708 5385 19742
rect 5419 19708 5453 19742
rect 5487 19708 5521 19742
rect 5555 19708 5589 19742
rect 5623 19708 5657 19742
rect 5691 19708 5725 19742
rect 5759 19708 5793 19742
rect 5827 19708 5861 19742
rect 5895 19708 5929 19742
rect 5963 19708 5997 19742
rect 6031 19708 6065 19742
rect 6099 19708 6133 19742
rect 6167 19708 6201 19742
rect 6235 19708 6269 19742
rect 6303 19708 6337 19742
rect 6371 19708 6405 19742
rect 6439 19708 6473 19742
rect 6507 19708 6541 19742
rect 6575 19708 6609 19742
rect 6643 19708 6677 19742
rect 6711 19708 6745 19742
rect 6779 19708 6813 19742
rect 6847 19708 6881 19742
rect 6915 19708 6949 19742
rect 6983 19708 7017 19742
rect 7051 19708 7085 19742
rect 7119 19708 7153 19742
rect 7187 19708 7221 19742
rect 7255 19708 7289 19742
rect 7323 19708 7357 19742
rect 7391 19708 7425 19742
rect 7459 19708 7493 19742
rect 7527 19708 7561 19742
rect 7595 19708 7629 19742
rect 7663 19708 7697 19742
rect 7731 19708 7765 19742
rect 7799 19708 7833 19742
rect 7867 19708 7901 19742
rect 7935 19708 7969 19742
rect 8003 19708 8037 19742
rect 8071 19708 8105 19742
rect 8139 19708 8173 19742
rect 8207 19708 8241 19742
rect 8275 19708 8309 19742
rect 8343 19708 8377 19742
rect 8411 19708 8445 19742
rect 8479 19708 8513 19742
rect 8547 19708 8581 19742
rect 8615 19708 8649 19742
rect 8683 19708 8717 19742
rect 8751 19708 8785 19742
rect 8819 19708 8853 19742
rect 8887 19708 8921 19742
rect 8955 19708 8989 19742
rect 9023 19708 9057 19742
rect 9091 19708 9125 19742
rect 9159 19708 9193 19742
rect 9227 19708 9261 19742
rect 9295 19708 9329 19742
rect 9363 19708 9397 19742
rect 9431 19708 9465 19742
rect 9499 19708 9533 19742
rect 9567 19708 9601 19742
rect 9635 19708 9669 19742
rect 9703 19708 9737 19742
rect 9771 19708 9805 19742
rect 9839 19708 9873 19742
rect 9907 19708 9941 19742
rect 9975 19708 10009 19742
rect 10043 19708 10077 19742
rect 10111 19708 10145 19742
rect 10179 19708 10213 19742
rect 10247 19708 10281 19742
rect 10315 19708 10349 19742
rect 10383 19708 10417 19742
rect 10451 19708 10485 19742
rect 10519 19708 10553 19742
rect 10587 19708 10621 19742
rect 10655 19708 10689 19742
rect 10723 19708 10757 19742
rect 10791 19708 10825 19742
rect 10859 19708 10893 19742
rect 10927 19708 10961 19742
rect 10995 19708 11029 19742
rect 11063 19708 11097 19742
rect 11131 19708 11165 19742
rect 11199 19708 11233 19742
rect 11267 19708 11301 19742
rect 11335 19708 11369 19742
rect 11403 19708 11437 19742
rect 11471 19708 11505 19742
rect 11539 19708 11573 19742
rect 11607 19708 11641 19742
rect 11675 19708 11709 19742
rect 11743 19708 11777 19742
rect 11811 19708 11845 19742
rect 11879 19708 11913 19742
rect 11947 19708 11981 19742
rect 12015 19708 12049 19742
rect 12083 19708 12117 19742
rect 12151 19708 12185 19742
rect 12219 19708 12253 19742
rect 12287 19708 12321 19742
rect 12355 19708 12389 19742
rect 12423 19708 12457 19742
rect 12491 19708 12525 19742
rect 12559 19708 12593 19742
rect 12627 19708 12661 19742
rect 12695 19708 12729 19742
rect 12763 19708 12797 19742
rect 12831 19708 12865 19742
rect 12899 19708 12933 19742
rect 12967 19708 13001 19742
rect 13035 19708 13069 19742
rect 13103 19708 13137 19742
rect 13171 19708 13205 19742
rect 13239 19708 13273 19742
rect 4943 18009 4977 18043
rect 5011 18009 5045 18043
rect 5079 18009 5113 18043
rect 5147 18009 5181 18043
rect 5215 18009 5249 18043
rect 5283 18009 5317 18043
rect 5351 18009 5385 18043
rect 5419 18009 5453 18043
rect 5487 18009 5521 18043
rect 5555 18009 5589 18043
rect 5623 18009 5657 18043
rect 5691 18009 5725 18043
rect 5759 18009 5793 18043
rect 5827 18009 5861 18043
rect 5895 18009 5929 18043
rect 5963 18009 5997 18043
rect 6031 18009 6065 18043
rect 6099 18009 6133 18043
rect 6167 18009 6201 18043
rect 6235 18009 6269 18043
rect 6303 18009 6337 18043
rect 6371 18009 6405 18043
rect 6439 18009 6473 18043
rect 6507 18009 6541 18043
rect 6575 18009 6609 18043
rect 6643 18009 6677 18043
rect 6711 18009 6745 18043
rect 6779 18009 6813 18043
rect 6847 18009 6881 18043
rect 6915 18009 6949 18043
rect 6983 18009 7017 18043
rect 7051 18009 7085 18043
rect 7119 18009 7153 18043
rect 7187 18009 7221 18043
rect 7255 18009 7289 18043
rect 7323 18009 7357 18043
rect 7391 18009 7425 18043
rect 7459 18009 7493 18043
rect 7527 18009 7561 18043
rect 7595 18009 7629 18043
rect 7663 18009 7697 18043
rect 7731 18009 7765 18043
rect 7799 18009 7833 18043
rect 7867 18009 7901 18043
rect 7935 18009 7969 18043
rect 8003 18009 8037 18043
rect 8071 18009 8105 18043
rect 8139 18009 8173 18043
rect 8207 18009 8241 18043
rect 8275 18009 8309 18043
rect 8343 18009 8377 18043
rect 8411 18009 8445 18043
rect 8479 18009 8513 18043
rect 8547 18009 8581 18043
rect 8615 18009 8649 18043
rect 8683 18009 8717 18043
rect 8751 18009 8785 18043
rect 8819 18009 8853 18043
rect 8887 18009 8921 18043
rect 8955 18009 8989 18043
rect 9023 18009 9057 18043
rect 9091 18009 9125 18043
rect 9159 18009 9193 18043
rect 9227 18009 9261 18043
rect 9295 18009 9329 18043
rect 9363 18009 9397 18043
rect 9431 18009 9465 18043
rect 9499 18009 9533 18043
rect 9567 18009 9601 18043
rect 9635 18009 9669 18043
rect 9703 18009 9737 18043
rect 9771 18009 9805 18043
rect 9839 18009 9873 18043
rect 9907 18009 9941 18043
rect 9975 18009 10009 18043
rect 10043 18009 10077 18043
rect 10111 18009 10145 18043
rect 10179 18009 10213 18043
rect 10247 18009 10281 18043
rect 10315 18009 10349 18043
rect 10383 18009 10417 18043
rect 10451 18009 10485 18043
rect 10519 18009 10553 18043
rect 10587 18009 10621 18043
rect 10655 18009 10689 18043
rect 10723 18009 10757 18043
rect 10791 18009 10825 18043
rect 10859 18009 10893 18043
rect 10927 18009 10961 18043
rect 10995 18009 11029 18043
rect 11063 18009 11097 18043
rect 11131 18009 11165 18043
rect 11199 18009 11233 18043
rect 11267 18009 11301 18043
rect 11335 18009 11369 18043
rect 11403 18009 11437 18043
rect 11471 18009 11505 18043
rect 11539 18009 11573 18043
rect 11607 18009 11641 18043
rect 11675 18009 11709 18043
rect 11743 18009 11777 18043
rect 11811 18009 11845 18043
rect 11879 18009 11913 18043
rect 11947 18009 11981 18043
rect 12015 18009 12049 18043
rect 12083 18009 12117 18043
rect 12151 18009 12185 18043
rect 12219 18009 12253 18043
rect 12287 18009 12321 18043
rect 12355 18009 12389 18043
rect 12423 18009 12457 18043
rect 12491 18009 12525 18043
rect 12559 18009 12593 18043
rect 12627 18009 12661 18043
rect 12695 18009 12729 18043
rect 12763 18009 12797 18043
rect 12831 18009 12865 18043
rect 12899 18009 12933 18043
rect 12967 18009 13001 18043
rect 13035 18009 13069 18043
rect 13103 18009 13137 18043
rect 13171 18009 13205 18043
rect 13239 18009 13273 18043
rect 2615 16209 2649 16243
rect 2683 16209 2717 16243
rect 2751 16209 2785 16243
rect 2819 16209 2853 16243
rect 2887 16209 2921 16243
rect 2955 16209 2989 16243
rect 3023 16209 3057 16243
rect 3091 16209 3125 16243
rect 3159 16209 3193 16243
rect 3227 16209 3261 16243
rect 3295 16209 3329 16243
rect 3363 16209 3397 16243
rect 3431 16209 3465 16243
rect 3499 16209 3533 16243
rect 3567 16209 3601 16243
rect 3635 16209 3669 16243
rect 3703 16209 3737 16243
rect 3771 16209 3805 16243
rect 3839 16209 3873 16243
rect 3907 16209 3941 16243
rect 3975 16209 4009 16243
rect 4043 16209 4077 16243
rect 4111 16209 4145 16243
rect 4179 16209 4213 16243
rect 4247 16209 4281 16243
rect 4315 16209 4349 16243
rect 4383 16209 4417 16243
rect 4451 16209 4485 16243
rect 4519 16209 4553 16243
rect 4587 16209 4621 16243
rect 4655 16209 4689 16243
rect 4723 16209 4757 16243
rect 4791 16209 4825 16243
rect 4859 16209 4893 16243
rect 4927 16209 4961 16243
rect 4995 16209 5029 16243
rect 5063 16209 5097 16243
rect 5131 16209 5165 16243
rect 5199 16209 5233 16243
rect 5267 16209 5301 16243
rect 5335 16209 5369 16243
rect 5403 16209 5437 16243
rect 5471 16209 5505 16243
rect 5539 16209 5573 16243
rect 5607 16209 5641 16243
rect 5675 16209 5709 16243
rect 5743 16209 5777 16243
rect 5811 16209 5845 16243
rect 5879 16209 5913 16243
rect 5947 16209 5981 16243
rect 6015 16209 6049 16243
rect 6083 16209 6117 16243
rect 6151 16209 6185 16243
rect 6219 16209 6253 16243
rect 6287 16209 6321 16243
rect 6355 16209 6389 16243
rect 6423 16209 6457 16243
rect 6491 16209 6525 16243
rect 6559 16209 6593 16243
rect 6627 16209 6661 16243
rect 6695 16209 6729 16243
rect 6763 16209 6797 16243
rect 6831 16209 6865 16243
rect 6899 16209 6933 16243
rect 6967 16209 7001 16243
rect 7035 16209 7069 16243
rect 7103 16209 7137 16243
rect 7171 16209 7205 16243
rect 7239 16209 7273 16243
rect 7307 16209 7341 16243
rect 7375 16209 7409 16243
rect 7443 16209 7477 16243
rect 7511 16209 7545 16243
rect 7579 16209 7613 16243
rect 7647 16209 7681 16243
rect 7715 16209 7749 16243
rect 7783 16209 7817 16243
rect 7851 16209 7885 16243
rect 7919 16209 7953 16243
rect 7987 16209 8021 16243
rect 8055 16209 8089 16243
rect 8123 16209 8157 16243
rect 8191 16209 8225 16243
rect 8259 16209 8293 16243
rect 8327 16209 8361 16243
rect 8395 16209 8429 16243
rect 8463 16209 8497 16243
rect 8531 16209 8565 16243
rect 8599 16209 8633 16243
rect 8667 16209 8701 16243
rect 8735 16209 8769 16243
rect 8803 16209 8837 16243
rect 8871 16209 8905 16243
rect 8939 16209 8973 16243
rect 9007 16209 9041 16243
rect 9075 16209 9109 16243
rect 9143 16209 9177 16243
rect 9211 16209 9245 16243
rect 9279 16209 9313 16243
rect 9347 16209 9381 16243
rect 9415 16209 9449 16243
rect 9483 16209 9517 16243
rect 9551 16209 9585 16243
rect 9619 16209 9653 16243
rect 9687 16209 9721 16243
rect 9755 16209 9789 16243
rect 9823 16209 9857 16243
rect 9891 16209 9925 16243
rect 9959 16209 9993 16243
rect 10027 16209 10061 16243
rect 10095 16209 10129 16243
rect 10163 16209 10197 16243
rect 10231 16209 10265 16243
rect 10299 16209 10333 16243
rect 10367 16209 10401 16243
rect 10435 16209 10469 16243
rect 10503 16209 10537 16243
rect 10571 16209 10605 16243
rect 10639 16209 10673 16243
rect 10707 16209 10741 16243
rect 10775 16209 10809 16243
rect 10843 16209 10877 16243
rect 10911 16209 10945 16243
rect 10979 16209 11013 16243
rect 11047 16209 11081 16243
rect 11115 16209 11149 16243
rect 11183 16209 11217 16243
rect 11251 16209 11285 16243
rect 11319 16209 11353 16243
rect 11387 16209 11421 16243
rect 11455 16209 11489 16243
rect 11523 16209 11557 16243
rect 11591 16209 11625 16243
rect 11659 16209 11693 16243
rect 11727 16209 11761 16243
rect 11795 16209 11829 16243
rect 11863 16209 11897 16243
rect 11931 16209 11965 16243
rect 11999 16209 12033 16243
rect 12067 16209 12101 16243
rect 12135 16209 12169 16243
rect 12203 16209 12237 16243
rect 12271 16209 12305 16243
rect 12339 16209 12373 16243
rect 12407 16209 12441 16243
rect 12475 16209 12509 16243
rect 12543 16209 12577 16243
rect 12611 16209 12645 16243
rect 12679 16209 12713 16243
rect 12747 16209 12781 16243
rect 12815 16209 12849 16243
rect 12883 16209 12917 16243
rect 12951 16209 12985 16243
rect 13019 16209 13053 16243
rect 13087 16209 13121 16243
rect 13155 16209 13189 16243
rect 13223 16209 13257 16243
rect 2888 13290 2922 13324
rect 2957 13290 2991 13324
rect 3026 13290 3060 13324
rect 3095 13290 3129 13324
rect 3164 13290 3198 13324
rect 3233 13290 3267 13324
rect 3302 13290 3336 13324
rect 3371 13290 3405 13324
rect 3440 13290 3474 13324
rect 3509 13290 3543 13324
rect 3578 13290 3612 13324
rect 3647 13290 3681 13324
rect 3716 13290 3750 13324
rect 3785 13290 3819 13324
rect 3854 13290 3888 13324
rect 3923 13290 3957 13324
rect 3992 13290 4026 13324
rect 4061 13290 4095 13324
rect 4130 13290 4164 13324
rect 4199 13290 4233 13324
rect 4268 13290 4302 13324
rect 4337 13290 4371 13324
rect 4406 13290 4440 13324
rect 4475 13290 4509 13324
rect 4544 13290 4578 13324
rect 4613 13290 4647 13324
rect 4682 13290 4716 13324
rect 4751 13290 4785 13324
rect 4820 13290 4854 13324
rect 4889 13290 4923 13324
rect 4958 13290 4992 13324
rect 5027 13290 5061 13324
rect 5096 13290 5130 13324
rect 5165 13290 5199 13324
rect 5234 13290 5268 13324
rect 5303 13290 5337 13324
rect 5372 13290 5406 13324
rect 5441 13290 5475 13324
rect 5510 13290 5544 13324
rect 5579 13290 5613 13324
rect 5648 13290 5682 13324
rect 5717 13290 5751 13324
rect 5786 13290 5820 13324
rect 5855 13290 5889 13324
rect 5924 13290 5958 13324
rect 5993 13290 6027 13324
rect 6062 13290 6096 13324
rect 6131 13290 6165 13324
rect 6200 13290 6234 13324
rect 6268 13290 6302 13324
rect 6336 13290 6370 13324
rect 6404 13290 6438 13324
rect 6472 13290 6506 13324
rect 6540 13290 6574 13324
rect 6608 13290 6642 13324
rect 6676 13290 6710 13324
rect 6744 13290 6778 13324
rect 6812 13290 6846 13324
rect 6880 13290 6914 13324
rect 6948 13290 6982 13324
rect 7016 13290 7050 13324
rect 7084 13290 7118 13324
rect 7152 13290 7186 13324
rect 7220 13290 7254 13324
rect 7288 13290 7322 13324
rect 7356 13290 7390 13324
rect 7424 13290 7458 13324
rect 7492 13290 7526 13324
rect 7560 13290 7594 13324
rect 7628 13290 7662 13324
rect 7696 13290 7730 13324
rect 7764 13290 7798 13324
rect 7832 13290 7866 13324
rect 7900 13290 7934 13324
rect 7968 13290 8002 13324
rect 8036 13290 8070 13324
rect 8104 13290 8138 13324
rect 8172 13290 8206 13324
rect 8240 13290 8274 13324
rect 8308 13290 8342 13324
rect 8376 13290 8410 13324
rect 8444 13290 8478 13324
rect 8512 13290 8546 13324
rect 8580 13290 8614 13324
rect 8648 13290 8682 13324
rect 8716 13290 8750 13324
rect 8784 13290 8818 13324
rect 8852 13290 8886 13324
rect 8920 13290 8954 13324
rect 8988 13290 9022 13324
rect 9056 13290 9090 13324
rect 9124 13290 9158 13324
rect 9192 13290 9226 13324
rect 9260 13290 9294 13324
rect 9328 13290 9362 13324
rect 9396 13290 9430 13324
rect 9464 13290 9498 13324
rect 9532 13290 9566 13324
rect 9600 13290 9634 13324
rect 9668 13290 9702 13324
rect 9736 13290 9770 13324
rect 9804 13290 9838 13324
rect 9872 13290 9906 13324
rect 9940 13290 9974 13324
rect 10008 13290 10042 13324
rect 10076 13290 10110 13324
rect 10144 13290 10178 13324
rect 10212 13290 10246 13324
rect 10280 13290 10314 13324
rect 10348 13290 10382 13324
rect 10416 13290 10450 13324
rect 10484 13290 10518 13324
rect 10552 13290 10586 13324
rect 10620 13290 10654 13324
rect 10688 13290 10722 13324
rect 10756 13290 10790 13324
rect 10824 13290 10858 13324
rect 10892 13290 10926 13324
rect 10960 13290 10994 13324
rect 11028 13290 11062 13324
rect 11096 13290 11130 13324
rect 11164 13290 11198 13324
rect 11232 13290 11266 13324
rect 11300 13290 11334 13324
rect 11368 13290 11402 13324
rect 11436 13290 11470 13324
rect 11504 13290 11538 13324
rect 11572 13290 11606 13324
rect 11640 13290 11674 13324
rect 11708 13290 11742 13324
rect 11776 13290 11810 13324
rect 11844 13290 11878 13324
rect 11912 13290 11946 13324
rect 11980 13290 12014 13324
rect 12048 13290 12082 13324
rect 12116 13290 12150 13324
rect 12184 13290 12218 13324
rect 12252 13290 12286 13324
rect 12320 13290 12354 13324
rect 12388 13290 12422 13324
rect 12456 13290 12490 13324
rect 12524 13290 12558 13324
rect 12592 13290 12626 13324
rect 12660 13290 12694 13324
rect 12728 13290 12762 13324
rect 12796 13290 12830 13324
rect 12864 13290 12898 13324
rect 12932 13290 12966 13324
rect 13000 13290 13034 13324
rect 13068 13290 13102 13324
rect 2888 12820 2922 12854
rect 2957 12820 2991 12854
rect 3026 12820 3060 12854
rect 3095 12820 3129 12854
rect 3164 12820 3198 12854
rect 3233 12820 3267 12854
rect 3302 12820 3336 12854
rect 3371 12820 3405 12854
rect 3440 12820 3474 12854
rect 3509 12820 3543 12854
rect 3578 12820 3612 12854
rect 3647 12820 3681 12854
rect 3716 12820 3750 12854
rect 3785 12820 3819 12854
rect 3854 12820 3888 12854
rect 3923 12820 3957 12854
rect 3992 12820 4026 12854
rect 4061 12820 4095 12854
rect 4130 12820 4164 12854
rect 4199 12820 4233 12854
rect 4268 12820 4302 12854
rect 4337 12820 4371 12854
rect 4406 12820 4440 12854
rect 4475 12820 4509 12854
rect 4544 12820 4578 12854
rect 4613 12820 4647 12854
rect 4682 12820 4716 12854
rect 4751 12820 4785 12854
rect 4820 12820 4854 12854
rect 4889 12820 4923 12854
rect 4958 12820 4992 12854
rect 5027 12820 5061 12854
rect 5096 12820 5130 12854
rect 5165 12820 5199 12854
rect 5234 12820 5268 12854
rect 5303 12820 5337 12854
rect 5372 12820 5406 12854
rect 5441 12820 5475 12854
rect 5510 12820 5544 12854
rect 5579 12820 5613 12854
rect 5648 12820 5682 12854
rect 5717 12820 5751 12854
rect 5786 12820 5820 12854
rect 5855 12820 5889 12854
rect 5924 12820 5958 12854
rect 5993 12820 6027 12854
rect 6062 12820 6096 12854
rect 6131 12820 6165 12854
rect 6200 12820 6234 12854
rect 6268 12820 6302 12854
rect 6336 12820 6370 12854
rect 6404 12820 6438 12854
rect 6472 12820 6506 12854
rect 6540 12820 6574 12854
rect 6608 12820 6642 12854
rect 6676 12820 6710 12854
rect 6744 12820 6778 12854
rect 6812 12820 6846 12854
rect 6880 12820 6914 12854
rect 6948 12820 6982 12854
rect 7016 12820 7050 12854
rect 7084 12820 7118 12854
rect 7152 12820 7186 12854
rect 7220 12820 7254 12854
rect 7288 12820 7322 12854
rect 7356 12820 7390 12854
rect 7424 12820 7458 12854
rect 7492 12820 7526 12854
rect 7560 12820 7594 12854
rect 7628 12820 7662 12854
rect 7696 12820 7730 12854
rect 7764 12820 7798 12854
rect 7832 12820 7866 12854
rect 7900 12820 7934 12854
rect 7968 12820 8002 12854
rect 8036 12820 8070 12854
rect 8104 12820 8138 12854
rect 8172 12820 8206 12854
rect 8240 12820 8274 12854
rect 8308 12820 8342 12854
rect 8376 12820 8410 12854
rect 8444 12820 8478 12854
rect 8512 12820 8546 12854
rect 8580 12820 8614 12854
rect 8648 12820 8682 12854
rect 8716 12820 8750 12854
rect 8784 12820 8818 12854
rect 8852 12820 8886 12854
rect 8920 12820 8954 12854
rect 8988 12820 9022 12854
rect 9056 12820 9090 12854
rect 9124 12820 9158 12854
rect 9192 12820 9226 12854
rect 9260 12820 9294 12854
rect 9328 12820 9362 12854
rect 9396 12820 9430 12854
rect 9464 12820 9498 12854
rect 9532 12820 9566 12854
rect 9600 12820 9634 12854
rect 9668 12820 9702 12854
rect 9736 12820 9770 12854
rect 9804 12820 9838 12854
rect 9872 12820 9906 12854
rect 9940 12820 9974 12854
rect 10008 12820 10042 12854
rect 10076 12820 10110 12854
rect 10144 12820 10178 12854
rect 10212 12820 10246 12854
rect 10280 12820 10314 12854
rect 10348 12820 10382 12854
rect 10416 12820 10450 12854
rect 10484 12820 10518 12854
rect 10552 12820 10586 12854
rect 10620 12820 10654 12854
rect 10688 12820 10722 12854
rect 10756 12820 10790 12854
rect 10824 12820 10858 12854
rect 10892 12820 10926 12854
rect 10960 12820 10994 12854
rect 11028 12820 11062 12854
rect 11096 12820 11130 12854
rect 11164 12820 11198 12854
rect 11232 12820 11266 12854
rect 11300 12820 11334 12854
rect 11368 12820 11402 12854
rect 11436 12820 11470 12854
rect 11504 12820 11538 12854
rect 11572 12820 11606 12854
rect 11640 12820 11674 12854
rect 11708 12820 11742 12854
rect 11776 12820 11810 12854
rect 11844 12820 11878 12854
rect 11912 12820 11946 12854
rect 11980 12820 12014 12854
rect 12048 12820 12082 12854
rect 12116 12820 12150 12854
rect 12184 12820 12218 12854
rect 12252 12820 12286 12854
rect 12320 12820 12354 12854
rect 12388 12820 12422 12854
rect 12456 12820 12490 12854
rect 12524 12820 12558 12854
rect 12592 12820 12626 12854
rect 12660 12820 12694 12854
rect 12728 12820 12762 12854
rect 12796 12820 12830 12854
rect 12864 12820 12898 12854
rect 12932 12820 12966 12854
rect 13000 12820 13034 12854
rect 13068 12820 13102 12854
rect 2888 11290 2922 11324
rect 2957 11290 2991 11324
rect 3026 11290 3060 11324
rect 3095 11290 3129 11324
rect 3164 11290 3198 11324
rect 3233 11290 3267 11324
rect 3302 11290 3336 11324
rect 3371 11290 3405 11324
rect 3440 11290 3474 11324
rect 3509 11290 3543 11324
rect 3578 11290 3612 11324
rect 3647 11290 3681 11324
rect 3716 11290 3750 11324
rect 3785 11290 3819 11324
rect 3854 11290 3888 11324
rect 3923 11290 3957 11324
rect 3992 11290 4026 11324
rect 4061 11290 4095 11324
rect 4130 11290 4164 11324
rect 4199 11290 4233 11324
rect 4268 11290 4302 11324
rect 4337 11290 4371 11324
rect 4406 11290 4440 11324
rect 4475 11290 4509 11324
rect 4544 11290 4578 11324
rect 4613 11290 4647 11324
rect 4682 11290 4716 11324
rect 4751 11290 4785 11324
rect 4820 11290 4854 11324
rect 4889 11290 4923 11324
rect 4958 11290 4992 11324
rect 5027 11290 5061 11324
rect 5096 11290 5130 11324
rect 5165 11290 5199 11324
rect 5234 11290 5268 11324
rect 5303 11290 5337 11324
rect 5372 11290 5406 11324
rect 5441 11290 5475 11324
rect 5510 11290 5544 11324
rect 5579 11290 5613 11324
rect 5648 11290 5682 11324
rect 5717 11290 5751 11324
rect 5786 11290 5820 11324
rect 5855 11290 5889 11324
rect 5924 11290 5958 11324
rect 5993 11290 6027 11324
rect 6062 11290 6096 11324
rect 6131 11290 6165 11324
rect 6200 11290 6234 11324
rect 6268 11290 6302 11324
rect 6336 11290 6370 11324
rect 6404 11290 6438 11324
rect 6472 11290 6506 11324
rect 6540 11290 6574 11324
rect 6608 11290 6642 11324
rect 6676 11290 6710 11324
rect 6744 11290 6778 11324
rect 6812 11290 6846 11324
rect 6880 11290 6914 11324
rect 6948 11290 6982 11324
rect 7016 11290 7050 11324
rect 7084 11290 7118 11324
rect 7152 11290 7186 11324
rect 7220 11290 7254 11324
rect 7288 11290 7322 11324
rect 7356 11290 7390 11324
rect 7424 11290 7458 11324
rect 7492 11290 7526 11324
rect 7560 11290 7594 11324
rect 7628 11290 7662 11324
rect 7696 11290 7730 11324
rect 7764 11290 7798 11324
rect 7832 11290 7866 11324
rect 7900 11290 7934 11324
rect 7968 11290 8002 11324
rect 8036 11290 8070 11324
rect 8104 11290 8138 11324
rect 8172 11290 8206 11324
rect 8240 11290 8274 11324
rect 8308 11290 8342 11324
rect 8376 11290 8410 11324
rect 8444 11290 8478 11324
rect 8512 11290 8546 11324
rect 8580 11290 8614 11324
rect 8648 11290 8682 11324
rect 8716 11290 8750 11324
rect 8784 11290 8818 11324
rect 8852 11290 8886 11324
rect 8920 11290 8954 11324
rect 8988 11290 9022 11324
rect 9056 11290 9090 11324
rect 9124 11290 9158 11324
rect 9192 11290 9226 11324
rect 9260 11290 9294 11324
rect 9328 11290 9362 11324
rect 9396 11290 9430 11324
rect 9464 11290 9498 11324
rect 9532 11290 9566 11324
rect 9600 11290 9634 11324
rect 9668 11290 9702 11324
rect 9736 11290 9770 11324
rect 9804 11290 9838 11324
rect 9872 11290 9906 11324
rect 9940 11290 9974 11324
rect 10008 11290 10042 11324
rect 10076 11290 10110 11324
rect 10144 11290 10178 11324
rect 10212 11290 10246 11324
rect 10280 11290 10314 11324
rect 10348 11290 10382 11324
rect 10416 11290 10450 11324
rect 10484 11290 10518 11324
rect 10552 11290 10586 11324
rect 10620 11290 10654 11324
rect 10688 11290 10722 11324
rect 10756 11290 10790 11324
rect 10824 11290 10858 11324
rect 10892 11290 10926 11324
rect 10960 11290 10994 11324
rect 11028 11290 11062 11324
rect 11096 11290 11130 11324
rect 11164 11290 11198 11324
rect 11232 11290 11266 11324
rect 11300 11290 11334 11324
rect 11368 11290 11402 11324
rect 11436 11290 11470 11324
rect 11504 11290 11538 11324
rect 11572 11290 11606 11324
rect 11640 11290 11674 11324
rect 11708 11290 11742 11324
rect 11776 11290 11810 11324
rect 11844 11290 11878 11324
rect 11912 11290 11946 11324
rect 11980 11290 12014 11324
rect 12048 11290 12082 11324
rect 12116 11290 12150 11324
rect 12184 11290 12218 11324
rect 12252 11290 12286 11324
rect 12320 11290 12354 11324
rect 12388 11290 12422 11324
rect 12456 11290 12490 11324
rect 12524 11290 12558 11324
rect 12592 11290 12626 11324
rect 12660 11290 12694 11324
rect 12728 11290 12762 11324
rect 12796 11290 12830 11324
rect 12864 11290 12898 11324
rect 12932 11290 12966 11324
rect 13000 11290 13034 11324
rect 13068 11290 13102 11324
rect 2888 10820 2922 10854
rect 2957 10820 2991 10854
rect 3026 10820 3060 10854
rect 3095 10820 3129 10854
rect 3164 10820 3198 10854
rect 3233 10820 3267 10854
rect 3302 10820 3336 10854
rect 3371 10820 3405 10854
rect 3440 10820 3474 10854
rect 3509 10820 3543 10854
rect 3578 10820 3612 10854
rect 3647 10820 3681 10854
rect 3716 10820 3750 10854
rect 3785 10820 3819 10854
rect 3854 10820 3888 10854
rect 3923 10820 3957 10854
rect 3992 10820 4026 10854
rect 4061 10820 4095 10854
rect 4130 10820 4164 10854
rect 4199 10820 4233 10854
rect 4268 10820 4302 10854
rect 4337 10820 4371 10854
rect 4406 10820 4440 10854
rect 4475 10820 4509 10854
rect 4544 10820 4578 10854
rect 4613 10820 4647 10854
rect 4682 10820 4716 10854
rect 4751 10820 4785 10854
rect 4820 10820 4854 10854
rect 4889 10820 4923 10854
rect 4958 10820 4992 10854
rect 5027 10820 5061 10854
rect 5096 10820 5130 10854
rect 5165 10820 5199 10854
rect 5234 10820 5268 10854
rect 5303 10820 5337 10854
rect 5372 10820 5406 10854
rect 5441 10820 5475 10854
rect 5510 10820 5544 10854
rect 5579 10820 5613 10854
rect 5648 10820 5682 10854
rect 5717 10820 5751 10854
rect 5786 10820 5820 10854
rect 5855 10820 5889 10854
rect 5924 10820 5958 10854
rect 5993 10820 6027 10854
rect 6062 10820 6096 10854
rect 6131 10820 6165 10854
rect 6200 10820 6234 10854
rect 6268 10820 6302 10854
rect 6336 10820 6370 10854
rect 6404 10820 6438 10854
rect 6472 10820 6506 10854
rect 6540 10820 6574 10854
rect 6608 10820 6642 10854
rect 6676 10820 6710 10854
rect 6744 10820 6778 10854
rect 6812 10820 6846 10854
rect 6880 10820 6914 10854
rect 6948 10820 6982 10854
rect 7016 10820 7050 10854
rect 7084 10820 7118 10854
rect 7152 10820 7186 10854
rect 7220 10820 7254 10854
rect 7288 10820 7322 10854
rect 7356 10820 7390 10854
rect 7424 10820 7458 10854
rect 7492 10820 7526 10854
rect 7560 10820 7594 10854
rect 7628 10820 7662 10854
rect 7696 10820 7730 10854
rect 7764 10820 7798 10854
rect 7832 10820 7866 10854
rect 7900 10820 7934 10854
rect 7968 10820 8002 10854
rect 8036 10820 8070 10854
rect 8104 10820 8138 10854
rect 8172 10820 8206 10854
rect 8240 10820 8274 10854
rect 8308 10820 8342 10854
rect 8376 10820 8410 10854
rect 8444 10820 8478 10854
rect 8512 10820 8546 10854
rect 8580 10820 8614 10854
rect 8648 10820 8682 10854
rect 8716 10820 8750 10854
rect 8784 10820 8818 10854
rect 8852 10820 8886 10854
rect 8920 10820 8954 10854
rect 8988 10820 9022 10854
rect 9056 10820 9090 10854
rect 9124 10820 9158 10854
rect 9192 10820 9226 10854
rect 9260 10820 9294 10854
rect 9328 10820 9362 10854
rect 9396 10820 9430 10854
rect 9464 10820 9498 10854
rect 9532 10820 9566 10854
rect 9600 10820 9634 10854
rect 9668 10820 9702 10854
rect 9736 10820 9770 10854
rect 9804 10820 9838 10854
rect 9872 10820 9906 10854
rect 9940 10820 9974 10854
rect 10008 10820 10042 10854
rect 10076 10820 10110 10854
rect 10144 10820 10178 10854
rect 10212 10820 10246 10854
rect 10280 10820 10314 10854
rect 10348 10820 10382 10854
rect 10416 10820 10450 10854
rect 10484 10820 10518 10854
rect 10552 10820 10586 10854
rect 10620 10820 10654 10854
rect 10688 10820 10722 10854
rect 10756 10820 10790 10854
rect 10824 10820 10858 10854
rect 10892 10820 10926 10854
rect 10960 10820 10994 10854
rect 11028 10820 11062 10854
rect 11096 10820 11130 10854
rect 11164 10820 11198 10854
rect 11232 10820 11266 10854
rect 11300 10820 11334 10854
rect 11368 10820 11402 10854
rect 11436 10820 11470 10854
rect 11504 10820 11538 10854
rect 11572 10820 11606 10854
rect 11640 10820 11674 10854
rect 11708 10820 11742 10854
rect 11776 10820 11810 10854
rect 11844 10820 11878 10854
rect 11912 10820 11946 10854
rect 11980 10820 12014 10854
rect 12048 10820 12082 10854
rect 12116 10820 12150 10854
rect 12184 10820 12218 10854
rect 12252 10820 12286 10854
rect 12320 10820 12354 10854
rect 12388 10820 12422 10854
rect 12456 10820 12490 10854
rect 12524 10820 12558 10854
rect 12592 10820 12626 10854
rect 12660 10820 12694 10854
rect 12728 10820 12762 10854
rect 12796 10820 12830 10854
rect 12864 10820 12898 10854
rect 12932 10820 12966 10854
rect 13000 10820 13034 10854
rect 13068 10820 13102 10854
rect 2888 9290 2922 9324
rect 2957 9290 2991 9324
rect 3026 9290 3060 9324
rect 3095 9290 3129 9324
rect 3164 9290 3198 9324
rect 3233 9290 3267 9324
rect 3302 9290 3336 9324
rect 3371 9290 3405 9324
rect 3440 9290 3474 9324
rect 3509 9290 3543 9324
rect 3578 9290 3612 9324
rect 3647 9290 3681 9324
rect 3716 9290 3750 9324
rect 3785 9290 3819 9324
rect 3854 9290 3888 9324
rect 3923 9290 3957 9324
rect 3992 9290 4026 9324
rect 4061 9290 4095 9324
rect 4130 9290 4164 9324
rect 4199 9290 4233 9324
rect 4268 9290 4302 9324
rect 4337 9290 4371 9324
rect 4406 9290 4440 9324
rect 4475 9290 4509 9324
rect 4544 9290 4578 9324
rect 4613 9290 4647 9324
rect 4682 9290 4716 9324
rect 4751 9290 4785 9324
rect 4820 9290 4854 9324
rect 4889 9290 4923 9324
rect 4958 9290 4992 9324
rect 5027 9290 5061 9324
rect 5096 9290 5130 9324
rect 5165 9290 5199 9324
rect 5234 9290 5268 9324
rect 5303 9290 5337 9324
rect 5372 9290 5406 9324
rect 5441 9290 5475 9324
rect 5510 9290 5544 9324
rect 5579 9290 5613 9324
rect 5648 9290 5682 9324
rect 5717 9290 5751 9324
rect 5786 9290 5820 9324
rect 5855 9290 5889 9324
rect 5924 9290 5958 9324
rect 5993 9290 6027 9324
rect 6062 9290 6096 9324
rect 6131 9290 6165 9324
rect 6200 9290 6234 9324
rect 6268 9290 6302 9324
rect 6336 9290 6370 9324
rect 6404 9290 6438 9324
rect 6472 9290 6506 9324
rect 6540 9290 6574 9324
rect 6608 9290 6642 9324
rect 6676 9290 6710 9324
rect 6744 9290 6778 9324
rect 6812 9290 6846 9324
rect 6880 9290 6914 9324
rect 6948 9290 6982 9324
rect 7016 9290 7050 9324
rect 7084 9290 7118 9324
rect 7152 9290 7186 9324
rect 7220 9290 7254 9324
rect 7288 9290 7322 9324
rect 7356 9290 7390 9324
rect 7424 9290 7458 9324
rect 7492 9290 7526 9324
rect 7560 9290 7594 9324
rect 7628 9290 7662 9324
rect 7696 9290 7730 9324
rect 7764 9290 7798 9324
rect 7832 9290 7866 9324
rect 7900 9290 7934 9324
rect 7968 9290 8002 9324
rect 8036 9290 8070 9324
rect 8104 9290 8138 9324
rect 8172 9290 8206 9324
rect 8240 9290 8274 9324
rect 8308 9290 8342 9324
rect 8376 9290 8410 9324
rect 8444 9290 8478 9324
rect 8512 9290 8546 9324
rect 8580 9290 8614 9324
rect 8648 9290 8682 9324
rect 8716 9290 8750 9324
rect 8784 9290 8818 9324
rect 8852 9290 8886 9324
rect 8920 9290 8954 9324
rect 8988 9290 9022 9324
rect 9056 9290 9090 9324
rect 9124 9290 9158 9324
rect 9192 9290 9226 9324
rect 9260 9290 9294 9324
rect 9328 9290 9362 9324
rect 9396 9290 9430 9324
rect 9464 9290 9498 9324
rect 9532 9290 9566 9324
rect 9600 9290 9634 9324
rect 9668 9290 9702 9324
rect 9736 9290 9770 9324
rect 9804 9290 9838 9324
rect 9872 9290 9906 9324
rect 9940 9290 9974 9324
rect 10008 9290 10042 9324
rect 10076 9290 10110 9324
rect 10144 9290 10178 9324
rect 10212 9290 10246 9324
rect 10280 9290 10314 9324
rect 10348 9290 10382 9324
rect 10416 9290 10450 9324
rect 10484 9290 10518 9324
rect 10552 9290 10586 9324
rect 10620 9290 10654 9324
rect 10688 9290 10722 9324
rect 10756 9290 10790 9324
rect 10824 9290 10858 9324
rect 10892 9290 10926 9324
rect 10960 9290 10994 9324
rect 11028 9290 11062 9324
rect 11096 9290 11130 9324
rect 11164 9290 11198 9324
rect 11232 9290 11266 9324
rect 11300 9290 11334 9324
rect 11368 9290 11402 9324
rect 11436 9290 11470 9324
rect 11504 9290 11538 9324
rect 11572 9290 11606 9324
rect 11640 9290 11674 9324
rect 11708 9290 11742 9324
rect 11776 9290 11810 9324
rect 11844 9290 11878 9324
rect 11912 9290 11946 9324
rect 11980 9290 12014 9324
rect 12048 9290 12082 9324
rect 12116 9290 12150 9324
rect 12184 9290 12218 9324
rect 12252 9290 12286 9324
rect 12320 9290 12354 9324
rect 12388 9290 12422 9324
rect 12456 9290 12490 9324
rect 12524 9290 12558 9324
rect 12592 9290 12626 9324
rect 12660 9290 12694 9324
rect 12728 9290 12762 9324
rect 12796 9290 12830 9324
rect 12864 9290 12898 9324
rect 12932 9290 12966 9324
rect 13000 9290 13034 9324
rect 13068 9290 13102 9324
rect 2888 8820 2922 8854
rect 2957 8820 2991 8854
rect 3026 8820 3060 8854
rect 3095 8820 3129 8854
rect 3164 8820 3198 8854
rect 3233 8820 3267 8854
rect 3302 8820 3336 8854
rect 3371 8820 3405 8854
rect 3440 8820 3474 8854
rect 3509 8820 3543 8854
rect 3578 8820 3612 8854
rect 3647 8820 3681 8854
rect 3716 8820 3750 8854
rect 3785 8820 3819 8854
rect 3854 8820 3888 8854
rect 3923 8820 3957 8854
rect 3992 8820 4026 8854
rect 4061 8820 4095 8854
rect 4130 8820 4164 8854
rect 4199 8820 4233 8854
rect 4268 8820 4302 8854
rect 4337 8820 4371 8854
rect 4406 8820 4440 8854
rect 4475 8820 4509 8854
rect 4544 8820 4578 8854
rect 4613 8820 4647 8854
rect 4682 8820 4716 8854
rect 4751 8820 4785 8854
rect 4820 8820 4854 8854
rect 4889 8820 4923 8854
rect 4958 8820 4992 8854
rect 5027 8820 5061 8854
rect 5096 8820 5130 8854
rect 5165 8820 5199 8854
rect 5234 8820 5268 8854
rect 5303 8820 5337 8854
rect 5372 8820 5406 8854
rect 5441 8820 5475 8854
rect 5510 8820 5544 8854
rect 5579 8820 5613 8854
rect 5648 8820 5682 8854
rect 5717 8820 5751 8854
rect 5786 8820 5820 8854
rect 5855 8820 5889 8854
rect 5924 8820 5958 8854
rect 5993 8820 6027 8854
rect 6062 8820 6096 8854
rect 6131 8820 6165 8854
rect 6200 8820 6234 8854
rect 6268 8820 6302 8854
rect 6336 8820 6370 8854
rect 6404 8820 6438 8854
rect 6472 8820 6506 8854
rect 6540 8820 6574 8854
rect 6608 8820 6642 8854
rect 6676 8820 6710 8854
rect 6744 8820 6778 8854
rect 6812 8820 6846 8854
rect 6880 8820 6914 8854
rect 6948 8820 6982 8854
rect 7016 8820 7050 8854
rect 7084 8820 7118 8854
rect 7152 8820 7186 8854
rect 7220 8820 7254 8854
rect 7288 8820 7322 8854
rect 7356 8820 7390 8854
rect 7424 8820 7458 8854
rect 7492 8820 7526 8854
rect 7560 8820 7594 8854
rect 7628 8820 7662 8854
rect 7696 8820 7730 8854
rect 7764 8820 7798 8854
rect 7832 8820 7866 8854
rect 7900 8820 7934 8854
rect 7968 8820 8002 8854
rect 8036 8820 8070 8854
rect 8104 8820 8138 8854
rect 8172 8820 8206 8854
rect 8240 8820 8274 8854
rect 8308 8820 8342 8854
rect 8376 8820 8410 8854
rect 8444 8820 8478 8854
rect 8512 8820 8546 8854
rect 8580 8820 8614 8854
rect 8648 8820 8682 8854
rect 8716 8820 8750 8854
rect 8784 8820 8818 8854
rect 8852 8820 8886 8854
rect 8920 8820 8954 8854
rect 8988 8820 9022 8854
rect 9056 8820 9090 8854
rect 9124 8820 9158 8854
rect 9192 8820 9226 8854
rect 9260 8820 9294 8854
rect 9328 8820 9362 8854
rect 9396 8820 9430 8854
rect 9464 8820 9498 8854
rect 9532 8820 9566 8854
rect 9600 8820 9634 8854
rect 9668 8820 9702 8854
rect 9736 8820 9770 8854
rect 9804 8820 9838 8854
rect 9872 8820 9906 8854
rect 9940 8820 9974 8854
rect 10008 8820 10042 8854
rect 10076 8820 10110 8854
rect 10144 8820 10178 8854
rect 10212 8820 10246 8854
rect 10280 8820 10314 8854
rect 10348 8820 10382 8854
rect 10416 8820 10450 8854
rect 10484 8820 10518 8854
rect 10552 8820 10586 8854
rect 10620 8820 10654 8854
rect 10688 8820 10722 8854
rect 10756 8820 10790 8854
rect 10824 8820 10858 8854
rect 10892 8820 10926 8854
rect 10960 8820 10994 8854
rect 11028 8820 11062 8854
rect 11096 8820 11130 8854
rect 11164 8820 11198 8854
rect 11232 8820 11266 8854
rect 11300 8820 11334 8854
rect 11368 8820 11402 8854
rect 11436 8820 11470 8854
rect 11504 8820 11538 8854
rect 11572 8820 11606 8854
rect 11640 8820 11674 8854
rect 11708 8820 11742 8854
rect 11776 8820 11810 8854
rect 11844 8820 11878 8854
rect 11912 8820 11946 8854
rect 11980 8820 12014 8854
rect 12048 8820 12082 8854
rect 12116 8820 12150 8854
rect 12184 8820 12218 8854
rect 12252 8820 12286 8854
rect 12320 8820 12354 8854
rect 12388 8820 12422 8854
rect 12456 8820 12490 8854
rect 12524 8820 12558 8854
rect 12592 8820 12626 8854
rect 12660 8820 12694 8854
rect 12728 8820 12762 8854
rect 12796 8820 12830 8854
rect 12864 8820 12898 8854
rect 12932 8820 12966 8854
rect 13000 8820 13034 8854
rect 13068 8820 13102 8854
rect 2888 7290 2922 7324
rect 2957 7290 2991 7324
rect 3026 7290 3060 7324
rect 3095 7290 3129 7324
rect 3164 7290 3198 7324
rect 3233 7290 3267 7324
rect 3302 7290 3336 7324
rect 3371 7290 3405 7324
rect 3440 7290 3474 7324
rect 3509 7290 3543 7324
rect 3578 7290 3612 7324
rect 3647 7290 3681 7324
rect 3716 7290 3750 7324
rect 3785 7290 3819 7324
rect 3854 7290 3888 7324
rect 3923 7290 3957 7324
rect 3992 7290 4026 7324
rect 4061 7290 4095 7324
rect 4130 7290 4164 7324
rect 4199 7290 4233 7324
rect 4268 7290 4302 7324
rect 4337 7290 4371 7324
rect 4406 7290 4440 7324
rect 4475 7290 4509 7324
rect 4544 7290 4578 7324
rect 4613 7290 4647 7324
rect 4682 7290 4716 7324
rect 4751 7290 4785 7324
rect 4820 7290 4854 7324
rect 4889 7290 4923 7324
rect 4958 7290 4992 7324
rect 5027 7290 5061 7324
rect 5096 7290 5130 7324
rect 5165 7290 5199 7324
rect 5234 7290 5268 7324
rect 5303 7290 5337 7324
rect 5372 7290 5406 7324
rect 5441 7290 5475 7324
rect 5510 7290 5544 7324
rect 5579 7290 5613 7324
rect 5648 7290 5682 7324
rect 5717 7290 5751 7324
rect 5786 7290 5820 7324
rect 5855 7290 5889 7324
rect 5924 7290 5958 7324
rect 5993 7290 6027 7324
rect 6062 7290 6096 7324
rect 6131 7290 6165 7324
rect 6200 7290 6234 7324
rect 6268 7290 6302 7324
rect 6336 7290 6370 7324
rect 6404 7290 6438 7324
rect 6472 7290 6506 7324
rect 6540 7290 6574 7324
rect 6608 7290 6642 7324
rect 6676 7290 6710 7324
rect 6744 7290 6778 7324
rect 6812 7290 6846 7324
rect 6880 7290 6914 7324
rect 6948 7290 6982 7324
rect 7016 7290 7050 7324
rect 7084 7290 7118 7324
rect 7152 7290 7186 7324
rect 7220 7290 7254 7324
rect 7288 7290 7322 7324
rect 7356 7290 7390 7324
rect 7424 7290 7458 7324
rect 7492 7290 7526 7324
rect 7560 7290 7594 7324
rect 7628 7290 7662 7324
rect 7696 7290 7730 7324
rect 7764 7290 7798 7324
rect 7832 7290 7866 7324
rect 7900 7290 7934 7324
rect 7968 7290 8002 7324
rect 8036 7290 8070 7324
rect 8104 7290 8138 7324
rect 8172 7290 8206 7324
rect 8240 7290 8274 7324
rect 8308 7290 8342 7324
rect 8376 7290 8410 7324
rect 8444 7290 8478 7324
rect 8512 7290 8546 7324
rect 8580 7290 8614 7324
rect 8648 7290 8682 7324
rect 8716 7290 8750 7324
rect 8784 7290 8818 7324
rect 8852 7290 8886 7324
rect 8920 7290 8954 7324
rect 8988 7290 9022 7324
rect 9056 7290 9090 7324
rect 9124 7290 9158 7324
rect 9192 7290 9226 7324
rect 9260 7290 9294 7324
rect 9328 7290 9362 7324
rect 9396 7290 9430 7324
rect 9464 7290 9498 7324
rect 9532 7290 9566 7324
rect 9600 7290 9634 7324
rect 9668 7290 9702 7324
rect 9736 7290 9770 7324
rect 9804 7290 9838 7324
rect 9872 7290 9906 7324
rect 9940 7290 9974 7324
rect 10008 7290 10042 7324
rect 10076 7290 10110 7324
rect 10144 7290 10178 7324
rect 10212 7290 10246 7324
rect 10280 7290 10314 7324
rect 10348 7290 10382 7324
rect 10416 7290 10450 7324
rect 10484 7290 10518 7324
rect 10552 7290 10586 7324
rect 10620 7290 10654 7324
rect 10688 7290 10722 7324
rect 10756 7290 10790 7324
rect 10824 7290 10858 7324
rect 10892 7290 10926 7324
rect 10960 7290 10994 7324
rect 11028 7290 11062 7324
rect 11096 7290 11130 7324
rect 11164 7290 11198 7324
rect 11232 7290 11266 7324
rect 11300 7290 11334 7324
rect 11368 7290 11402 7324
rect 11436 7290 11470 7324
rect 11504 7290 11538 7324
rect 11572 7290 11606 7324
rect 11640 7290 11674 7324
rect 11708 7290 11742 7324
rect 11776 7290 11810 7324
rect 11844 7290 11878 7324
rect 11912 7290 11946 7324
rect 11980 7290 12014 7324
rect 12048 7290 12082 7324
rect 12116 7290 12150 7324
rect 12184 7290 12218 7324
rect 12252 7290 12286 7324
rect 12320 7290 12354 7324
rect 12388 7290 12422 7324
rect 12456 7290 12490 7324
rect 12524 7290 12558 7324
rect 12592 7290 12626 7324
rect 12660 7290 12694 7324
rect 12728 7290 12762 7324
rect 12796 7290 12830 7324
rect 12864 7290 12898 7324
rect 12932 7290 12966 7324
rect 13000 7290 13034 7324
rect 13068 7290 13102 7324
rect 2888 6820 2922 6854
rect 2957 6820 2991 6854
rect 3026 6820 3060 6854
rect 3095 6820 3129 6854
rect 3164 6820 3198 6854
rect 3233 6820 3267 6854
rect 3302 6820 3336 6854
rect 3371 6820 3405 6854
rect 3440 6820 3474 6854
rect 3509 6820 3543 6854
rect 3578 6820 3612 6854
rect 3647 6820 3681 6854
rect 3716 6820 3750 6854
rect 3785 6820 3819 6854
rect 3854 6820 3888 6854
rect 3923 6820 3957 6854
rect 3992 6820 4026 6854
rect 4061 6820 4095 6854
rect 4130 6820 4164 6854
rect 4199 6820 4233 6854
rect 4268 6820 4302 6854
rect 4337 6820 4371 6854
rect 4406 6820 4440 6854
rect 4475 6820 4509 6854
rect 4544 6820 4578 6854
rect 4613 6820 4647 6854
rect 4682 6820 4716 6854
rect 4751 6820 4785 6854
rect 4820 6820 4854 6854
rect 4889 6820 4923 6854
rect 4958 6820 4992 6854
rect 5027 6820 5061 6854
rect 5096 6820 5130 6854
rect 5165 6820 5199 6854
rect 5234 6820 5268 6854
rect 5303 6820 5337 6854
rect 5372 6820 5406 6854
rect 5441 6820 5475 6854
rect 5510 6820 5544 6854
rect 5579 6820 5613 6854
rect 5648 6820 5682 6854
rect 5717 6820 5751 6854
rect 5786 6820 5820 6854
rect 5855 6820 5889 6854
rect 5924 6820 5958 6854
rect 5993 6820 6027 6854
rect 6062 6820 6096 6854
rect 6131 6820 6165 6854
rect 6200 6820 6234 6854
rect 6268 6820 6302 6854
rect 6336 6820 6370 6854
rect 6404 6820 6438 6854
rect 6472 6820 6506 6854
rect 6540 6820 6574 6854
rect 6608 6820 6642 6854
rect 6676 6820 6710 6854
rect 6744 6820 6778 6854
rect 6812 6820 6846 6854
rect 6880 6820 6914 6854
rect 6948 6820 6982 6854
rect 7016 6820 7050 6854
rect 7084 6820 7118 6854
rect 7152 6820 7186 6854
rect 7220 6820 7254 6854
rect 7288 6820 7322 6854
rect 7356 6820 7390 6854
rect 7424 6820 7458 6854
rect 7492 6820 7526 6854
rect 7560 6820 7594 6854
rect 7628 6820 7662 6854
rect 7696 6820 7730 6854
rect 7764 6820 7798 6854
rect 7832 6820 7866 6854
rect 7900 6820 7934 6854
rect 7968 6820 8002 6854
rect 8036 6820 8070 6854
rect 8104 6820 8138 6854
rect 8172 6820 8206 6854
rect 8240 6820 8274 6854
rect 8308 6820 8342 6854
rect 8376 6820 8410 6854
rect 8444 6820 8478 6854
rect 8512 6820 8546 6854
rect 8580 6820 8614 6854
rect 8648 6820 8682 6854
rect 8716 6820 8750 6854
rect 8784 6820 8818 6854
rect 8852 6820 8886 6854
rect 8920 6820 8954 6854
rect 8988 6820 9022 6854
rect 9056 6820 9090 6854
rect 9124 6820 9158 6854
rect 9192 6820 9226 6854
rect 9260 6820 9294 6854
rect 9328 6820 9362 6854
rect 9396 6820 9430 6854
rect 9464 6820 9498 6854
rect 9532 6820 9566 6854
rect 9600 6820 9634 6854
rect 9668 6820 9702 6854
rect 9736 6820 9770 6854
rect 9804 6820 9838 6854
rect 9872 6820 9906 6854
rect 9940 6820 9974 6854
rect 10008 6820 10042 6854
rect 10076 6820 10110 6854
rect 10144 6820 10178 6854
rect 10212 6820 10246 6854
rect 10280 6820 10314 6854
rect 10348 6820 10382 6854
rect 10416 6820 10450 6854
rect 10484 6820 10518 6854
rect 10552 6820 10586 6854
rect 10620 6820 10654 6854
rect 10688 6820 10722 6854
rect 10756 6820 10790 6854
rect 10824 6820 10858 6854
rect 10892 6820 10926 6854
rect 10960 6820 10994 6854
rect 11028 6820 11062 6854
rect 11096 6820 11130 6854
rect 11164 6820 11198 6854
rect 11232 6820 11266 6854
rect 11300 6820 11334 6854
rect 11368 6820 11402 6854
rect 11436 6820 11470 6854
rect 11504 6820 11538 6854
rect 11572 6820 11606 6854
rect 11640 6820 11674 6854
rect 11708 6820 11742 6854
rect 11776 6820 11810 6854
rect 11844 6820 11878 6854
rect 11912 6820 11946 6854
rect 11980 6820 12014 6854
rect 12048 6820 12082 6854
rect 12116 6820 12150 6854
rect 12184 6820 12218 6854
rect 12252 6820 12286 6854
rect 12320 6820 12354 6854
rect 12388 6820 12422 6854
rect 12456 6820 12490 6854
rect 12524 6820 12558 6854
rect 12592 6820 12626 6854
rect 12660 6820 12694 6854
rect 12728 6820 12762 6854
rect 12796 6820 12830 6854
rect 12864 6820 12898 6854
rect 12932 6820 12966 6854
rect 13000 6820 13034 6854
rect 13068 6820 13102 6854
rect 1887 4500 1921 4534
rect 1955 4500 1989 4534
rect 64 3806 98 3840
rect 64 3738 98 3772
rect 430 1852 464 1886
rect 503 1852 537 1886
rect 576 1852 610 1886
rect 649 1852 683 1886
rect 722 1852 756 1886
rect 795 1852 829 1886
rect 868 1852 902 1886
rect 940 1852 974 1886
rect 1012 1852 1046 1886
rect 1084 1852 1118 1886
rect 1156 1852 1190 1886
rect 1228 1852 1262 1886
rect 430 322 464 356
rect 503 322 537 356
rect 576 322 610 356
rect 649 322 683 356
rect 722 322 756 356
rect 795 322 829 356
rect 868 322 902 356
rect 940 322 974 356
rect 1012 322 1046 356
rect 1084 322 1118 356
rect 1156 322 1190 356
rect 1228 322 1262 356
rect 13683 1864 13717 1898
rect 13756 1864 13790 1898
rect 13829 1864 13863 1898
rect 13902 1864 13936 1898
rect 13975 1864 14009 1898
rect 14048 1864 14082 1898
rect 14121 1864 14155 1898
rect 14193 1864 14227 1898
rect 14265 1864 14299 1898
rect 14337 1864 14371 1898
rect 14409 1864 14443 1898
rect 14481 1864 14515 1898
rect 13683 334 13717 368
rect 13756 334 13790 368
rect 13829 334 13863 368
rect 13902 334 13936 368
rect 13975 334 14009 368
rect 14048 334 14082 368
rect 14121 334 14155 368
rect 14193 334 14227 368
rect 14265 334 14299 368
rect 14337 334 14371 368
rect 14409 334 14443 368
rect 14481 334 14515 368
<< locali >>
rect 14809 39522 14917 39556
rect 1831 39474 2163 39476
rect 10189 39474 10228 39476
rect 10262 39474 10301 39476
rect 10335 39474 10374 39476
rect 10408 39474 10447 39476
rect 10481 39474 10520 39476
rect 10554 39474 10593 39476
rect 10627 39474 10666 39476
rect 10700 39474 10739 39476
rect 10773 39474 10812 39476
rect 10846 39474 10885 39476
rect 10919 39474 10958 39476
rect 10992 39474 11031 39476
rect 11065 39474 11104 39476
rect 11138 39474 11177 39476
rect 11211 39474 11250 39476
rect 11284 39474 11323 39476
rect 11357 39474 11396 39476
rect 11430 39474 11469 39476
rect 11503 39474 11542 39476
rect 11576 39474 11615 39476
rect 11649 39474 11688 39476
rect 11722 39474 11761 39476
rect 11795 39474 11834 39476
rect 11868 39474 11907 39476
rect 11941 39474 11980 39476
rect 12014 39474 12053 39476
rect 12087 39474 12126 39476
rect 12160 39474 12199 39476
rect 12233 39474 12272 39476
rect 12306 39474 12345 39476
rect 12379 39474 12418 39476
rect 12452 39474 12491 39476
rect 12525 39474 12564 39476
rect 12598 39474 12637 39476
rect 12671 39474 12710 39476
rect 12744 39474 12783 39476
rect 12817 39474 12856 39476
rect 12890 39474 12929 39476
rect 12963 39474 13002 39476
rect 13036 39474 13075 39476
rect 13109 39474 13148 39476
rect 13182 39474 13221 39476
rect 13255 39474 13294 39476
rect 13328 39474 13367 39476
rect 13401 39474 13440 39476
rect 13474 39474 13513 39476
rect 13547 39474 13586 39476
rect 13620 39474 13659 39476
rect 13693 39474 13732 39476
rect 13766 39474 13944 39476
rect 1831 39470 2076 39474
rect 1668 39238 1684 39284
rect 1718 39238 1734 39284
rect 1668 39212 1734 39238
rect 1668 39170 1684 39212
rect 1718 39170 1734 39212
rect 1831 34108 1944 39470
rect 2050 39440 2076 39470
rect 2110 39440 2144 39474
rect 2050 39372 2144 39440
rect 13874 39470 13944 39474
rect 14775 39418 14951 39522
rect 14809 39384 14917 39418
rect 2050 39370 2163 39372
rect 10189 39370 10228 39372
rect 10262 39370 10301 39372
rect 10335 39370 10374 39372
rect 10408 39370 10447 39372
rect 10481 39370 10520 39372
rect 10554 39370 10593 39372
rect 10627 39370 10666 39372
rect 10700 39370 10739 39372
rect 10773 39370 10812 39372
rect 10846 39370 10885 39372
rect 10919 39370 10958 39372
rect 10992 39370 11031 39372
rect 11065 39370 11104 39372
rect 11138 39370 11177 39372
rect 11211 39370 11250 39372
rect 11284 39370 11323 39372
rect 11357 39370 11396 39372
rect 11430 39370 11469 39372
rect 11503 39370 11542 39372
rect 11576 39370 11615 39372
rect 11649 39370 11688 39372
rect 11722 39370 11761 39372
rect 11795 39370 11834 39372
rect 11868 39370 11907 39372
rect 11941 39370 11980 39372
rect 12014 39370 12053 39372
rect 12087 39370 12126 39372
rect 12160 39370 12199 39372
rect 12233 39370 12272 39372
rect 12306 39370 12345 39372
rect 12379 39370 12418 39372
rect 12452 39370 12491 39372
rect 12525 39370 12564 39372
rect 12598 39370 12637 39372
rect 12671 39370 12710 39372
rect 12744 39370 12783 39372
rect 12817 39370 12856 39372
rect 12890 39370 12929 39372
rect 12963 39370 13002 39372
rect 13036 39370 13075 39372
rect 13109 39370 13148 39372
rect 13182 39370 13221 39372
rect 13255 39370 13294 39372
rect 13328 39370 13367 39372
rect 13401 39370 13440 39372
rect 13474 39370 13513 39372
rect 13547 39370 13586 39372
rect 13620 39370 13659 39372
rect 13693 39370 13732 39372
rect 13766 39370 13838 39372
rect 2050 34108 2056 39370
rect 1831 34069 1946 34108
rect 2048 34069 2056 34108
rect 1831 34035 1944 34069
rect 2050 34035 2056 34069
rect 1831 33996 1946 34035
rect 2048 33996 2056 34035
rect 1831 33962 1944 33996
rect 2050 33962 2056 33996
rect 1831 33923 1946 33962
rect 2048 33923 2056 33962
rect 1831 33889 1944 33923
rect 2050 33889 2056 33923
rect 1831 33850 1946 33889
rect 2048 33850 2056 33889
rect 1831 33816 1944 33850
rect 2050 33816 2056 33850
rect 1831 33777 1946 33816
rect 2048 33777 2056 33816
rect 1831 33743 1944 33777
rect 2050 33743 2056 33777
rect 1831 33704 1946 33743
rect 2048 33704 2056 33743
rect 1831 33670 1944 33704
rect 2050 33670 2056 33704
rect 1831 21393 1946 33670
rect 1871 19864 1909 19898
rect 1943 19864 1946 19898
rect 1837 19821 1946 19864
rect 1871 19787 1909 19821
rect 1943 19787 1946 19821
rect 1837 19744 1946 19787
rect 1871 19710 1909 19744
rect 1943 19710 1946 19744
rect 1837 19667 1946 19710
rect 1871 19633 1909 19667
rect 1943 19633 1946 19667
rect 1837 19477 1946 19633
rect 2048 19477 2056 33670
rect 2213 39171 13699 39177
rect 2213 39119 2291 39171
rect 9957 39153 9996 39171
rect 10030 39153 10069 39171
rect 10103 39153 10142 39171
rect 10176 39153 10215 39171
rect 10249 39153 10288 39171
rect 9957 39119 9978 39153
rect 10030 39137 10047 39153
rect 10103 39137 10116 39153
rect 10176 39137 10185 39153
rect 10249 39137 10254 39153
rect 10012 39119 10047 39137
rect 10081 39119 10116 39137
rect 10150 39119 10185 39137
rect 10219 39119 10254 39137
rect 10322 39153 10361 39171
rect 10395 39153 10434 39171
rect 10468 39153 10507 39171
rect 10541 39153 10580 39171
rect 10614 39153 10653 39171
rect 10687 39153 10726 39171
rect 10760 39153 10799 39171
rect 10833 39153 10872 39171
rect 10906 39153 10945 39171
rect 10979 39153 11018 39171
rect 11052 39153 11091 39171
rect 11125 39153 11164 39171
rect 11198 39153 11237 39171
rect 11271 39153 11310 39171
rect 11344 39153 11383 39171
rect 11417 39153 11456 39171
rect 11490 39153 11529 39171
rect 11563 39153 11602 39171
rect 11636 39153 11675 39171
rect 11709 39153 11748 39171
rect 11782 39153 11821 39171
rect 11855 39153 11894 39171
rect 11928 39153 11967 39171
rect 12001 39153 12040 39171
rect 12074 39153 12113 39171
rect 12147 39153 12186 39171
rect 12220 39153 12259 39171
rect 12293 39153 12332 39171
rect 12366 39153 12405 39171
rect 12439 39153 12478 39171
rect 12512 39153 12551 39171
rect 12585 39153 12624 39171
rect 12658 39153 12697 39171
rect 12731 39153 12770 39171
rect 12804 39153 12843 39171
rect 12877 39153 12916 39171
rect 12950 39153 12989 39171
rect 13095 39153 13137 39171
rect 13171 39153 13213 39171
rect 13247 39153 13289 39171
rect 13323 39153 13365 39171
rect 13399 39153 13441 39171
rect 10322 39137 10323 39153
rect 10288 39119 10323 39137
rect 10357 39137 10361 39153
rect 10426 39137 10434 39153
rect 10495 39137 10507 39153
rect 10564 39137 10580 39153
rect 10633 39137 10653 39153
rect 10702 39137 10726 39153
rect 10771 39137 10799 39153
rect 10840 39137 10872 39153
rect 10357 39119 10392 39137
rect 10426 39119 10461 39137
rect 10495 39119 10530 39137
rect 10564 39119 10599 39137
rect 10633 39119 10668 39137
rect 10702 39119 10737 39137
rect 10771 39119 10806 39137
rect 10840 39119 10875 39137
rect 10909 39119 10944 39153
rect 10979 39137 11013 39153
rect 11052 39137 11082 39153
rect 11125 39137 11151 39153
rect 11198 39137 11220 39153
rect 11271 39137 11289 39153
rect 11344 39137 11358 39153
rect 11417 39137 11427 39153
rect 11490 39137 11496 39153
rect 11563 39137 11565 39153
rect 10978 39119 11013 39137
rect 11047 39119 11082 39137
rect 11116 39119 11151 39137
rect 11185 39119 11220 39137
rect 11254 39119 11289 39137
rect 11323 39119 11358 39137
rect 11392 39119 11427 39137
rect 11461 39119 11496 39137
rect 11530 39119 11565 39137
rect 11599 39137 11602 39153
rect 11668 39137 11675 39153
rect 11737 39137 11748 39153
rect 11806 39137 11821 39153
rect 11875 39137 11894 39153
rect 11944 39137 11967 39153
rect 12013 39137 12040 39153
rect 12082 39137 12113 39153
rect 11599 39119 11634 39137
rect 11668 39119 11703 39137
rect 11737 39119 11772 39137
rect 11806 39119 11841 39137
rect 11875 39119 11910 39137
rect 11944 39119 11979 39137
rect 12013 39119 12048 39137
rect 12082 39119 12117 39137
rect 12151 39119 12186 39153
rect 12220 39119 12255 39153
rect 12293 39137 12324 39153
rect 12366 39137 12393 39153
rect 12439 39137 12462 39153
rect 12512 39137 12531 39153
rect 12585 39137 12600 39153
rect 12658 39137 12669 39153
rect 12731 39137 12738 39153
rect 12804 39137 12807 39153
rect 12289 39119 12324 39137
rect 12358 39119 12393 39137
rect 12427 39119 12462 39137
rect 12496 39119 12531 39137
rect 12565 39119 12600 39137
rect 12634 39119 12669 39137
rect 12703 39119 12738 39137
rect 12772 39119 12807 39137
rect 12841 39137 12843 39153
rect 12910 39137 12916 39153
rect 12841 39119 12876 39137
rect 12910 39119 12945 39137
rect 12979 39119 12989 39153
rect 13117 39137 13137 39153
rect 13186 39137 13213 39153
rect 13255 39137 13289 39153
rect 13117 39119 13152 39137
rect 13186 39119 13221 39137
rect 13255 39119 13290 39137
rect 13324 39119 13359 39153
rect 13399 39137 13428 39153
rect 13475 39137 13517 39171
rect 13551 39137 13593 39171
rect 13627 39137 13699 39171
rect 13393 39119 13428 39137
rect 13462 39129 13699 39137
rect 13462 39119 13515 39129
rect 2213 39099 2274 39119
rect 2213 39065 2219 39099
rect 2253 39065 2274 39099
rect 2213 39026 2274 39065
rect 2213 38992 2219 39026
rect 2253 38992 2274 39026
rect 9957 39099 12989 39119
rect 9957 39065 9996 39099
rect 10030 39065 10069 39099
rect 10103 39065 10142 39099
rect 10176 39065 10215 39099
rect 10249 39065 10288 39099
rect 10322 39065 10361 39099
rect 10395 39065 10434 39099
rect 10468 39065 10507 39099
rect 10541 39065 10580 39099
rect 10614 39065 10653 39099
rect 10687 39065 10726 39099
rect 10760 39065 10799 39099
rect 10833 39065 10872 39099
rect 10906 39065 10945 39099
rect 10979 39065 11018 39099
rect 11052 39065 11091 39099
rect 11125 39065 11164 39099
rect 11198 39065 11237 39099
rect 11271 39065 11310 39099
rect 11344 39065 11383 39099
rect 11417 39065 11456 39099
rect 11490 39065 11529 39099
rect 11563 39065 11602 39099
rect 11636 39065 11675 39099
rect 11709 39065 11748 39099
rect 11782 39065 11821 39099
rect 11855 39065 11894 39099
rect 11928 39065 11967 39099
rect 12001 39065 12040 39099
rect 12074 39065 12113 39099
rect 12147 39065 12186 39099
rect 12220 39065 12259 39099
rect 12293 39065 12332 39099
rect 12366 39065 12405 39099
rect 12439 39065 12478 39099
rect 12512 39065 12551 39099
rect 12585 39065 12624 39099
rect 12658 39065 12697 39099
rect 12731 39065 12770 39099
rect 12804 39065 12843 39099
rect 12877 39065 12916 39099
rect 12950 39065 12989 39099
rect 9957 39027 12989 39065
rect 13095 39099 13515 39119
rect 13617 39099 13699 39129
rect 13095 39065 13137 39099
rect 13171 39065 13213 39099
rect 13247 39065 13289 39099
rect 13323 39065 13365 39099
rect 13399 39065 13441 39099
rect 13475 39065 13515 39099
rect 13095 39027 13515 39065
rect 9957 38993 9978 39027
rect 10030 38993 10047 39027
rect 10103 38993 10116 39027
rect 10176 38993 10185 39027
rect 10249 38993 10254 39027
rect 10322 38993 10323 39027
rect 10357 38993 10361 39027
rect 10426 38993 10434 39027
rect 10495 38993 10507 39027
rect 10564 38993 10580 39027
rect 10633 38993 10653 39027
rect 10702 38993 10726 39027
rect 10771 38993 10799 39027
rect 10840 38993 10872 39027
rect 10909 38993 10944 39027
rect 10979 38993 11013 39027
rect 11052 38993 11082 39027
rect 11125 38993 11151 39027
rect 11198 38993 11220 39027
rect 11271 38993 11289 39027
rect 11344 38993 11358 39027
rect 11417 38993 11427 39027
rect 11490 38993 11496 39027
rect 11563 38993 11565 39027
rect 11599 38993 11602 39027
rect 11668 38993 11675 39027
rect 11737 38993 11748 39027
rect 11806 38993 11821 39027
rect 11875 38993 11894 39027
rect 11944 38993 11967 39027
rect 12013 38993 12040 39027
rect 12082 38993 12113 39027
rect 12151 38993 12186 39027
rect 12220 38993 12255 39027
rect 12293 38993 12324 39027
rect 12366 38993 12393 39027
rect 12439 38993 12462 39027
rect 12512 38993 12531 39027
rect 12585 38993 12600 39027
rect 12658 38993 12669 39027
rect 12731 38993 12738 39027
rect 12804 38993 12807 39027
rect 12841 38993 12843 39027
rect 12910 38993 12916 39027
rect 12979 38993 12989 39027
rect 13117 38993 13137 39027
rect 13186 38993 13213 39027
rect 13255 38993 13290 39027
rect 13324 38993 13359 39027
rect 13401 38993 13428 39027
rect 13478 38993 13515 39027
rect 2213 38953 2274 38992
rect 2444 38987 13515 38993
rect 2213 38919 2219 38953
rect 2253 38919 2274 38953
rect 2213 38880 2274 38919
rect 2213 38846 2219 38880
rect 2253 38846 2274 38880
rect 2213 38807 2274 38846
rect 2872 38820 2884 38854
rect 2922 38820 2957 38854
rect 2991 38820 3026 38854
rect 3064 38820 3095 38854
rect 3137 38820 3164 38854
rect 3210 38820 3233 38854
rect 3283 38820 3302 38854
rect 3356 38820 3371 38854
rect 3429 38820 3440 38854
rect 3502 38820 3509 38854
rect 3575 38820 3578 38854
rect 3612 38820 3614 38854
rect 3681 38820 3687 38854
rect 3750 38820 3760 38854
rect 3819 38820 3833 38854
rect 3888 38820 3906 38854
rect 3957 38820 3979 38854
rect 4026 38820 4052 38854
rect 4095 38820 4125 38854
rect 4164 38820 4198 38854
rect 4233 38820 4268 38854
rect 4305 38820 4337 38854
rect 4378 38820 4406 38854
rect 4451 38820 4475 38854
rect 4524 38820 4544 38854
rect 4597 38820 4613 38854
rect 4670 38820 4682 38854
rect 4743 38820 4751 38854
rect 4816 38820 4820 38854
rect 4854 38820 4855 38854
rect 4923 38820 4928 38854
rect 4992 38820 5001 38854
rect 5061 38820 5074 38854
rect 5130 38820 5147 38854
rect 5199 38820 5220 38854
rect 5268 38820 5293 38854
rect 5337 38820 5366 38854
rect 5406 38820 5439 38854
rect 5475 38820 5510 38854
rect 5546 38820 5579 38854
rect 5618 38820 5648 38854
rect 5690 38820 5717 38854
rect 5762 38820 5786 38854
rect 5834 38820 5855 38854
rect 5906 38820 5924 38854
rect 5978 38820 5993 38854
rect 6050 38820 6062 38854
rect 6122 38820 6131 38854
rect 6194 38820 6200 38854
rect 6266 38820 6268 38854
rect 6302 38820 6304 38854
rect 6370 38820 6376 38854
rect 6438 38820 6448 38854
rect 6506 38820 6520 38854
rect 6574 38820 6592 38854
rect 6642 38820 6664 38854
rect 6710 38820 6736 38854
rect 6778 38820 6808 38854
rect 6846 38820 6880 38854
rect 6914 38820 6948 38854
rect 6986 38820 7016 38854
rect 7058 38820 7084 38854
rect 7130 38820 7152 38854
rect 7202 38820 7220 38854
rect 7274 38820 7288 38854
rect 7346 38820 7356 38854
rect 7418 38820 7424 38854
rect 7490 38820 7492 38854
rect 7526 38820 7528 38854
rect 7594 38820 7600 38854
rect 7662 38820 7672 38854
rect 7730 38820 7744 38854
rect 7798 38820 7816 38854
rect 7866 38820 7888 38854
rect 7934 38820 7960 38854
rect 8002 38820 8032 38854
rect 8070 38820 8104 38854
rect 8138 38820 8172 38854
rect 8210 38820 8240 38854
rect 8282 38820 8308 38854
rect 8354 38820 8376 38854
rect 8426 38820 8444 38854
rect 8498 38820 8512 38854
rect 8570 38820 8580 38854
rect 8642 38820 8648 38854
rect 8714 38820 8716 38854
rect 8750 38820 8752 38854
rect 8818 38820 8824 38854
rect 8886 38820 8896 38854
rect 8954 38820 8968 38854
rect 9022 38820 9040 38854
rect 9090 38820 9112 38854
rect 9158 38820 9184 38854
rect 9226 38820 9256 38854
rect 9294 38820 9328 38854
rect 9362 38820 9396 38854
rect 9434 38820 9464 38854
rect 9506 38820 9532 38854
rect 9578 38820 9600 38854
rect 9650 38820 9668 38854
rect 9722 38820 9736 38854
rect 9794 38820 9804 38854
rect 9866 38820 9872 38854
rect 9938 38820 9940 38854
rect 9974 38820 9976 38854
rect 10042 38820 10048 38854
rect 10110 38820 10120 38854
rect 10178 38820 10192 38854
rect 10246 38820 10264 38854
rect 10314 38820 10336 38854
rect 10382 38820 10408 38854
rect 10450 38820 10480 38854
rect 10518 38820 10552 38854
rect 10586 38820 10620 38854
rect 10658 38820 10688 38854
rect 10730 38820 10756 38854
rect 10802 38820 10824 38854
rect 10874 38820 10892 38854
rect 10946 38820 10960 38854
rect 11018 38820 11028 38854
rect 11090 38820 11096 38854
rect 11162 38820 11164 38854
rect 11198 38820 11200 38854
rect 11266 38820 11272 38854
rect 11334 38820 11344 38854
rect 11402 38820 11416 38854
rect 11470 38820 11488 38854
rect 11538 38820 11560 38854
rect 11606 38820 11632 38854
rect 11674 38820 11704 38854
rect 11742 38820 11776 38854
rect 11810 38820 11844 38854
rect 11882 38820 11912 38854
rect 11954 38820 11980 38854
rect 12026 38820 12048 38854
rect 12098 38820 12116 38854
rect 12170 38820 12184 38854
rect 12242 38820 12252 38854
rect 12314 38820 12320 38854
rect 12386 38820 12388 38854
rect 12422 38820 12424 38854
rect 12490 38820 12496 38854
rect 12558 38820 12568 38854
rect 12626 38820 12640 38854
rect 12694 38820 12712 38854
rect 12762 38820 12784 38854
rect 12830 38820 12856 38854
rect 12898 38820 12928 38854
rect 12966 38820 13000 38854
rect 13034 38820 13068 38854
rect 13106 38820 13118 38854
rect 2213 38773 2219 38807
rect 2253 38773 2274 38807
rect 2213 38734 2274 38773
rect 2213 38700 2219 38734
rect 2253 38700 2274 38734
rect 2958 38714 3060 38726
rect 3512 38714 3614 38726
rect 4066 38714 4168 38726
rect 4620 38714 4722 38726
rect 5174 38714 5276 38726
rect 5728 38714 5830 38726
rect 6282 38714 6384 38726
rect 6836 38714 6938 38726
rect 7390 38714 7492 38726
rect 7944 38714 8046 38726
rect 8498 38714 8600 38726
rect 9052 38714 9154 38726
rect 9606 38714 9708 38726
rect 10160 38714 10262 38726
rect 10714 38714 10816 38726
rect 11268 38714 11370 38726
rect 11822 38714 11924 38726
rect 12376 38714 12478 38726
rect 12930 38714 13032 38726
rect 2213 38661 2274 38700
rect 2213 38627 2219 38661
rect 2253 38627 2274 38661
rect 2213 38588 2274 38627
rect 2213 38554 2219 38588
rect 2253 38554 2274 38588
rect 2213 38515 2274 38554
rect 2213 38481 2219 38515
rect 2253 38481 2274 38515
rect 2213 38442 2274 38481
rect 2213 38408 2219 38442
rect 2253 38408 2274 38442
rect 2213 38369 2274 38408
rect 2213 38335 2219 38369
rect 2253 38335 2274 38369
rect 2213 38296 2274 38335
rect 2213 38262 2219 38296
rect 2253 38262 2274 38296
rect 2213 38223 2274 38262
rect 2213 38189 2219 38223
rect 2253 38189 2274 38223
rect 2213 38150 2274 38189
rect 2213 38116 2219 38150
rect 2253 38116 2274 38150
rect 2213 38077 2274 38116
rect 2213 38043 2219 38077
rect 2253 38043 2274 38077
rect 2213 38004 2274 38043
rect 2213 37970 2219 38004
rect 2253 37970 2274 38004
rect 2213 37931 2274 37970
rect 2213 37897 2219 37931
rect 2253 37897 2274 37931
rect 2213 37858 2274 37897
rect 2213 37824 2219 37858
rect 2253 37824 2274 37858
rect 2213 37785 2274 37824
rect 2213 37751 2219 37785
rect 2253 37751 2274 37785
rect 2213 37712 2274 37751
rect 2213 37678 2219 37712
rect 2253 37678 2274 37712
rect 2213 37639 2274 37678
rect 2213 37605 2219 37639
rect 2253 37605 2274 37639
rect 2213 37566 2274 37605
rect 2213 37532 2219 37566
rect 2253 37532 2274 37566
rect 2213 37493 2274 37532
rect 2213 37459 2219 37493
rect 2253 37459 2274 37493
rect 2213 37420 2274 37459
rect 2213 37386 2219 37420
rect 2253 37386 2274 37420
rect 2213 37347 2274 37386
rect 2713 38680 2751 38714
rect 2679 38641 2785 38680
rect 2713 38607 2751 38641
rect 2679 38568 2785 38607
rect 2713 38534 2751 38568
rect 2679 38495 2785 38534
rect 2713 38461 2751 38495
rect 2679 38422 2785 38461
rect 2990 38680 3028 38714
rect 2956 38641 3062 38680
rect 2990 38607 3028 38641
rect 2956 38568 3062 38607
rect 2990 38534 3028 38568
rect 2956 38495 3062 38534
rect 2990 38461 3028 38495
rect 2956 38422 3062 38461
rect 3267 38680 3305 38714
rect 3233 38641 3339 38680
rect 3267 38607 3305 38641
rect 3233 38568 3339 38607
rect 3267 38534 3305 38568
rect 3233 38495 3339 38534
rect 3267 38461 3305 38495
rect 3233 38422 3339 38461
rect 3544 38680 3582 38714
rect 3510 38641 3616 38680
rect 3544 38607 3582 38641
rect 3510 38568 3616 38607
rect 3544 38534 3582 38568
rect 3510 38495 3616 38534
rect 3544 38461 3582 38495
rect 3510 38422 3616 38461
rect 3821 38680 3859 38714
rect 3787 38641 3893 38680
rect 3821 38607 3859 38641
rect 3787 38568 3893 38607
rect 3821 38534 3859 38568
rect 3787 38495 3893 38534
rect 3821 38461 3859 38495
rect 3787 38422 3893 38461
rect 4098 38680 4136 38714
rect 4064 38641 4170 38680
rect 4098 38607 4136 38641
rect 4064 38568 4170 38607
rect 4098 38534 4136 38568
rect 4064 38495 4170 38534
rect 4098 38461 4136 38495
rect 4064 38422 4170 38461
rect 4375 38680 4413 38714
rect 4341 38641 4447 38680
rect 4375 38607 4413 38641
rect 4341 38568 4447 38607
rect 4375 38534 4413 38568
rect 4341 38495 4447 38534
rect 4375 38461 4413 38495
rect 4341 38422 4447 38461
rect 4652 38680 4690 38714
rect 4618 38641 4724 38680
rect 4652 38607 4690 38641
rect 4618 38568 4724 38607
rect 4652 38534 4690 38568
rect 4618 38495 4724 38534
rect 4652 38461 4690 38495
rect 4618 38422 4724 38461
rect 4929 38680 4967 38714
rect 4895 38641 5001 38680
rect 4929 38607 4967 38641
rect 4895 38568 5001 38607
rect 4929 38534 4967 38568
rect 4895 38495 5001 38534
rect 4929 38461 4967 38495
rect 4895 38422 5001 38461
rect 5206 38680 5244 38714
rect 5172 38641 5278 38680
rect 5206 38607 5244 38641
rect 5172 38568 5278 38607
rect 5206 38534 5244 38568
rect 5172 38495 5278 38534
rect 5206 38461 5244 38495
rect 5172 38422 5278 38461
rect 5483 38680 5521 38714
rect 5449 38641 5555 38680
rect 5483 38607 5521 38641
rect 5449 38568 5555 38607
rect 5483 38534 5521 38568
rect 5449 38495 5555 38534
rect 5483 38461 5521 38495
rect 5449 38422 5555 38461
rect 5760 38680 5798 38714
rect 5726 38641 5832 38680
rect 5760 38607 5798 38641
rect 5726 38568 5832 38607
rect 5760 38534 5798 38568
rect 5726 38495 5832 38534
rect 5760 38461 5798 38495
rect 5726 38422 5832 38461
rect 6037 38680 6075 38714
rect 6003 38641 6109 38680
rect 6037 38607 6075 38641
rect 6003 38568 6109 38607
rect 6037 38534 6075 38568
rect 6003 38495 6109 38534
rect 6037 38461 6075 38495
rect 6003 38422 6109 38461
rect 6314 38680 6352 38714
rect 6280 38641 6386 38680
rect 6314 38607 6352 38641
rect 6280 38568 6386 38607
rect 6314 38534 6352 38568
rect 6280 38495 6386 38534
rect 6314 38461 6352 38495
rect 6280 38422 6386 38461
rect 6591 38680 6629 38714
rect 6557 38641 6663 38680
rect 6591 38607 6629 38641
rect 6557 38568 6663 38607
rect 6591 38534 6629 38568
rect 6557 38495 6663 38534
rect 6591 38461 6629 38495
rect 6557 38422 6663 38461
rect 6868 38680 6906 38714
rect 6834 38641 6940 38680
rect 6868 38607 6906 38641
rect 6834 38568 6940 38607
rect 6868 38534 6906 38568
rect 6834 38495 6940 38534
rect 6868 38461 6906 38495
rect 6834 38422 6940 38461
rect 7145 38680 7183 38714
rect 7111 38641 7217 38680
rect 7145 38607 7183 38641
rect 7111 38568 7217 38607
rect 7145 38534 7183 38568
rect 7111 38495 7217 38534
rect 7145 38461 7183 38495
rect 7111 38422 7217 38461
rect 7422 38680 7460 38714
rect 7388 38641 7494 38680
rect 7422 38607 7460 38641
rect 7388 38568 7494 38607
rect 7422 38534 7460 38568
rect 7388 38495 7494 38534
rect 7422 38461 7460 38495
rect 7388 38422 7494 38461
rect 7699 38680 7737 38714
rect 7665 38641 7771 38680
rect 7699 38607 7737 38641
rect 7665 38568 7771 38607
rect 7699 38534 7737 38568
rect 7665 38495 7771 38534
rect 7699 38461 7737 38495
rect 7665 38422 7771 38461
rect 7976 38680 8014 38714
rect 7942 38641 8048 38680
rect 7976 38607 8014 38641
rect 7942 38568 8048 38607
rect 7976 38534 8014 38568
rect 7942 38495 8048 38534
rect 7976 38461 8014 38495
rect 7942 38422 8048 38461
rect 8253 38680 8291 38714
rect 8219 38641 8325 38680
rect 8253 38607 8291 38641
rect 8219 38568 8325 38607
rect 8253 38534 8291 38568
rect 8219 38495 8325 38534
rect 8253 38461 8291 38495
rect 8219 38422 8325 38461
rect 8530 38680 8568 38714
rect 8496 38641 8602 38680
rect 8530 38607 8568 38641
rect 8496 38568 8602 38607
rect 8530 38534 8568 38568
rect 8496 38495 8602 38534
rect 8530 38461 8568 38495
rect 8496 38422 8602 38461
rect 8807 38680 8845 38714
rect 8773 38641 8879 38680
rect 8807 38607 8845 38641
rect 8773 38568 8879 38607
rect 8807 38534 8845 38568
rect 8773 38495 8879 38534
rect 8807 38461 8845 38495
rect 8773 38422 8879 38461
rect 9084 38680 9122 38714
rect 9050 38641 9156 38680
rect 9084 38607 9122 38641
rect 9050 38568 9156 38607
rect 9084 38534 9122 38568
rect 9050 38495 9156 38534
rect 9084 38461 9122 38495
rect 9050 38422 9156 38461
rect 9361 38680 9399 38714
rect 9327 38641 9433 38680
rect 9361 38607 9399 38641
rect 9327 38568 9433 38607
rect 9361 38534 9399 38568
rect 9327 38495 9433 38534
rect 9361 38461 9399 38495
rect 9327 38422 9433 38461
rect 9638 38680 9676 38714
rect 9604 38641 9710 38680
rect 9638 38607 9676 38641
rect 9604 38568 9710 38607
rect 9638 38534 9676 38568
rect 9604 38495 9710 38534
rect 9638 38461 9676 38495
rect 9604 38422 9710 38461
rect 9915 38680 9953 38714
rect 9881 38641 9987 38680
rect 9915 38607 9953 38641
rect 9881 38568 9987 38607
rect 9915 38534 9953 38568
rect 9881 38495 9987 38534
rect 9915 38461 9953 38495
rect 9881 38422 9987 38461
rect 10192 38680 10230 38714
rect 10158 38641 10264 38680
rect 10192 38607 10230 38641
rect 10158 38568 10264 38607
rect 10192 38534 10230 38568
rect 10158 38495 10264 38534
rect 10192 38461 10230 38495
rect 10158 38422 10264 38461
rect 10469 38680 10507 38714
rect 10435 38641 10541 38680
rect 10469 38607 10507 38641
rect 10435 38568 10541 38607
rect 10469 38534 10507 38568
rect 10435 38495 10541 38534
rect 10469 38461 10507 38495
rect 10435 38422 10541 38461
rect 10746 38680 10784 38714
rect 10712 38641 10818 38680
rect 10746 38607 10784 38641
rect 10712 38568 10818 38607
rect 10746 38534 10784 38568
rect 10712 38495 10818 38534
rect 10746 38461 10784 38495
rect 10712 38422 10818 38461
rect 11023 38680 11061 38714
rect 10989 38641 11095 38680
rect 11023 38607 11061 38641
rect 10989 38568 11095 38607
rect 11023 38534 11061 38568
rect 10989 38495 11095 38534
rect 11023 38461 11061 38495
rect 10989 38422 11095 38461
rect 11300 38680 11338 38714
rect 11266 38641 11372 38680
rect 11300 38607 11338 38641
rect 11266 38568 11372 38607
rect 11300 38534 11338 38568
rect 11266 38495 11372 38534
rect 11300 38461 11338 38495
rect 11266 38422 11372 38461
rect 11577 38680 11615 38714
rect 11543 38641 11649 38680
rect 11577 38607 11615 38641
rect 11543 38568 11649 38607
rect 11577 38534 11615 38568
rect 11543 38495 11649 38534
rect 11577 38461 11615 38495
rect 11543 38422 11649 38461
rect 11854 38680 11892 38714
rect 11820 38641 11926 38680
rect 11854 38607 11892 38641
rect 11820 38568 11926 38607
rect 11854 38534 11892 38568
rect 11820 38495 11926 38534
rect 11854 38461 11892 38495
rect 11820 38422 11926 38461
rect 12131 38680 12169 38714
rect 12097 38641 12203 38680
rect 12131 38607 12169 38641
rect 12097 38568 12203 38607
rect 12131 38534 12169 38568
rect 12097 38495 12203 38534
rect 12131 38461 12169 38495
rect 12097 38422 12203 38461
rect 12408 38680 12446 38714
rect 12374 38641 12480 38680
rect 12408 38607 12446 38641
rect 12374 38568 12480 38607
rect 12408 38534 12446 38568
rect 12374 38495 12480 38534
rect 12408 38461 12446 38495
rect 12374 38422 12480 38461
rect 12685 38680 12723 38714
rect 12651 38641 12757 38680
rect 12685 38607 12723 38641
rect 12651 38568 12757 38607
rect 12685 38534 12723 38568
rect 12651 38495 12757 38534
rect 12685 38461 12723 38495
rect 12651 38422 12757 38461
rect 12962 38680 13000 38714
rect 12928 38641 13034 38680
rect 12962 38607 13000 38641
rect 12928 38568 13034 38607
rect 12962 38534 13000 38568
rect 12928 38495 13034 38534
rect 12962 38461 13000 38495
rect 12928 38422 13034 38461
rect 13239 38680 13277 38714
rect 13205 38641 13311 38680
rect 13239 38607 13277 38641
rect 13205 38568 13311 38607
rect 13239 38534 13277 38568
rect 13205 38495 13311 38534
rect 13239 38461 13277 38495
rect 13205 38422 13311 38461
rect 2958 37368 3060 37380
rect 3512 37368 3614 37380
rect 4066 37368 4168 37380
rect 4620 37368 4722 37380
rect 5174 37368 5276 37380
rect 5728 37368 5830 37380
rect 6282 37368 6384 37380
rect 6836 37368 6938 37380
rect 7390 37368 7492 37380
rect 7944 37368 8046 37380
rect 8498 37368 8600 37380
rect 9052 37368 9154 37380
rect 9606 37368 9708 37380
rect 10160 37368 10262 37380
rect 10714 37368 10816 37380
rect 11268 37368 11370 37380
rect 11822 37368 11924 37380
rect 12376 37368 12478 37380
rect 12930 37368 13032 37380
rect 2213 37313 2219 37347
rect 2253 37313 2274 37347
rect 2213 37274 2274 37313
rect 2213 37240 2219 37274
rect 2253 37240 2274 37274
rect 2213 37201 2274 37240
rect 2213 37167 2219 37201
rect 2253 37167 2274 37201
rect 2213 37128 2274 37167
rect 2213 37094 2219 37128
rect 2253 37094 2274 37128
rect 2213 37055 2274 37094
rect 2213 37021 2219 37055
rect 2253 37021 2274 37055
rect 2213 36982 2274 37021
rect 2213 36948 2219 36982
rect 2253 36948 2274 36982
rect 2213 36909 2274 36948
rect 2213 36875 2219 36909
rect 2253 36875 2274 36909
rect 2213 36836 2274 36875
rect 2213 36802 2219 36836
rect 2253 36802 2274 36836
rect 2481 37290 2482 37324
rect 2516 37290 2568 37324
rect 2602 37290 2654 37324
rect 2688 37290 2740 37324
rect 2774 37290 2826 37324
rect 2860 37290 2888 37324
rect 2922 37290 2957 37324
rect 2991 37290 3026 37324
rect 3060 37290 3095 37324
rect 3129 37290 3164 37324
rect 3198 37290 3233 37324
rect 3267 37290 3302 37324
rect 3336 37290 3371 37324
rect 3405 37290 3440 37324
rect 3474 37290 3509 37324
rect 3543 37290 3578 37324
rect 3612 37290 3647 37324
rect 3681 37290 3716 37324
rect 3750 37290 3785 37324
rect 3819 37290 3854 37324
rect 3888 37290 3923 37324
rect 3957 37290 3992 37324
rect 4026 37290 4061 37324
rect 4095 37290 4130 37324
rect 4164 37290 4199 37324
rect 4233 37290 4268 37324
rect 4302 37290 4337 37324
rect 4371 37290 4406 37324
rect 4440 37290 4475 37324
rect 4509 37290 4544 37324
rect 4578 37290 4613 37324
rect 4647 37290 4682 37324
rect 4716 37290 4751 37324
rect 4785 37290 4820 37324
rect 4854 37290 4889 37324
rect 4923 37290 4958 37324
rect 4992 37290 5027 37324
rect 5061 37290 5096 37324
rect 5130 37290 5165 37324
rect 5199 37290 5234 37324
rect 5268 37290 5303 37324
rect 5337 37290 5372 37324
rect 5406 37290 5441 37324
rect 5475 37290 5510 37324
rect 5544 37290 5579 37324
rect 5613 37290 5648 37324
rect 5682 37290 5717 37324
rect 5751 37290 5786 37324
rect 5820 37290 5855 37324
rect 5889 37290 5924 37324
rect 5958 37290 5993 37324
rect 6027 37290 6062 37324
rect 6096 37290 6131 37324
rect 6165 37290 6200 37324
rect 6234 37290 6268 37324
rect 6302 37290 6336 37324
rect 6370 37290 6404 37324
rect 6438 37290 6472 37324
rect 6506 37290 6540 37324
rect 6574 37290 6608 37324
rect 6642 37290 6676 37324
rect 6710 37290 6744 37324
rect 6778 37290 6812 37324
rect 6846 37290 6880 37324
rect 6914 37290 6948 37324
rect 6982 37290 7016 37324
rect 7050 37290 7084 37324
rect 7118 37290 7152 37324
rect 7186 37290 7220 37324
rect 7254 37290 7288 37324
rect 7322 37290 7356 37324
rect 7390 37290 7424 37324
rect 7458 37290 7492 37324
rect 7526 37290 7560 37324
rect 7594 37290 7628 37324
rect 7662 37290 7696 37324
rect 7730 37290 7764 37324
rect 7798 37290 7832 37324
rect 7866 37290 7900 37324
rect 7934 37290 7968 37324
rect 8002 37290 8036 37324
rect 8070 37290 8104 37324
rect 8138 37290 8172 37324
rect 8206 37290 8240 37324
rect 8274 37290 8308 37324
rect 8342 37290 8376 37324
rect 8410 37290 8444 37324
rect 8478 37290 8512 37324
rect 8546 37290 8580 37324
rect 8614 37290 8648 37324
rect 8682 37290 8716 37324
rect 8750 37290 8784 37324
rect 8818 37290 8852 37324
rect 8886 37290 8920 37324
rect 8954 37290 8988 37324
rect 9022 37290 9056 37324
rect 9090 37290 9124 37324
rect 9158 37290 9192 37324
rect 9226 37290 9260 37324
rect 9294 37290 9328 37324
rect 9362 37290 9396 37324
rect 9430 37290 9464 37324
rect 9498 37290 9532 37324
rect 9566 37290 9600 37324
rect 9634 37290 9668 37324
rect 9702 37290 9736 37324
rect 9770 37290 9804 37324
rect 9838 37290 9872 37324
rect 9906 37290 9940 37324
rect 9974 37290 10008 37324
rect 10042 37290 10076 37324
rect 10110 37290 10144 37324
rect 10178 37290 10212 37324
rect 10246 37290 10280 37324
rect 10314 37290 10348 37324
rect 10382 37290 10416 37324
rect 10450 37290 10484 37324
rect 10518 37290 10552 37324
rect 10586 37290 10620 37324
rect 10654 37290 10688 37324
rect 10722 37290 10756 37324
rect 10790 37290 10824 37324
rect 10858 37290 10892 37324
rect 10926 37290 10960 37324
rect 10994 37290 11028 37324
rect 11062 37290 11096 37324
rect 11130 37290 11164 37324
rect 11198 37290 11232 37324
rect 11266 37290 11300 37324
rect 11334 37290 11368 37324
rect 11402 37290 11436 37324
rect 11470 37290 11504 37324
rect 11538 37290 11572 37324
rect 11606 37290 11640 37324
rect 11674 37290 11708 37324
rect 11742 37290 11776 37324
rect 11810 37290 11844 37324
rect 11878 37290 11912 37324
rect 11946 37290 11980 37324
rect 12014 37290 12048 37324
rect 12082 37290 12116 37324
rect 12150 37290 12184 37324
rect 12218 37290 12252 37324
rect 12286 37290 12320 37324
rect 12354 37290 12388 37324
rect 12422 37290 12456 37324
rect 12490 37290 12524 37324
rect 12558 37290 12592 37324
rect 12626 37290 12660 37324
rect 12694 37290 12728 37324
rect 12762 37290 12796 37324
rect 12830 37290 12864 37324
rect 12898 37290 12932 37324
rect 12966 37290 13000 37324
rect 13034 37290 13068 37324
rect 13102 37290 13315 37324
rect 2481 37247 13315 37290
rect 2481 37213 2482 37247
rect 2516 37213 2568 37247
rect 2602 37213 2654 37247
rect 2688 37213 2740 37247
rect 2774 37213 2826 37247
rect 2860 37213 13315 37247
rect 2481 37170 13315 37213
rect 2481 37136 2482 37170
rect 2516 37136 2568 37170
rect 2602 37136 2654 37170
rect 2688 37136 2740 37170
rect 2774 37136 2826 37170
rect 2860 37136 13315 37170
rect 2481 37093 13315 37136
rect 2481 37059 2482 37093
rect 2516 37059 2568 37093
rect 2602 37059 2654 37093
rect 2688 37059 2740 37093
rect 2774 37059 2826 37093
rect 2860 37059 13315 37093
rect 2481 37016 13315 37059
rect 2481 36982 2482 37016
rect 2516 36982 2568 37016
rect 2602 36982 2654 37016
rect 2688 36982 2740 37016
rect 2774 36982 2826 37016
rect 2860 36982 13315 37016
rect 2481 36939 13315 36982
rect 2481 36905 2482 36939
rect 2516 36905 2568 36939
rect 2602 36905 2654 36939
rect 2688 36905 2740 36939
rect 2774 36905 2826 36939
rect 2860 36905 13315 36939
rect 2481 36862 13315 36905
rect 2481 36828 2482 36862
rect 2516 36828 2568 36862
rect 2602 36828 2654 36862
rect 2688 36828 2740 36862
rect 2774 36828 2826 36862
rect 2860 36854 13315 36862
rect 2860 36828 2888 36854
rect 2486 36820 2888 36828
rect 2922 36820 2957 36854
rect 2991 36820 3026 36854
rect 3060 36820 3095 36854
rect 3129 36820 3164 36854
rect 3198 36820 3233 36854
rect 3267 36820 3302 36854
rect 3336 36820 3371 36854
rect 3405 36820 3440 36854
rect 3474 36820 3509 36854
rect 3543 36820 3578 36854
rect 3612 36820 3647 36854
rect 3681 36820 3716 36854
rect 3750 36820 3785 36854
rect 3819 36820 3854 36854
rect 3888 36820 3923 36854
rect 3957 36820 3992 36854
rect 4026 36820 4061 36854
rect 4095 36820 4130 36854
rect 4164 36820 4199 36854
rect 4233 36820 4268 36854
rect 4302 36820 4337 36854
rect 4371 36820 4406 36854
rect 4440 36820 4475 36854
rect 4509 36820 4544 36854
rect 4578 36820 4613 36854
rect 4647 36820 4682 36854
rect 4716 36820 4751 36854
rect 4785 36820 4820 36854
rect 4854 36820 4889 36854
rect 4923 36820 4958 36854
rect 4992 36820 5027 36854
rect 5061 36820 5096 36854
rect 5130 36820 5165 36854
rect 5199 36820 5234 36854
rect 5268 36820 5303 36854
rect 5337 36820 5372 36854
rect 5406 36820 5441 36854
rect 5475 36820 5510 36854
rect 5544 36820 5579 36854
rect 5613 36820 5648 36854
rect 5682 36820 5717 36854
rect 5751 36820 5786 36854
rect 5820 36820 5855 36854
rect 5889 36820 5924 36854
rect 5958 36820 5993 36854
rect 6027 36820 6062 36854
rect 6096 36820 6131 36854
rect 6165 36820 6200 36854
rect 6234 36820 6268 36854
rect 6302 36820 6336 36854
rect 6370 36820 6404 36854
rect 6438 36820 6472 36854
rect 6506 36820 6540 36854
rect 6574 36820 6608 36854
rect 6642 36820 6676 36854
rect 6710 36820 6744 36854
rect 6778 36820 6812 36854
rect 6846 36820 6880 36854
rect 6914 36820 6948 36854
rect 6982 36820 7016 36854
rect 7050 36820 7084 36854
rect 7118 36820 7152 36854
rect 7186 36820 7220 36854
rect 7254 36820 7288 36854
rect 7322 36820 7356 36854
rect 7390 36820 7424 36854
rect 7458 36820 7492 36854
rect 7526 36820 7560 36854
rect 7594 36820 7628 36854
rect 7662 36820 7696 36854
rect 7730 36820 7764 36854
rect 7798 36820 7832 36854
rect 7866 36820 7900 36854
rect 7934 36820 7968 36854
rect 8002 36820 8036 36854
rect 8070 36820 8104 36854
rect 8138 36820 8172 36854
rect 8206 36820 8240 36854
rect 8274 36820 8308 36854
rect 8342 36820 8376 36854
rect 8410 36820 8444 36854
rect 8478 36820 8512 36854
rect 8546 36820 8580 36854
rect 8614 36820 8648 36854
rect 8682 36820 8716 36854
rect 8750 36820 8784 36854
rect 8818 36820 8852 36854
rect 8886 36820 8920 36854
rect 8954 36820 8988 36854
rect 9022 36820 9056 36854
rect 9090 36820 9124 36854
rect 9158 36820 9192 36854
rect 9226 36820 9260 36854
rect 9294 36820 9328 36854
rect 9362 36820 9396 36854
rect 9430 36820 9464 36854
rect 9498 36820 9532 36854
rect 9566 36820 9600 36854
rect 9634 36820 9668 36854
rect 9702 36820 9736 36854
rect 9770 36820 9804 36854
rect 9838 36820 9872 36854
rect 9906 36820 9940 36854
rect 9974 36820 10008 36854
rect 10042 36820 10076 36854
rect 10110 36820 10144 36854
rect 10178 36820 10212 36854
rect 10246 36820 10280 36854
rect 10314 36820 10348 36854
rect 10382 36820 10416 36854
rect 10450 36820 10484 36854
rect 10518 36820 10552 36854
rect 10586 36820 10620 36854
rect 10654 36820 10688 36854
rect 10722 36820 10756 36854
rect 10790 36820 10824 36854
rect 10858 36820 10892 36854
rect 10926 36820 10960 36854
rect 10994 36820 11028 36854
rect 11062 36820 11096 36854
rect 11130 36820 11164 36854
rect 11198 36820 11232 36854
rect 11266 36820 11300 36854
rect 11334 36820 11368 36854
rect 11402 36820 11436 36854
rect 11470 36820 11504 36854
rect 11538 36820 11572 36854
rect 11606 36820 11640 36854
rect 11674 36820 11708 36854
rect 11742 36820 11776 36854
rect 11810 36820 11844 36854
rect 11878 36820 11912 36854
rect 11946 36820 11980 36854
rect 12014 36820 12048 36854
rect 12082 36820 12116 36854
rect 12150 36820 12184 36854
rect 12218 36820 12252 36854
rect 12286 36820 12320 36854
rect 12354 36820 12388 36854
rect 12422 36820 12456 36854
rect 12490 36820 12524 36854
rect 12558 36820 12592 36854
rect 12626 36820 12660 36854
rect 12694 36820 12728 36854
rect 12762 36820 12796 36854
rect 12830 36820 12864 36854
rect 12898 36820 12932 36854
rect 12966 36820 13000 36854
rect 13034 36820 13068 36854
rect 13102 36820 13315 36854
rect 2213 36763 2274 36802
rect 2213 36729 2219 36763
rect 2253 36729 2274 36763
rect 2213 36690 2274 36729
rect 3512 36714 3614 36726
rect 4066 36714 4168 36726
rect 4620 36714 4722 36726
rect 5174 36714 5276 36726
rect 5728 36714 5830 36726
rect 6282 36714 6384 36726
rect 6836 36714 6938 36726
rect 7390 36714 7492 36726
rect 7944 36714 8046 36726
rect 8498 36714 8600 36726
rect 9052 36714 9154 36726
rect 9606 36714 9708 36726
rect 10160 36714 10262 36726
rect 10714 36714 10816 36726
rect 11268 36714 11370 36726
rect 11822 36714 11924 36726
rect 12376 36714 12478 36726
rect 12930 36714 13032 36726
rect 2213 36656 2219 36690
rect 2253 36656 2274 36690
rect 2213 36617 2274 36656
rect 2213 36583 2219 36617
rect 2253 36583 2274 36617
rect 2213 36544 2274 36583
rect 2213 36510 2219 36544
rect 2253 36510 2274 36544
rect 2213 36471 2274 36510
rect 2213 36437 2219 36471
rect 2253 36437 2274 36471
rect 2213 36398 2274 36437
rect 2213 36364 2219 36398
rect 2253 36364 2274 36398
rect 2213 36325 2274 36364
rect 2213 36291 2219 36325
rect 2253 36291 2274 36325
rect 2213 36252 2274 36291
rect 2213 36218 2219 36252
rect 2253 36218 2274 36252
rect 2213 36179 2274 36218
rect 2213 36145 2219 36179
rect 2253 36145 2274 36179
rect 2213 36106 2274 36145
rect 2213 36072 2219 36106
rect 2253 36072 2274 36106
rect 2213 36033 2274 36072
rect 2213 35999 2219 36033
rect 2253 35999 2274 36033
rect 2213 35960 2274 35999
rect 2213 35926 2219 35960
rect 2253 35926 2274 35960
rect 2213 35887 2274 35926
rect 2213 35853 2219 35887
rect 2253 35853 2274 35887
rect 2213 35814 2274 35853
rect 2213 35780 2219 35814
rect 2253 35780 2274 35814
rect 2213 35741 2274 35780
rect 2213 35707 2219 35741
rect 2253 35707 2274 35741
rect 2213 35668 2274 35707
rect 2213 35634 2219 35668
rect 2253 35634 2274 35668
rect 2213 35595 2274 35634
rect 2213 35561 2219 35595
rect 2253 35561 2274 35595
rect 2213 35522 2274 35561
rect 2213 33688 2219 35522
rect 3267 36680 3305 36714
rect 3233 36641 3339 36680
rect 3267 36607 3305 36641
rect 3233 36568 3339 36607
rect 3267 36534 3305 36568
rect 3233 36495 3339 36534
rect 3267 36461 3305 36495
rect 3233 36422 3339 36461
rect 3544 36680 3582 36714
rect 3510 36641 3616 36680
rect 3544 36607 3582 36641
rect 3510 36568 3616 36607
rect 3544 36534 3582 36568
rect 3510 36495 3616 36534
rect 3544 36461 3582 36495
rect 3510 36422 3616 36461
rect 3821 36680 3859 36714
rect 3787 36641 3893 36680
rect 3821 36607 3859 36641
rect 3787 36568 3893 36607
rect 3821 36534 3859 36568
rect 3787 36495 3893 36534
rect 3821 36461 3859 36495
rect 3787 36422 3893 36461
rect 4098 36680 4136 36714
rect 4064 36641 4170 36680
rect 4098 36607 4136 36641
rect 4064 36568 4170 36607
rect 4098 36534 4136 36568
rect 4064 36495 4170 36534
rect 4098 36461 4136 36495
rect 4064 36422 4170 36461
rect 4375 36680 4413 36714
rect 4341 36641 4447 36680
rect 4375 36607 4413 36641
rect 4341 36568 4447 36607
rect 4375 36534 4413 36568
rect 4341 36495 4447 36534
rect 4375 36461 4413 36495
rect 4341 36422 4447 36461
rect 4652 36680 4690 36714
rect 4618 36641 4724 36680
rect 4652 36607 4690 36641
rect 4618 36568 4724 36607
rect 4652 36534 4690 36568
rect 4618 36495 4724 36534
rect 4652 36461 4690 36495
rect 4618 36422 4724 36461
rect 4929 36680 4967 36714
rect 4895 36641 5001 36680
rect 4929 36607 4967 36641
rect 4895 36568 5001 36607
rect 4929 36534 4967 36568
rect 4895 36495 5001 36534
rect 4929 36461 4967 36495
rect 4895 36422 5001 36461
rect 5206 36680 5244 36714
rect 5172 36641 5278 36680
rect 5206 36607 5244 36641
rect 5172 36568 5278 36607
rect 5206 36534 5244 36568
rect 5172 36495 5278 36534
rect 5206 36461 5244 36495
rect 5172 36422 5278 36461
rect 5483 36680 5521 36714
rect 5449 36641 5555 36680
rect 5483 36607 5521 36641
rect 5449 36568 5555 36607
rect 5483 36534 5521 36568
rect 5449 36495 5555 36534
rect 5483 36461 5521 36495
rect 5449 36422 5555 36461
rect 5760 36680 5798 36714
rect 5726 36641 5832 36680
rect 5760 36607 5798 36641
rect 5726 36568 5832 36607
rect 5760 36534 5798 36568
rect 5726 36495 5832 36534
rect 5760 36461 5798 36495
rect 5726 36422 5832 36461
rect 6037 36680 6075 36714
rect 6003 36641 6109 36680
rect 6037 36607 6075 36641
rect 6003 36568 6109 36607
rect 6037 36534 6075 36568
rect 6003 36495 6109 36534
rect 6037 36461 6075 36495
rect 6003 36422 6109 36461
rect 6314 36680 6352 36714
rect 6280 36641 6386 36680
rect 6314 36607 6352 36641
rect 6280 36568 6386 36607
rect 6314 36534 6352 36568
rect 6280 36495 6386 36534
rect 6314 36461 6352 36495
rect 6280 36422 6386 36461
rect 6591 36680 6629 36714
rect 6557 36641 6663 36680
rect 6591 36607 6629 36641
rect 6557 36568 6663 36607
rect 6591 36534 6629 36568
rect 6557 36495 6663 36534
rect 6591 36461 6629 36495
rect 6557 36422 6663 36461
rect 6868 36680 6906 36714
rect 6834 36641 6940 36680
rect 6868 36607 6906 36641
rect 6834 36568 6940 36607
rect 6868 36534 6906 36568
rect 6834 36495 6940 36534
rect 6868 36461 6906 36495
rect 6834 36422 6940 36461
rect 7145 36680 7183 36714
rect 7111 36641 7217 36680
rect 7145 36607 7183 36641
rect 7111 36568 7217 36607
rect 7145 36534 7183 36568
rect 7111 36495 7217 36534
rect 7145 36461 7183 36495
rect 7111 36422 7217 36461
rect 7422 36680 7460 36714
rect 7388 36641 7494 36680
rect 7422 36607 7460 36641
rect 7388 36568 7494 36607
rect 7422 36534 7460 36568
rect 7388 36495 7494 36534
rect 7422 36461 7460 36495
rect 7388 36422 7494 36461
rect 7699 36680 7737 36714
rect 7665 36641 7771 36680
rect 7699 36607 7737 36641
rect 7665 36568 7771 36607
rect 7699 36534 7737 36568
rect 7665 36495 7771 36534
rect 7699 36461 7737 36495
rect 7665 36422 7771 36461
rect 7976 36680 8014 36714
rect 7942 36641 8048 36680
rect 7976 36607 8014 36641
rect 7942 36568 8048 36607
rect 7976 36534 8014 36568
rect 7942 36495 8048 36534
rect 7976 36461 8014 36495
rect 7942 36422 8048 36461
rect 8253 36680 8291 36714
rect 8219 36641 8325 36680
rect 8253 36607 8291 36641
rect 8219 36568 8325 36607
rect 8253 36534 8291 36568
rect 8219 36495 8325 36534
rect 8253 36461 8291 36495
rect 8219 36422 8325 36461
rect 8530 36680 8568 36714
rect 8496 36641 8602 36680
rect 8530 36607 8568 36641
rect 8496 36568 8602 36607
rect 8530 36534 8568 36568
rect 8496 36495 8602 36534
rect 8530 36461 8568 36495
rect 8496 36422 8602 36461
rect 8807 36680 8845 36714
rect 8773 36641 8879 36680
rect 8807 36607 8845 36641
rect 8773 36568 8879 36607
rect 8807 36534 8845 36568
rect 8773 36495 8879 36534
rect 8807 36461 8845 36495
rect 8773 36422 8879 36461
rect 9084 36680 9122 36714
rect 9050 36641 9156 36680
rect 9084 36607 9122 36641
rect 9050 36568 9156 36607
rect 9084 36534 9122 36568
rect 9050 36495 9156 36534
rect 9084 36461 9122 36495
rect 9050 36422 9156 36461
rect 9361 36680 9399 36714
rect 9327 36641 9433 36680
rect 9361 36607 9399 36641
rect 9327 36568 9433 36607
rect 9361 36534 9399 36568
rect 9327 36495 9433 36534
rect 9361 36461 9399 36495
rect 9327 36422 9433 36461
rect 9638 36680 9676 36714
rect 9604 36641 9710 36680
rect 9638 36607 9676 36641
rect 9604 36568 9710 36607
rect 9638 36534 9676 36568
rect 9604 36495 9710 36534
rect 9638 36461 9676 36495
rect 9604 36422 9710 36461
rect 9915 36680 9953 36714
rect 9881 36641 9987 36680
rect 9915 36607 9953 36641
rect 9881 36568 9987 36607
rect 9915 36534 9953 36568
rect 9881 36495 9987 36534
rect 9915 36461 9953 36495
rect 9881 36422 9987 36461
rect 10192 36680 10230 36714
rect 10158 36641 10264 36680
rect 10192 36607 10230 36641
rect 10158 36568 10264 36607
rect 10192 36534 10230 36568
rect 10158 36495 10264 36534
rect 10192 36461 10230 36495
rect 10158 36422 10264 36461
rect 10469 36680 10507 36714
rect 10435 36641 10541 36680
rect 10469 36607 10507 36641
rect 10435 36568 10541 36607
rect 10469 36534 10507 36568
rect 10435 36495 10541 36534
rect 10469 36461 10507 36495
rect 10435 36422 10541 36461
rect 10746 36680 10784 36714
rect 10712 36641 10818 36680
rect 10746 36607 10784 36641
rect 10712 36568 10818 36607
rect 10746 36534 10784 36568
rect 10712 36495 10818 36534
rect 10746 36461 10784 36495
rect 10712 36422 10818 36461
rect 11023 36680 11061 36714
rect 10989 36641 11095 36680
rect 11023 36607 11061 36641
rect 10989 36568 11095 36607
rect 11023 36534 11061 36568
rect 10989 36495 11095 36534
rect 11023 36461 11061 36495
rect 10989 36422 11095 36461
rect 11300 36680 11338 36714
rect 11266 36641 11372 36680
rect 11300 36607 11338 36641
rect 11266 36568 11372 36607
rect 11300 36534 11338 36568
rect 11266 36495 11372 36534
rect 11300 36461 11338 36495
rect 11266 36422 11372 36461
rect 11577 36680 11615 36714
rect 11543 36641 11649 36680
rect 11577 36607 11615 36641
rect 11543 36568 11649 36607
rect 11577 36534 11615 36568
rect 11543 36495 11649 36534
rect 11577 36461 11615 36495
rect 11543 36422 11649 36461
rect 11854 36680 11892 36714
rect 11820 36641 11926 36680
rect 11854 36607 11892 36641
rect 11820 36568 11926 36607
rect 11854 36534 11892 36568
rect 11820 36495 11926 36534
rect 11854 36461 11892 36495
rect 11820 36422 11926 36461
rect 12131 36680 12169 36714
rect 12097 36641 12203 36680
rect 12131 36607 12169 36641
rect 12097 36568 12203 36607
rect 12131 36534 12169 36568
rect 12097 36495 12203 36534
rect 12131 36461 12169 36495
rect 12097 36422 12203 36461
rect 12408 36680 12446 36714
rect 12374 36641 12480 36680
rect 12408 36607 12446 36641
rect 12374 36568 12480 36607
rect 12408 36534 12446 36568
rect 12374 36495 12480 36534
rect 12408 36461 12446 36495
rect 12374 36422 12480 36461
rect 12685 36680 12723 36714
rect 12651 36641 12757 36680
rect 12685 36607 12723 36641
rect 12651 36568 12757 36607
rect 12685 36534 12723 36568
rect 12651 36495 12757 36534
rect 12685 36461 12723 36495
rect 12651 36422 12757 36461
rect 12962 36680 13000 36714
rect 12928 36641 13034 36680
rect 12962 36607 13000 36641
rect 12928 36568 13034 36607
rect 12962 36534 13000 36568
rect 12928 36495 13034 36534
rect 12962 36461 13000 36495
rect 12928 36422 13034 36461
rect 13239 36680 13277 36714
rect 13205 36641 13311 36680
rect 13239 36607 13277 36641
rect 13205 36568 13311 36607
rect 13239 36534 13277 36568
rect 13205 36495 13311 36534
rect 13239 36461 13277 36495
rect 13205 36422 13311 36461
rect 3512 35368 3614 35380
rect 4066 35368 4168 35380
rect 4620 35368 4722 35380
rect 5174 35368 5276 35380
rect 5728 35368 5830 35380
rect 6282 35368 6384 35380
rect 6836 35368 6938 35380
rect 7390 35368 7492 35380
rect 7944 35368 8046 35380
rect 8498 35368 8600 35380
rect 9052 35368 9154 35380
rect 9606 35368 9708 35380
rect 10160 35368 10262 35380
rect 10714 35368 10816 35380
rect 11268 35368 11370 35380
rect 11822 35368 11924 35380
rect 12376 35368 12478 35380
rect 12930 35368 13032 35380
rect 2667 35321 2888 35324
rect 2667 35287 2674 35321
rect 2708 35287 2750 35321
rect 2784 35287 2826 35321
rect 2860 35290 2888 35321
rect 2922 35290 2957 35324
rect 2991 35290 3026 35324
rect 3060 35290 3095 35324
rect 3129 35290 3164 35324
rect 3198 35290 3233 35324
rect 3267 35290 3302 35324
rect 3336 35290 3371 35324
rect 3405 35290 3440 35324
rect 3474 35290 3509 35324
rect 3543 35290 3578 35324
rect 3612 35290 3647 35324
rect 3681 35290 3716 35324
rect 3750 35290 3785 35324
rect 3819 35290 3854 35324
rect 3888 35290 3923 35324
rect 3957 35290 3992 35324
rect 4026 35290 4061 35324
rect 4095 35290 4130 35324
rect 4164 35290 4199 35324
rect 4233 35290 4268 35324
rect 4302 35290 4337 35324
rect 4371 35290 4406 35324
rect 4440 35290 4475 35324
rect 4509 35290 4544 35324
rect 4578 35290 4613 35324
rect 4647 35290 4682 35324
rect 4716 35290 4751 35324
rect 4785 35290 4820 35324
rect 4854 35290 4889 35324
rect 4923 35290 4958 35324
rect 4992 35290 5027 35324
rect 5061 35290 5096 35324
rect 5130 35290 5165 35324
rect 5199 35290 5234 35324
rect 5268 35290 5303 35324
rect 5337 35290 5372 35324
rect 5406 35290 5441 35324
rect 5475 35290 5510 35324
rect 5544 35290 5579 35324
rect 5613 35290 5648 35324
rect 5682 35290 5717 35324
rect 5751 35290 5786 35324
rect 5820 35290 5855 35324
rect 5889 35290 5924 35324
rect 5958 35290 5993 35324
rect 6027 35290 6062 35324
rect 6096 35290 6131 35324
rect 6165 35290 6200 35324
rect 6234 35290 6268 35324
rect 6302 35290 6336 35324
rect 6370 35290 6404 35324
rect 6438 35290 6472 35324
rect 6506 35290 6540 35324
rect 6574 35290 6608 35324
rect 6642 35290 6676 35324
rect 6710 35290 6744 35324
rect 6778 35290 6812 35324
rect 6846 35290 6880 35324
rect 6914 35290 6948 35324
rect 6982 35290 7016 35324
rect 7050 35290 7084 35324
rect 7118 35290 7152 35324
rect 7186 35290 7220 35324
rect 7254 35290 7288 35324
rect 7322 35290 7356 35324
rect 7390 35290 7424 35324
rect 7458 35290 7492 35324
rect 7526 35290 7560 35324
rect 7594 35290 7628 35324
rect 7662 35290 7696 35324
rect 7730 35290 7764 35324
rect 7798 35290 7832 35324
rect 7866 35290 7900 35324
rect 7934 35290 7968 35324
rect 8002 35290 8036 35324
rect 8070 35290 8104 35324
rect 8138 35290 8172 35324
rect 8206 35290 8240 35324
rect 8274 35290 8308 35324
rect 8342 35290 8376 35324
rect 8410 35290 8444 35324
rect 8478 35290 8512 35324
rect 8546 35290 8580 35324
rect 8614 35290 8648 35324
rect 8682 35290 8716 35324
rect 8750 35290 8784 35324
rect 8818 35290 8852 35324
rect 8886 35290 8920 35324
rect 8954 35290 8988 35324
rect 9022 35290 9056 35324
rect 9090 35290 9124 35324
rect 9158 35290 9192 35324
rect 9226 35290 9260 35324
rect 9294 35290 9328 35324
rect 9362 35290 9396 35324
rect 9430 35290 9464 35324
rect 9498 35290 9532 35324
rect 9566 35290 9600 35324
rect 9634 35290 9668 35324
rect 9702 35290 9736 35324
rect 9770 35290 9804 35324
rect 9838 35290 9872 35324
rect 9906 35290 9940 35324
rect 9974 35290 10008 35324
rect 10042 35290 10076 35324
rect 10110 35290 10144 35324
rect 10178 35290 10212 35324
rect 10246 35290 10280 35324
rect 10314 35290 10348 35324
rect 10382 35290 10416 35324
rect 10450 35290 10484 35324
rect 10518 35290 10552 35324
rect 10586 35290 10620 35324
rect 10654 35290 10688 35324
rect 10722 35290 10756 35324
rect 10790 35290 10824 35324
rect 10858 35290 10892 35324
rect 10926 35290 10960 35324
rect 10994 35290 11028 35324
rect 11062 35290 11096 35324
rect 11130 35290 11164 35324
rect 11198 35290 11232 35324
rect 11266 35290 11300 35324
rect 11334 35290 11368 35324
rect 11402 35290 11436 35324
rect 11470 35290 11504 35324
rect 11538 35290 11572 35324
rect 11606 35290 11640 35324
rect 11674 35290 11708 35324
rect 11742 35290 11776 35324
rect 11810 35290 11844 35324
rect 11878 35290 11912 35324
rect 11946 35290 11980 35324
rect 12014 35290 12048 35324
rect 12082 35290 12116 35324
rect 12150 35290 12184 35324
rect 12218 35290 12252 35324
rect 12286 35290 12320 35324
rect 12354 35290 12388 35324
rect 12422 35290 12456 35324
rect 12490 35290 12524 35324
rect 12558 35290 12592 35324
rect 12626 35290 12660 35324
rect 12694 35290 12728 35324
rect 12762 35290 12796 35324
rect 12830 35290 12864 35324
rect 12898 35290 12932 35324
rect 12966 35290 13000 35324
rect 13034 35290 13068 35324
rect 13102 35290 13118 35324
rect 2860 35287 13118 35290
rect 2667 35244 13118 35287
rect 2667 35210 2674 35244
rect 2708 35210 2750 35244
rect 2784 35210 2826 35244
rect 2860 35210 13118 35244
rect 2667 35167 13118 35210
rect 2667 35133 2674 35167
rect 2708 35133 2750 35167
rect 2784 35133 2826 35167
rect 2860 35133 13118 35167
rect 2667 35089 13118 35133
rect 2667 35055 2674 35089
rect 2708 35055 2750 35089
rect 2784 35055 2826 35089
rect 2860 35055 13118 35089
rect 2667 35011 13118 35055
rect 2667 34977 2674 35011
rect 2708 34977 2750 35011
rect 2784 34977 2826 35011
rect 2860 34977 13118 35011
rect 2667 34933 13118 34977
rect 2667 34899 2674 34933
rect 2708 34899 2750 34933
rect 2784 34899 2826 34933
rect 2860 34899 13118 34933
rect 2667 34855 13118 34899
rect 2667 34821 2674 34855
rect 2708 34821 2750 34855
rect 2784 34821 2826 34855
rect 2860 34854 13118 34855
rect 2860 34821 3507 34854
rect 2667 34820 3507 34821
rect 3541 34820 3576 34854
rect 3610 34820 3645 34854
rect 3679 34820 3714 34854
rect 3748 34820 3783 34854
rect 3817 34820 3852 34854
rect 3886 34820 3921 34854
rect 3955 34820 3990 34854
rect 4024 34820 4059 34854
rect 4093 34820 4128 34854
rect 4162 34820 4197 34854
rect 4231 34820 4266 34854
rect 4300 34820 4335 34854
rect 4369 34820 4404 34854
rect 4438 34820 4473 34854
rect 4507 34820 4542 34854
rect 4576 34820 4611 34854
rect 4645 34820 4680 34854
rect 4714 34820 4749 34854
rect 4783 34820 4818 34854
rect 4852 34820 4887 34854
rect 4921 34820 4956 34854
rect 4990 34820 5025 34854
rect 5059 34820 5094 34854
rect 5128 34820 5163 34854
rect 5197 34820 5232 34854
rect 5266 34820 5301 34854
rect 5335 34820 5370 34854
rect 5404 34820 5439 34854
rect 5473 34820 5508 34854
rect 5542 34820 5577 34854
rect 5611 34820 5646 34854
rect 5680 34820 5715 34854
rect 5749 34820 5784 34854
rect 5818 34820 5853 34854
rect 5887 34820 5922 34854
rect 5956 34820 5991 34854
rect 6025 34820 6060 34854
rect 6094 34820 6129 34854
rect 6163 34820 6198 34854
rect 6232 34820 6267 34854
rect 6301 34820 6336 34854
rect 6370 34820 6405 34854
rect 6439 34820 6474 34854
rect 6508 34820 6543 34854
rect 6577 34820 6612 34854
rect 6646 34820 6681 34854
rect 6715 34820 6750 34854
rect 6784 34820 6819 34854
rect 6853 34820 6888 34854
rect 6922 34820 6957 34854
rect 6991 34820 7026 34854
rect 7060 34820 7095 34854
rect 7129 34820 7163 34854
rect 7197 34820 7231 34854
rect 7265 34820 7299 34854
rect 7333 34820 7367 34854
rect 7401 34820 7435 34854
rect 7469 34820 7503 34854
rect 7537 34820 7571 34854
rect 7605 34820 7639 34854
rect 7673 34820 7707 34854
rect 7741 34820 7775 34854
rect 7809 34820 7843 34854
rect 7877 34820 7911 34854
rect 7945 34820 7979 34854
rect 8013 34820 8047 34854
rect 8081 34820 8115 34854
rect 8149 34820 8183 34854
rect 8217 34820 8251 34854
rect 8285 34820 8319 34854
rect 8353 34820 8387 34854
rect 8421 34820 8455 34854
rect 8489 34820 8523 34854
rect 8557 34820 8591 34854
rect 8625 34820 8659 34854
rect 8693 34820 8727 34854
rect 8761 34820 8795 34854
rect 8829 34820 8863 34854
rect 8897 34820 8931 34854
rect 8965 34820 8999 34854
rect 9033 34820 9067 34854
rect 9101 34820 9135 34854
rect 9169 34820 9203 34854
rect 9237 34820 9271 34854
rect 9305 34820 9339 34854
rect 9373 34820 9407 34854
rect 9441 34820 9475 34854
rect 9509 34820 9543 34854
rect 9577 34820 9611 34854
rect 9645 34820 9679 34854
rect 9713 34820 9747 34854
rect 9781 34820 9815 34854
rect 9849 34820 9883 34854
rect 9917 34820 9951 34854
rect 9985 34820 10019 34854
rect 10053 34820 10087 34854
rect 10121 34820 10155 34854
rect 10189 34820 10223 34854
rect 10257 34820 10291 34854
rect 10325 34820 10359 34854
rect 10393 34820 10427 34854
rect 10461 34820 10495 34854
rect 10529 34820 10563 34854
rect 10597 34820 10631 34854
rect 10665 34820 10699 34854
rect 10733 34820 10767 34854
rect 10801 34820 10835 34854
rect 10869 34820 10903 34854
rect 10937 34820 10971 34854
rect 11005 34820 11039 34854
rect 11073 34820 11107 34854
rect 11141 34820 11175 34854
rect 11209 34820 11243 34854
rect 11277 34820 11311 34854
rect 11345 34820 11379 34854
rect 11413 34820 11447 34854
rect 11481 34820 11515 34854
rect 11549 34820 11583 34854
rect 11617 34820 11651 34854
rect 11685 34820 11719 34854
rect 11753 34820 11787 34854
rect 11821 34820 11855 34854
rect 11889 34820 11923 34854
rect 11957 34820 11991 34854
rect 12025 34820 12059 34854
rect 12093 34820 12127 34854
rect 12161 34820 12195 34854
rect 12229 34820 12263 34854
rect 12297 34820 12331 34854
rect 12365 34820 12399 34854
rect 12433 34820 12467 34854
rect 12501 34820 12535 34854
rect 12569 34820 12603 34854
rect 12637 34820 12671 34854
rect 12705 34820 12739 34854
rect 12773 34820 12807 34854
rect 12841 34820 12875 34854
rect 12909 34820 12943 34854
rect 12977 34820 13118 34854
rect 3593 34714 3695 34726
rect 4429 34714 4531 34726
rect 5265 34714 5367 34726
rect 6101 34714 6203 34726
rect 6937 34714 7039 34726
rect 7773 34714 7875 34726
rect 8609 34714 8711 34726
rect 9445 34714 9547 34726
rect 10281 34714 10383 34726
rect 11117 34714 11219 34726
rect 11953 34714 12055 34726
rect 12789 34714 12891 34726
rect 2213 33656 2274 33688
rect 2219 33644 2274 33656
rect 2253 33610 2274 33644
rect 2219 33571 2274 33610
rect 2253 33537 2274 33571
rect 2219 33498 2274 33537
rect 2253 33464 2274 33498
rect 2219 33425 2274 33464
rect 2253 33391 2274 33425
rect 2219 33352 2274 33391
rect 3207 34680 3245 34714
rect 3173 34641 3279 34680
rect 3207 34607 3245 34641
rect 3173 34568 3279 34607
rect 3207 34534 3245 34568
rect 3173 34495 3279 34534
rect 3207 34461 3245 34495
rect 3173 34422 3279 34461
rect 3625 34680 3663 34714
rect 3591 34641 3697 34680
rect 3625 34607 3663 34641
rect 3591 34568 3697 34607
rect 3625 34534 3663 34568
rect 3591 34495 3697 34534
rect 3625 34461 3663 34495
rect 3591 34422 3697 34461
rect 4043 34680 4081 34714
rect 4009 34641 4115 34680
rect 4043 34607 4081 34641
rect 4009 34568 4115 34607
rect 4043 34534 4081 34568
rect 4009 34495 4115 34534
rect 4043 34461 4081 34495
rect 4009 34422 4115 34461
rect 4461 34680 4499 34714
rect 4427 34641 4533 34680
rect 4461 34607 4499 34641
rect 4427 34568 4533 34607
rect 4461 34534 4499 34568
rect 4427 34495 4533 34534
rect 4461 34461 4499 34495
rect 4427 34422 4533 34461
rect 4879 34680 4917 34714
rect 4845 34641 4951 34680
rect 4879 34607 4917 34641
rect 4845 34568 4951 34607
rect 4879 34534 4917 34568
rect 4845 34495 4951 34534
rect 4879 34461 4917 34495
rect 4845 34422 4951 34461
rect 5297 34680 5335 34714
rect 5263 34641 5369 34680
rect 5297 34607 5335 34641
rect 5263 34568 5369 34607
rect 5297 34534 5335 34568
rect 5263 34495 5369 34534
rect 5297 34461 5335 34495
rect 5263 34422 5369 34461
rect 5715 34680 5753 34714
rect 5681 34641 5787 34680
rect 5715 34607 5753 34641
rect 5681 34568 5787 34607
rect 5715 34534 5753 34568
rect 5681 34495 5787 34534
rect 5715 34461 5753 34495
rect 5681 34422 5787 34461
rect 6133 34680 6171 34714
rect 6099 34641 6205 34680
rect 6133 34607 6171 34641
rect 6099 34568 6205 34607
rect 6133 34534 6171 34568
rect 6099 34495 6205 34534
rect 6133 34461 6171 34495
rect 6099 34422 6205 34461
rect 6551 34680 6589 34714
rect 6517 34641 6623 34680
rect 6551 34607 6589 34641
rect 6517 34568 6623 34607
rect 6551 34534 6589 34568
rect 6517 34495 6623 34534
rect 6551 34461 6589 34495
rect 6517 34422 6623 34461
rect 6969 34680 7007 34714
rect 6935 34641 7041 34680
rect 6969 34607 7007 34641
rect 6935 34568 7041 34607
rect 6969 34534 7007 34568
rect 6935 34495 7041 34534
rect 6969 34461 7007 34495
rect 6935 34422 7041 34461
rect 7387 34680 7425 34714
rect 7353 34641 7459 34680
rect 7387 34607 7425 34641
rect 7353 34568 7459 34607
rect 7387 34534 7425 34568
rect 7353 34495 7459 34534
rect 7387 34461 7425 34495
rect 7353 34422 7459 34461
rect 7805 34680 7843 34714
rect 7771 34641 7877 34680
rect 7805 34607 7843 34641
rect 7771 34568 7877 34607
rect 7805 34534 7843 34568
rect 7771 34495 7877 34534
rect 7805 34461 7843 34495
rect 7771 34422 7877 34461
rect 8223 34680 8261 34714
rect 8189 34641 8295 34680
rect 8223 34607 8261 34641
rect 8189 34568 8295 34607
rect 8223 34534 8261 34568
rect 8189 34495 8295 34534
rect 8223 34461 8261 34495
rect 8189 34422 8295 34461
rect 8641 34680 8679 34714
rect 8607 34641 8713 34680
rect 8641 34607 8679 34641
rect 8607 34568 8713 34607
rect 8641 34534 8679 34568
rect 8607 34495 8713 34534
rect 8641 34461 8679 34495
rect 8607 34422 8713 34461
rect 9059 34680 9097 34714
rect 9025 34641 9131 34680
rect 9059 34607 9097 34641
rect 9025 34568 9131 34607
rect 9059 34534 9097 34568
rect 9025 34495 9131 34534
rect 9059 34461 9097 34495
rect 9025 34422 9131 34461
rect 9477 34680 9515 34714
rect 9443 34641 9549 34680
rect 9477 34607 9515 34641
rect 9443 34568 9549 34607
rect 9477 34534 9515 34568
rect 9443 34495 9549 34534
rect 9477 34461 9515 34495
rect 9443 34422 9549 34461
rect 9895 34680 9933 34714
rect 9861 34641 9967 34680
rect 9895 34607 9933 34641
rect 9861 34568 9967 34607
rect 9895 34534 9933 34568
rect 9861 34495 9967 34534
rect 9895 34461 9933 34495
rect 9861 34422 9967 34461
rect 10313 34680 10351 34714
rect 10279 34641 10385 34680
rect 10313 34607 10351 34641
rect 10279 34568 10385 34607
rect 10313 34534 10351 34568
rect 10279 34495 10385 34534
rect 10313 34461 10351 34495
rect 10279 34422 10385 34461
rect 10731 34680 10769 34714
rect 10697 34641 10803 34680
rect 10731 34607 10769 34641
rect 10697 34568 10803 34607
rect 10731 34534 10769 34568
rect 10697 34495 10803 34534
rect 10731 34461 10769 34495
rect 10697 34422 10803 34461
rect 11149 34680 11187 34714
rect 11115 34641 11221 34680
rect 11149 34607 11187 34641
rect 11115 34568 11221 34607
rect 11149 34534 11187 34568
rect 11115 34495 11221 34534
rect 11149 34461 11187 34495
rect 11115 34422 11221 34461
rect 11567 34680 11605 34714
rect 11533 34641 11639 34680
rect 11567 34607 11605 34641
rect 11533 34568 11639 34607
rect 11567 34534 11605 34568
rect 11533 34495 11639 34534
rect 11567 34461 11605 34495
rect 11533 34422 11639 34461
rect 11985 34680 12023 34714
rect 11951 34641 12057 34680
rect 11985 34607 12023 34641
rect 11951 34568 12057 34607
rect 11985 34534 12023 34568
rect 11951 34495 12057 34534
rect 11985 34461 12023 34495
rect 11951 34422 12057 34461
rect 12403 34680 12441 34714
rect 12369 34641 12475 34680
rect 12403 34607 12441 34641
rect 12369 34568 12475 34607
rect 12403 34534 12441 34568
rect 12369 34495 12475 34534
rect 12403 34461 12441 34495
rect 12369 34422 12475 34461
rect 12821 34680 12859 34714
rect 12787 34641 12893 34680
rect 12821 34607 12859 34641
rect 12787 34568 12893 34607
rect 12821 34534 12859 34568
rect 12787 34495 12893 34534
rect 12821 34461 12859 34495
rect 12787 34422 12893 34461
rect 13239 34680 13277 34714
rect 13205 34641 13311 34680
rect 13239 34607 13277 34641
rect 13205 34568 13311 34607
rect 13239 34534 13277 34568
rect 13205 34495 13311 34534
rect 13239 34461 13277 34495
rect 13205 34422 13311 34461
rect 3593 33368 3695 33380
rect 4429 33368 4531 33380
rect 5265 33368 5367 33380
rect 6101 33368 6203 33380
rect 6937 33368 7039 33380
rect 7773 33368 7875 33380
rect 8609 33368 8711 33380
rect 9445 33368 9547 33380
rect 10281 33368 10383 33380
rect 11117 33368 11219 33380
rect 11953 33368 12055 33380
rect 12789 33368 12891 33380
rect 2253 33318 2274 33352
rect 2219 33279 2274 33318
rect 2253 33245 2274 33279
rect 2219 33206 2274 33245
rect 2253 33172 2274 33206
rect 2219 33133 2274 33172
rect 2253 33099 2274 33133
rect 2219 33060 2274 33099
rect 2253 33026 2274 33060
rect 2219 32987 2274 33026
rect 2253 32953 2274 32987
rect 2219 32914 2274 32953
rect 2253 32880 2274 32914
rect 2219 32841 2274 32880
rect 2253 32807 2274 32841
rect 2673 33322 3507 33324
rect 2673 33288 2674 33322
rect 2708 33288 2750 33322
rect 2784 33288 2826 33322
rect 2860 33290 3507 33322
rect 3541 33290 3576 33324
rect 3610 33290 3645 33324
rect 3679 33290 3714 33324
rect 3748 33290 3783 33324
rect 3817 33290 3852 33324
rect 3886 33290 3921 33324
rect 3955 33290 3990 33324
rect 4024 33290 4059 33324
rect 4093 33290 4128 33324
rect 4162 33290 4197 33324
rect 4231 33290 4266 33324
rect 4300 33290 4335 33324
rect 4369 33290 4404 33324
rect 4438 33290 4473 33324
rect 4507 33290 4542 33324
rect 4576 33290 4611 33324
rect 4645 33290 4680 33324
rect 4714 33290 4749 33324
rect 4783 33290 4818 33324
rect 4852 33290 4887 33324
rect 4921 33290 4956 33324
rect 4990 33290 5025 33324
rect 5059 33290 5094 33324
rect 5128 33290 5163 33324
rect 5197 33290 5232 33324
rect 5266 33290 5301 33324
rect 5335 33290 5370 33324
rect 5404 33290 5439 33324
rect 5473 33290 5508 33324
rect 5542 33290 5577 33324
rect 5611 33290 5646 33324
rect 5680 33290 5715 33324
rect 5749 33290 5784 33324
rect 5818 33290 5853 33324
rect 5887 33290 5922 33324
rect 5956 33290 5991 33324
rect 6025 33290 6060 33324
rect 6094 33290 6129 33324
rect 6163 33290 6198 33324
rect 6232 33290 6267 33324
rect 6301 33290 6336 33324
rect 6370 33290 6405 33324
rect 6439 33290 6474 33324
rect 6508 33290 6543 33324
rect 6577 33290 6612 33324
rect 6646 33290 6681 33324
rect 6715 33290 6750 33324
rect 6784 33290 6819 33324
rect 6853 33290 6888 33324
rect 6922 33290 6957 33324
rect 6991 33290 7026 33324
rect 7060 33290 7095 33324
rect 7129 33290 7163 33324
rect 7197 33290 7231 33324
rect 7265 33290 7299 33324
rect 7333 33290 7367 33324
rect 7401 33290 7435 33324
rect 7469 33290 7503 33324
rect 7537 33290 7571 33324
rect 7605 33290 7639 33324
rect 7673 33290 7707 33324
rect 7741 33290 7775 33324
rect 7809 33290 7843 33324
rect 7877 33290 7911 33324
rect 7945 33290 7979 33324
rect 8013 33290 8047 33324
rect 8081 33290 8115 33324
rect 8149 33290 8183 33324
rect 8217 33290 8251 33324
rect 8285 33290 8319 33324
rect 8353 33290 8387 33324
rect 8421 33290 8455 33324
rect 8489 33290 8523 33324
rect 8557 33290 8591 33324
rect 8625 33290 8659 33324
rect 8693 33290 8727 33324
rect 8761 33290 8795 33324
rect 8829 33290 8863 33324
rect 8897 33290 8931 33324
rect 8965 33290 8999 33324
rect 9033 33290 9067 33324
rect 9101 33290 9135 33324
rect 9169 33290 9203 33324
rect 9237 33290 9271 33324
rect 9305 33290 9339 33324
rect 9373 33290 9407 33324
rect 9441 33290 9475 33324
rect 9509 33290 9543 33324
rect 9577 33290 9611 33324
rect 9645 33290 9679 33324
rect 9713 33290 9747 33324
rect 9781 33290 9815 33324
rect 9849 33290 9883 33324
rect 9917 33290 9951 33324
rect 9985 33290 10019 33324
rect 10053 33290 10087 33324
rect 10121 33290 10155 33324
rect 10189 33290 10223 33324
rect 10257 33290 10291 33324
rect 10325 33290 10359 33324
rect 10393 33290 10427 33324
rect 10461 33290 10495 33324
rect 10529 33290 10563 33324
rect 10597 33290 10631 33324
rect 10665 33290 10699 33324
rect 10733 33290 10767 33324
rect 10801 33290 10835 33324
rect 10869 33290 10903 33324
rect 10937 33290 10971 33324
rect 11005 33290 11039 33324
rect 11073 33290 11107 33324
rect 11141 33290 11175 33324
rect 11209 33290 11243 33324
rect 11277 33290 11311 33324
rect 11345 33290 11379 33324
rect 11413 33290 11447 33324
rect 11481 33290 11515 33324
rect 11549 33290 11583 33324
rect 11617 33290 11651 33324
rect 11685 33290 11719 33324
rect 11753 33290 11787 33324
rect 11821 33290 11855 33324
rect 11889 33290 11923 33324
rect 11957 33290 11991 33324
rect 12025 33290 12059 33324
rect 12093 33290 12127 33324
rect 12161 33290 12195 33324
rect 12229 33290 12263 33324
rect 12297 33290 12331 33324
rect 12365 33290 12399 33324
rect 12433 33290 12467 33324
rect 12501 33290 12535 33324
rect 12569 33290 12603 33324
rect 12637 33290 12671 33324
rect 12705 33290 12739 33324
rect 12773 33290 12807 33324
rect 12841 33290 12875 33324
rect 12909 33290 12943 33324
rect 12977 33290 13118 33324
rect 2860 33288 13118 33290
rect 2673 33245 13118 33288
rect 2673 33211 2674 33245
rect 2708 33211 2750 33245
rect 2784 33211 2826 33245
rect 2860 33211 13118 33245
rect 2673 33168 13118 33211
rect 2673 33134 2674 33168
rect 2708 33134 2750 33168
rect 2784 33134 2826 33168
rect 2860 33134 13118 33168
rect 2673 33090 13118 33134
rect 2673 33056 2674 33090
rect 2708 33056 2750 33090
rect 2784 33056 2826 33090
rect 2860 33056 13118 33090
rect 2673 33012 13118 33056
rect 2673 32978 2674 33012
rect 2708 32978 2750 33012
rect 2784 32978 2826 33012
rect 2860 32978 13118 33012
rect 2673 32934 13118 32978
rect 2673 32900 2674 32934
rect 2708 32900 2750 32934
rect 2784 32900 2826 32934
rect 2860 32900 13118 32934
rect 2673 32856 13118 32900
rect 2673 32822 2674 32856
rect 2708 32822 2750 32856
rect 2784 32822 2826 32856
rect 2860 32854 13118 32856
rect 2860 32822 3507 32854
rect 2673 32820 3507 32822
rect 3541 32820 3576 32854
rect 3610 32820 3645 32854
rect 3679 32820 3714 32854
rect 3748 32820 3783 32854
rect 3817 32820 3852 32854
rect 3886 32820 3921 32854
rect 3955 32820 3990 32854
rect 4024 32820 4059 32854
rect 4093 32820 4128 32854
rect 4162 32820 4197 32854
rect 4231 32820 4266 32854
rect 4300 32820 4335 32854
rect 4369 32820 4404 32854
rect 4438 32820 4473 32854
rect 4507 32820 4542 32854
rect 4576 32820 4611 32854
rect 4645 32820 4680 32854
rect 4714 32820 4749 32854
rect 4783 32820 4818 32854
rect 4852 32820 4887 32854
rect 4921 32820 4956 32854
rect 4990 32820 5025 32854
rect 5059 32820 5094 32854
rect 5128 32820 5163 32854
rect 5197 32820 5232 32854
rect 5266 32820 5301 32854
rect 5335 32820 5370 32854
rect 5404 32820 5439 32854
rect 5473 32820 5508 32854
rect 5542 32820 5577 32854
rect 5611 32820 5646 32854
rect 5680 32820 5715 32854
rect 5749 32820 5784 32854
rect 5818 32820 5853 32854
rect 5887 32820 5922 32854
rect 5956 32820 5991 32854
rect 6025 32820 6060 32854
rect 6094 32820 6129 32854
rect 6163 32820 6198 32854
rect 6232 32820 6267 32854
rect 6301 32820 6336 32854
rect 6370 32820 6405 32854
rect 6439 32820 6474 32854
rect 6508 32820 6543 32854
rect 6577 32820 6612 32854
rect 6646 32820 6681 32854
rect 6715 32820 6750 32854
rect 6784 32820 6819 32854
rect 6853 32820 6888 32854
rect 6922 32820 6957 32854
rect 6991 32820 7026 32854
rect 7060 32820 7095 32854
rect 7129 32820 7163 32854
rect 7197 32820 7231 32854
rect 7265 32820 7299 32854
rect 7333 32820 7367 32854
rect 7401 32820 7435 32854
rect 7469 32820 7503 32854
rect 7537 32820 7571 32854
rect 7605 32820 7639 32854
rect 7673 32820 7707 32854
rect 7741 32820 7775 32854
rect 7809 32820 7843 32854
rect 7877 32820 7911 32854
rect 7945 32820 7979 32854
rect 8013 32820 8047 32854
rect 8081 32820 8115 32854
rect 8149 32820 8183 32854
rect 8217 32820 8251 32854
rect 8285 32820 8319 32854
rect 8353 32820 8387 32854
rect 8421 32820 8455 32854
rect 8489 32820 8523 32854
rect 8557 32820 8591 32854
rect 8625 32820 8659 32854
rect 8693 32820 8727 32854
rect 8761 32820 8795 32854
rect 8829 32820 8863 32854
rect 8897 32820 8931 32854
rect 8965 32820 8999 32854
rect 9033 32820 9067 32854
rect 9101 32820 9135 32854
rect 9169 32820 9203 32854
rect 9237 32820 9271 32854
rect 9305 32820 9339 32854
rect 9373 32820 9407 32854
rect 9441 32820 9475 32854
rect 9509 32820 9543 32854
rect 9577 32820 9611 32854
rect 9645 32820 9679 32854
rect 9713 32820 9747 32854
rect 9781 32820 9815 32854
rect 9849 32820 9883 32854
rect 9917 32820 9951 32854
rect 9985 32820 10019 32854
rect 10053 32820 10087 32854
rect 10121 32820 10155 32854
rect 10189 32820 10223 32854
rect 10257 32820 10291 32854
rect 10325 32820 10359 32854
rect 10393 32820 10427 32854
rect 10461 32820 10495 32854
rect 10529 32820 10563 32854
rect 10597 32820 10631 32854
rect 10665 32820 10699 32854
rect 10733 32820 10767 32854
rect 10801 32820 10835 32854
rect 10869 32820 10903 32854
rect 10937 32820 10971 32854
rect 11005 32820 11039 32854
rect 11073 32820 11107 32854
rect 11141 32820 11175 32854
rect 11209 32820 11243 32854
rect 11277 32820 11311 32854
rect 11345 32820 11379 32854
rect 11413 32820 11447 32854
rect 11481 32820 11515 32854
rect 11549 32820 11583 32854
rect 11617 32820 11651 32854
rect 11685 32820 11719 32854
rect 11753 32820 11787 32854
rect 11821 32820 11855 32854
rect 11889 32820 11923 32854
rect 11957 32820 11991 32854
rect 12025 32820 12059 32854
rect 12093 32820 12127 32854
rect 12161 32820 12195 32854
rect 12229 32820 12263 32854
rect 12297 32820 12331 32854
rect 12365 32820 12399 32854
rect 12433 32820 12467 32854
rect 12501 32820 12535 32854
rect 12569 32820 12603 32854
rect 12637 32820 12671 32854
rect 12705 32820 12739 32854
rect 12773 32820 12807 32854
rect 12841 32820 12875 32854
rect 12909 32820 12943 32854
rect 12977 32820 13118 32854
rect 2219 32768 2274 32807
rect 2253 32734 2274 32768
rect 2219 32695 2274 32734
rect 3593 32714 3695 32726
rect 4429 32714 4531 32726
rect 5265 32714 5367 32726
rect 6101 32714 6203 32726
rect 6937 32714 7039 32726
rect 7773 32714 7875 32726
rect 8609 32714 8711 32726
rect 9445 32714 9547 32726
rect 10281 32714 10383 32726
rect 11117 32714 11219 32726
rect 11953 32714 12055 32726
rect 12789 32714 12891 32726
rect 2253 32661 2274 32695
rect 2219 32622 2274 32661
rect 2253 32588 2274 32622
rect 2219 32549 2274 32588
rect 2253 32515 2274 32549
rect 2219 32476 2274 32515
rect 2253 32442 2274 32476
rect 2219 32403 2274 32442
rect 2253 32369 2274 32403
rect 2219 32330 2274 32369
rect 2253 32296 2274 32330
rect 2219 32257 2274 32296
rect 2253 32223 2274 32257
rect 2219 32184 2274 32223
rect 2253 32150 2274 32184
rect 2219 32111 2274 32150
rect 2253 32077 2274 32111
rect 2219 32038 2274 32077
rect 2253 32004 2274 32038
rect 2219 31965 2274 32004
rect 2253 31931 2274 31965
rect 2219 31892 2274 31931
rect 2253 31858 2274 31892
rect 2219 31819 2274 31858
rect 2253 31785 2274 31819
rect 2219 31746 2274 31785
rect 2253 31712 2274 31746
rect 2219 31673 2274 31712
rect 2253 31639 2274 31673
rect 2219 31600 2274 31639
rect 2253 31566 2274 31600
rect 2219 31527 2274 31566
rect 2253 31493 2274 31527
rect 2219 31454 2274 31493
rect 2253 31420 2274 31454
rect 2219 31381 2274 31420
rect 2253 31347 2274 31381
rect 3207 32680 3245 32714
rect 3173 32641 3279 32680
rect 3207 32607 3245 32641
rect 3173 32568 3279 32607
rect 3207 32534 3245 32568
rect 3173 32495 3279 32534
rect 3207 32461 3245 32495
rect 3173 32422 3279 32461
rect 3625 32680 3663 32714
rect 3591 32641 3697 32680
rect 3625 32607 3663 32641
rect 3591 32568 3697 32607
rect 3625 32534 3663 32568
rect 3591 32495 3697 32534
rect 3625 32461 3663 32495
rect 3591 32422 3697 32461
rect 4043 32680 4081 32714
rect 4009 32641 4115 32680
rect 4043 32607 4081 32641
rect 4009 32568 4115 32607
rect 4043 32534 4081 32568
rect 4009 32495 4115 32534
rect 4043 32461 4081 32495
rect 4009 32422 4115 32461
rect 4461 32680 4499 32714
rect 4427 32641 4533 32680
rect 4461 32607 4499 32641
rect 4427 32568 4533 32607
rect 4461 32534 4499 32568
rect 4427 32495 4533 32534
rect 4461 32461 4499 32495
rect 4427 32422 4533 32461
rect 4879 32680 4917 32714
rect 4845 32641 4951 32680
rect 4879 32607 4917 32641
rect 4845 32568 4951 32607
rect 4879 32534 4917 32568
rect 4845 32495 4951 32534
rect 4879 32461 4917 32495
rect 4845 32422 4951 32461
rect 5297 32680 5335 32714
rect 5263 32641 5369 32680
rect 5297 32607 5335 32641
rect 5263 32568 5369 32607
rect 5297 32534 5335 32568
rect 5263 32495 5369 32534
rect 5297 32461 5335 32495
rect 5263 32422 5369 32461
rect 5715 32680 5753 32714
rect 5681 32641 5787 32680
rect 5715 32607 5753 32641
rect 5681 32568 5787 32607
rect 5715 32534 5753 32568
rect 5681 32495 5787 32534
rect 5715 32461 5753 32495
rect 5681 32422 5787 32461
rect 6133 32680 6171 32714
rect 6099 32641 6205 32680
rect 6133 32607 6171 32641
rect 6099 32568 6205 32607
rect 6133 32534 6171 32568
rect 6099 32495 6205 32534
rect 6133 32461 6171 32495
rect 6099 32422 6205 32461
rect 6551 32680 6589 32714
rect 6517 32641 6623 32680
rect 6551 32607 6589 32641
rect 6517 32568 6623 32607
rect 6551 32534 6589 32568
rect 6517 32495 6623 32534
rect 6551 32461 6589 32495
rect 6517 32422 6623 32461
rect 6969 32680 7007 32714
rect 6935 32641 7041 32680
rect 6969 32607 7007 32641
rect 6935 32568 7041 32607
rect 6969 32534 7007 32568
rect 6935 32495 7041 32534
rect 6969 32461 7007 32495
rect 6935 32422 7041 32461
rect 7387 32680 7425 32714
rect 7353 32641 7459 32680
rect 7387 32607 7425 32641
rect 7353 32568 7459 32607
rect 7387 32534 7425 32568
rect 7353 32495 7459 32534
rect 7387 32461 7425 32495
rect 7353 32422 7459 32461
rect 7805 32680 7843 32714
rect 7771 32641 7877 32680
rect 7805 32607 7843 32641
rect 7771 32568 7877 32607
rect 7805 32534 7843 32568
rect 7771 32495 7877 32534
rect 7805 32461 7843 32495
rect 7771 32422 7877 32461
rect 8223 32680 8261 32714
rect 8189 32641 8295 32680
rect 8223 32607 8261 32641
rect 8189 32568 8295 32607
rect 8223 32534 8261 32568
rect 8189 32495 8295 32534
rect 8223 32461 8261 32495
rect 8189 32422 8295 32461
rect 8641 32680 8679 32714
rect 8607 32641 8713 32680
rect 8641 32607 8679 32641
rect 8607 32568 8713 32607
rect 8641 32534 8679 32568
rect 8607 32495 8713 32534
rect 8641 32461 8679 32495
rect 8607 32422 8713 32461
rect 9059 32680 9097 32714
rect 9025 32641 9131 32680
rect 9059 32607 9097 32641
rect 9025 32568 9131 32607
rect 9059 32534 9097 32568
rect 9025 32495 9131 32534
rect 9059 32461 9097 32495
rect 9025 32422 9131 32461
rect 9477 32680 9515 32714
rect 9443 32641 9549 32680
rect 9477 32607 9515 32641
rect 9443 32568 9549 32607
rect 9477 32534 9515 32568
rect 9443 32495 9549 32534
rect 9477 32461 9515 32495
rect 9443 32422 9549 32461
rect 9895 32680 9933 32714
rect 9861 32641 9967 32680
rect 9895 32607 9933 32641
rect 9861 32568 9967 32607
rect 9895 32534 9933 32568
rect 9861 32495 9967 32534
rect 9895 32461 9933 32495
rect 9861 32422 9967 32461
rect 10313 32680 10351 32714
rect 10279 32641 10385 32680
rect 10313 32607 10351 32641
rect 10279 32568 10385 32607
rect 10313 32534 10351 32568
rect 10279 32495 10385 32534
rect 10313 32461 10351 32495
rect 10279 32422 10385 32461
rect 10731 32680 10769 32714
rect 10697 32641 10803 32680
rect 10731 32607 10769 32641
rect 10697 32568 10803 32607
rect 10731 32534 10769 32568
rect 10697 32495 10803 32534
rect 10731 32461 10769 32495
rect 10697 32422 10803 32461
rect 11149 32680 11187 32714
rect 11115 32641 11221 32680
rect 11149 32607 11187 32641
rect 11115 32568 11221 32607
rect 11149 32534 11187 32568
rect 11115 32495 11221 32534
rect 11149 32461 11187 32495
rect 11115 32422 11221 32461
rect 11567 32680 11605 32714
rect 11533 32641 11639 32680
rect 11567 32607 11605 32641
rect 11533 32568 11639 32607
rect 11567 32534 11605 32568
rect 11533 32495 11639 32534
rect 11567 32461 11605 32495
rect 11533 32422 11639 32461
rect 11985 32680 12023 32714
rect 11951 32641 12057 32680
rect 11985 32607 12023 32641
rect 11951 32568 12057 32607
rect 11985 32534 12023 32568
rect 11951 32495 12057 32534
rect 11985 32461 12023 32495
rect 11951 32422 12057 32461
rect 12403 32680 12441 32714
rect 12369 32641 12475 32680
rect 12403 32607 12441 32641
rect 12369 32568 12475 32607
rect 12403 32534 12441 32568
rect 12369 32495 12475 32534
rect 12403 32461 12441 32495
rect 12369 32422 12475 32461
rect 12821 32680 12859 32714
rect 12787 32641 12893 32680
rect 12821 32607 12859 32641
rect 12787 32568 12893 32607
rect 12821 32534 12859 32568
rect 12787 32495 12893 32534
rect 12821 32461 12859 32495
rect 12787 32422 12893 32461
rect 13239 32680 13277 32714
rect 13205 32641 13311 32680
rect 13239 32607 13277 32641
rect 13205 32568 13311 32607
rect 13239 32534 13277 32568
rect 13205 32495 13311 32534
rect 13239 32461 13277 32495
rect 13205 32422 13311 32461
rect 3593 31368 3695 31380
rect 4429 31368 4531 31380
rect 5265 31368 5367 31380
rect 6101 31368 6203 31380
rect 6937 31368 7039 31380
rect 7773 31368 7875 31380
rect 8609 31368 8711 31380
rect 9445 31368 9547 31380
rect 10281 31368 10383 31380
rect 11117 31368 11219 31380
rect 11953 31368 12055 31380
rect 12789 31368 12891 31380
rect 2219 31308 2274 31347
rect 2253 31274 2274 31308
rect 2219 31235 2274 31274
rect 2253 31201 2274 31235
rect 2219 31162 2274 31201
rect 2253 31128 2274 31162
rect 2219 31089 2274 31128
rect 2253 31055 2274 31089
rect 2219 31016 2274 31055
rect 2253 30982 2274 31016
rect 2219 30943 2274 30982
rect 2253 30909 2274 30943
rect 2219 30871 2274 30909
rect 2253 30837 2274 30871
rect 2219 30799 2274 30837
rect 2673 31323 3507 31324
rect 2673 31289 2674 31323
rect 2708 31289 2750 31323
rect 2784 31289 2826 31323
rect 2860 31290 3507 31323
rect 3541 31290 3576 31324
rect 3610 31290 3645 31324
rect 3679 31290 3714 31324
rect 3748 31290 3783 31324
rect 3817 31290 3852 31324
rect 3886 31290 3921 31324
rect 3955 31290 3990 31324
rect 4024 31290 4059 31324
rect 4093 31290 4128 31324
rect 4162 31290 4197 31324
rect 4231 31290 4266 31324
rect 4300 31290 4335 31324
rect 4369 31290 4404 31324
rect 4438 31290 4473 31324
rect 4507 31290 4542 31324
rect 4576 31290 4611 31324
rect 4645 31290 4680 31324
rect 4714 31290 4749 31324
rect 4783 31290 4818 31324
rect 4852 31290 4887 31324
rect 4921 31290 4956 31324
rect 4990 31290 5025 31324
rect 5059 31290 5094 31324
rect 5128 31290 5163 31324
rect 5197 31290 5232 31324
rect 5266 31290 5301 31324
rect 5335 31290 5370 31324
rect 5404 31290 5439 31324
rect 5473 31290 5508 31324
rect 5542 31290 5577 31324
rect 5611 31290 5646 31324
rect 5680 31290 5715 31324
rect 5749 31290 5784 31324
rect 5818 31290 5853 31324
rect 5887 31290 5922 31324
rect 5956 31290 5991 31324
rect 6025 31290 6060 31324
rect 6094 31290 6129 31324
rect 6163 31290 6198 31324
rect 6232 31290 6267 31324
rect 6301 31290 6336 31324
rect 6370 31290 6405 31324
rect 6439 31290 6474 31324
rect 6508 31290 6543 31324
rect 6577 31290 6612 31324
rect 6646 31290 6681 31324
rect 6715 31290 6750 31324
rect 6784 31290 6819 31324
rect 6853 31290 6888 31324
rect 6922 31290 6957 31324
rect 6991 31290 7026 31324
rect 7060 31290 7095 31324
rect 7129 31290 7163 31324
rect 7197 31290 7231 31324
rect 7265 31290 7299 31324
rect 7333 31290 7367 31324
rect 7401 31290 7435 31324
rect 7469 31290 7503 31324
rect 7537 31290 7571 31324
rect 7605 31290 7639 31324
rect 7673 31290 7707 31324
rect 7741 31290 7775 31324
rect 7809 31290 7843 31324
rect 7877 31290 7911 31324
rect 7945 31290 7979 31324
rect 8013 31290 8047 31324
rect 8081 31290 8115 31324
rect 8149 31290 8183 31324
rect 8217 31290 8251 31324
rect 8285 31290 8319 31324
rect 8353 31290 8387 31324
rect 8421 31290 8455 31324
rect 8489 31290 8523 31324
rect 8557 31290 8591 31324
rect 8625 31290 8659 31324
rect 8693 31290 8727 31324
rect 8761 31290 8795 31324
rect 8829 31290 8863 31324
rect 8897 31290 8931 31324
rect 8965 31290 8999 31324
rect 9033 31290 9067 31324
rect 9101 31290 9135 31324
rect 9169 31290 9203 31324
rect 9237 31290 9271 31324
rect 9305 31290 9339 31324
rect 9373 31290 9407 31324
rect 9441 31290 9475 31324
rect 9509 31290 9543 31324
rect 9577 31290 9611 31324
rect 9645 31290 9679 31324
rect 9713 31290 9747 31324
rect 9781 31290 9815 31324
rect 9849 31290 9883 31324
rect 9917 31290 9951 31324
rect 9985 31290 10019 31324
rect 10053 31290 10087 31324
rect 10121 31290 10155 31324
rect 10189 31290 10223 31324
rect 10257 31290 10291 31324
rect 10325 31290 10359 31324
rect 10393 31290 10427 31324
rect 10461 31290 10495 31324
rect 10529 31290 10563 31324
rect 10597 31290 10631 31324
rect 10665 31290 10699 31324
rect 10733 31290 10767 31324
rect 10801 31290 10835 31324
rect 10869 31290 10903 31324
rect 10937 31290 10971 31324
rect 11005 31290 11039 31324
rect 11073 31290 11107 31324
rect 11141 31290 11175 31324
rect 11209 31290 11243 31324
rect 11277 31290 11311 31324
rect 11345 31290 11379 31324
rect 11413 31290 11447 31324
rect 11481 31290 11515 31324
rect 11549 31290 11583 31324
rect 11617 31290 11651 31324
rect 11685 31290 11719 31324
rect 11753 31290 11787 31324
rect 11821 31290 11855 31324
rect 11889 31290 11923 31324
rect 11957 31290 11991 31324
rect 12025 31290 12059 31324
rect 12093 31290 12127 31324
rect 12161 31290 12195 31324
rect 12229 31290 12263 31324
rect 12297 31290 12331 31324
rect 12365 31290 12399 31324
rect 12433 31290 12467 31324
rect 12501 31290 12535 31324
rect 12569 31290 12603 31324
rect 12637 31290 12671 31324
rect 12705 31290 12739 31324
rect 12773 31290 12807 31324
rect 12841 31290 12875 31324
rect 12909 31290 12943 31324
rect 12977 31290 13118 31324
rect 2860 31289 13118 31290
rect 2673 31246 13118 31289
rect 2673 31212 2674 31246
rect 2708 31212 2750 31246
rect 2784 31212 2826 31246
rect 2860 31212 13118 31246
rect 2673 31169 13118 31212
rect 2673 31135 2674 31169
rect 2708 31135 2750 31169
rect 2784 31135 2826 31169
rect 2860 31135 13118 31169
rect 2673 31091 13118 31135
rect 2673 31057 2674 31091
rect 2708 31057 2750 31091
rect 2784 31057 2826 31091
rect 2860 31057 13118 31091
rect 2673 31013 13118 31057
rect 2673 30979 2674 31013
rect 2708 30979 2750 31013
rect 2784 30979 2826 31013
rect 2860 30979 13118 31013
rect 2673 30935 13118 30979
rect 2673 30901 2674 30935
rect 2708 30901 2750 30935
rect 2784 30901 2826 30935
rect 2860 30901 13118 30935
rect 2673 30857 13118 30901
rect 2673 30823 2674 30857
rect 2708 30823 2750 30857
rect 2784 30823 2826 30857
rect 2860 30854 13118 30857
rect 2860 30823 3507 30854
rect 2673 30820 3507 30823
rect 3541 30820 3576 30854
rect 3610 30820 3645 30854
rect 3679 30820 3714 30854
rect 3748 30820 3783 30854
rect 3817 30820 3852 30854
rect 3886 30820 3921 30854
rect 3955 30820 3990 30854
rect 4024 30820 4059 30854
rect 4093 30820 4128 30854
rect 4162 30820 4197 30854
rect 4231 30820 4266 30854
rect 4300 30820 4335 30854
rect 4369 30820 4404 30854
rect 4438 30820 4473 30854
rect 4507 30820 4542 30854
rect 4576 30820 4611 30854
rect 4645 30820 4680 30854
rect 4714 30820 4749 30854
rect 4783 30820 4818 30854
rect 4852 30820 4887 30854
rect 4921 30820 4956 30854
rect 4990 30820 5025 30854
rect 5059 30820 5094 30854
rect 5128 30820 5163 30854
rect 5197 30820 5232 30854
rect 5266 30820 5301 30854
rect 5335 30820 5370 30854
rect 5404 30820 5439 30854
rect 5473 30820 5508 30854
rect 5542 30820 5577 30854
rect 5611 30820 5646 30854
rect 5680 30820 5715 30854
rect 5749 30820 5784 30854
rect 5818 30820 5853 30854
rect 5887 30820 5922 30854
rect 5956 30820 5991 30854
rect 6025 30820 6060 30854
rect 6094 30820 6129 30854
rect 6163 30820 6198 30854
rect 6232 30820 6267 30854
rect 6301 30820 6336 30854
rect 6370 30820 6405 30854
rect 6439 30820 6474 30854
rect 6508 30820 6543 30854
rect 6577 30820 6612 30854
rect 6646 30820 6681 30854
rect 6715 30820 6750 30854
rect 6784 30820 6819 30854
rect 6853 30820 6888 30854
rect 6922 30820 6957 30854
rect 6991 30820 7026 30854
rect 7060 30820 7095 30854
rect 7129 30820 7163 30854
rect 7197 30820 7231 30854
rect 7265 30820 7299 30854
rect 7333 30820 7367 30854
rect 7401 30820 7435 30854
rect 7469 30820 7503 30854
rect 7537 30820 7571 30854
rect 7605 30820 7639 30854
rect 7673 30820 7707 30854
rect 7741 30820 7775 30854
rect 7809 30820 7843 30854
rect 7877 30820 7911 30854
rect 7945 30820 7979 30854
rect 8013 30820 8047 30854
rect 8081 30820 8115 30854
rect 8149 30820 8183 30854
rect 8217 30820 8251 30854
rect 8285 30820 8319 30854
rect 8353 30820 8387 30854
rect 8421 30820 8455 30854
rect 8489 30820 8523 30854
rect 8557 30820 8591 30854
rect 8625 30820 8659 30854
rect 8693 30820 8727 30854
rect 8761 30820 8795 30854
rect 8829 30820 8863 30854
rect 8897 30820 8931 30854
rect 8965 30820 8999 30854
rect 9033 30820 9067 30854
rect 9101 30820 9135 30854
rect 9169 30820 9203 30854
rect 9237 30820 9271 30854
rect 9305 30820 9339 30854
rect 9373 30820 9407 30854
rect 9441 30820 9475 30854
rect 9509 30820 9543 30854
rect 9577 30820 9611 30854
rect 9645 30820 9679 30854
rect 9713 30820 9747 30854
rect 9781 30820 9815 30854
rect 9849 30820 9883 30854
rect 9917 30820 9951 30854
rect 9985 30820 10019 30854
rect 10053 30820 10087 30854
rect 10121 30820 10155 30854
rect 10189 30820 10223 30854
rect 10257 30820 10291 30854
rect 10325 30820 10359 30854
rect 10393 30820 10427 30854
rect 10461 30820 10495 30854
rect 10529 30820 10563 30854
rect 10597 30820 10631 30854
rect 10665 30820 10699 30854
rect 10733 30820 10767 30854
rect 10801 30820 10835 30854
rect 10869 30820 10903 30854
rect 10937 30820 10971 30854
rect 11005 30820 11039 30854
rect 11073 30820 11107 30854
rect 11141 30820 11175 30854
rect 11209 30820 11243 30854
rect 11277 30820 11311 30854
rect 11345 30820 11379 30854
rect 11413 30820 11447 30854
rect 11481 30820 11515 30854
rect 11549 30820 11583 30854
rect 11617 30820 11651 30854
rect 11685 30820 11719 30854
rect 11753 30820 11787 30854
rect 11821 30820 11855 30854
rect 11889 30820 11923 30854
rect 11957 30820 11991 30854
rect 12025 30820 12059 30854
rect 12093 30820 12127 30854
rect 12161 30820 12195 30854
rect 12229 30820 12263 30854
rect 12297 30820 12331 30854
rect 12365 30820 12399 30854
rect 12433 30820 12467 30854
rect 12501 30820 12535 30854
rect 12569 30820 12603 30854
rect 12637 30820 12671 30854
rect 12705 30820 12739 30854
rect 12773 30820 12807 30854
rect 12841 30820 12875 30854
rect 12909 30820 12943 30854
rect 12977 30820 13118 30854
rect 2253 30765 2274 30799
rect 2219 30727 2274 30765
rect 2253 30693 2274 30727
rect 3593 30714 3695 30726
rect 4429 30714 4531 30726
rect 5265 30714 5367 30726
rect 6101 30714 6203 30726
rect 6937 30714 7039 30726
rect 7773 30714 7875 30726
rect 8609 30714 8711 30726
rect 9445 30714 9547 30726
rect 10281 30714 10383 30726
rect 11117 30714 11219 30726
rect 11953 30714 12055 30726
rect 12789 30714 12891 30726
rect 2219 30655 2274 30693
rect 2253 30621 2274 30655
rect 2219 30583 2274 30621
rect 2253 30549 2274 30583
rect 2219 30511 2274 30549
rect 2253 30477 2274 30511
rect 2219 30439 2274 30477
rect 2253 30405 2274 30439
rect 2219 30367 2274 30405
rect 2253 30333 2274 30367
rect 2219 30295 2274 30333
rect 2253 30261 2274 30295
rect 2219 30223 2274 30261
rect 2253 30189 2274 30223
rect 2219 30151 2274 30189
rect 2253 30117 2274 30151
rect 2219 30079 2274 30117
rect 2253 30045 2274 30079
rect 2219 30007 2274 30045
rect 2253 29973 2274 30007
rect 2219 29935 2274 29973
rect 2253 29901 2274 29935
rect 2219 29863 2274 29901
rect 2253 29829 2274 29863
rect 2219 29791 2274 29829
rect 2253 29757 2274 29791
rect 2219 29719 2274 29757
rect 2253 29685 2274 29719
rect 2219 29647 2274 29685
rect 2253 29613 2274 29647
rect 2219 29575 2274 29613
rect 2253 29541 2274 29575
rect 2219 29503 2274 29541
rect 2253 29469 2274 29503
rect 2219 29431 2274 29469
rect 2253 29397 2274 29431
rect 2219 29359 2274 29397
rect 3207 30680 3245 30714
rect 3173 30641 3279 30680
rect 3207 30607 3245 30641
rect 3173 30568 3279 30607
rect 3207 30534 3245 30568
rect 3173 30495 3279 30534
rect 3207 30461 3245 30495
rect 3173 30422 3279 30461
rect 3625 30680 3663 30714
rect 3591 30641 3697 30680
rect 3625 30607 3663 30641
rect 3591 30568 3697 30607
rect 3625 30534 3663 30568
rect 3591 30495 3697 30534
rect 3625 30461 3663 30495
rect 3591 30422 3697 30461
rect 4043 30680 4081 30714
rect 4009 30641 4115 30680
rect 4043 30607 4081 30641
rect 4009 30568 4115 30607
rect 4043 30534 4081 30568
rect 4009 30495 4115 30534
rect 4043 30461 4081 30495
rect 4009 30422 4115 30461
rect 4461 30680 4499 30714
rect 4427 30641 4533 30680
rect 4461 30607 4499 30641
rect 4427 30568 4533 30607
rect 4461 30534 4499 30568
rect 4427 30495 4533 30534
rect 4461 30461 4499 30495
rect 4427 30422 4533 30461
rect 4879 30680 4917 30714
rect 4845 30641 4951 30680
rect 4879 30607 4917 30641
rect 4845 30568 4951 30607
rect 4879 30534 4917 30568
rect 4845 30495 4951 30534
rect 4879 30461 4917 30495
rect 4845 30422 4951 30461
rect 5297 30680 5335 30714
rect 5263 30641 5369 30680
rect 5297 30607 5335 30641
rect 5263 30568 5369 30607
rect 5297 30534 5335 30568
rect 5263 30495 5369 30534
rect 5297 30461 5335 30495
rect 5263 30422 5369 30461
rect 5715 30680 5753 30714
rect 5681 30641 5787 30680
rect 5715 30607 5753 30641
rect 5681 30568 5787 30607
rect 5715 30534 5753 30568
rect 5681 30495 5787 30534
rect 5715 30461 5753 30495
rect 5681 30422 5787 30461
rect 6133 30680 6171 30714
rect 6099 30641 6205 30680
rect 6133 30607 6171 30641
rect 6099 30568 6205 30607
rect 6133 30534 6171 30568
rect 6099 30495 6205 30534
rect 6133 30461 6171 30495
rect 6099 30422 6205 30461
rect 6551 30680 6589 30714
rect 6517 30641 6623 30680
rect 6551 30607 6589 30641
rect 6517 30568 6623 30607
rect 6551 30534 6589 30568
rect 6517 30495 6623 30534
rect 6551 30461 6589 30495
rect 6517 30422 6623 30461
rect 6969 30680 7007 30714
rect 6935 30641 7041 30680
rect 6969 30607 7007 30641
rect 6935 30568 7041 30607
rect 6969 30534 7007 30568
rect 6935 30495 7041 30534
rect 6969 30461 7007 30495
rect 6935 30422 7041 30461
rect 7387 30680 7425 30714
rect 7353 30641 7459 30680
rect 7387 30607 7425 30641
rect 7353 30568 7459 30607
rect 7387 30534 7425 30568
rect 7353 30495 7459 30534
rect 7387 30461 7425 30495
rect 7353 30422 7459 30461
rect 7805 30680 7843 30714
rect 7771 30641 7877 30680
rect 7805 30607 7843 30641
rect 7771 30568 7877 30607
rect 7805 30534 7843 30568
rect 7771 30495 7877 30534
rect 7805 30461 7843 30495
rect 7771 30422 7877 30461
rect 8223 30680 8261 30714
rect 8189 30641 8295 30680
rect 8223 30607 8261 30641
rect 8189 30568 8295 30607
rect 8223 30534 8261 30568
rect 8189 30495 8295 30534
rect 8223 30461 8261 30495
rect 8189 30422 8295 30461
rect 8641 30680 8679 30714
rect 8607 30641 8713 30680
rect 8641 30607 8679 30641
rect 8607 30568 8713 30607
rect 8641 30534 8679 30568
rect 8607 30495 8713 30534
rect 8641 30461 8679 30495
rect 8607 30422 8713 30461
rect 9059 30680 9097 30714
rect 9025 30641 9131 30680
rect 9059 30607 9097 30641
rect 9025 30568 9131 30607
rect 9059 30534 9097 30568
rect 9025 30495 9131 30534
rect 9059 30461 9097 30495
rect 9025 30422 9131 30461
rect 9477 30680 9515 30714
rect 9443 30641 9549 30680
rect 9477 30607 9515 30641
rect 9443 30568 9549 30607
rect 9477 30534 9515 30568
rect 9443 30495 9549 30534
rect 9477 30461 9515 30495
rect 9443 30422 9549 30461
rect 9895 30680 9933 30714
rect 9861 30641 9967 30680
rect 9895 30607 9933 30641
rect 9861 30568 9967 30607
rect 9895 30534 9933 30568
rect 9861 30495 9967 30534
rect 9895 30461 9933 30495
rect 9861 30422 9967 30461
rect 10313 30680 10351 30714
rect 10279 30641 10385 30680
rect 10313 30607 10351 30641
rect 10279 30568 10385 30607
rect 10313 30534 10351 30568
rect 10279 30495 10385 30534
rect 10313 30461 10351 30495
rect 10279 30422 10385 30461
rect 10731 30680 10769 30714
rect 10697 30641 10803 30680
rect 10731 30607 10769 30641
rect 10697 30568 10803 30607
rect 10731 30534 10769 30568
rect 10697 30495 10803 30534
rect 10731 30461 10769 30495
rect 10697 30422 10803 30461
rect 11149 30680 11187 30714
rect 11115 30641 11221 30680
rect 11149 30607 11187 30641
rect 11115 30568 11221 30607
rect 11149 30534 11187 30568
rect 11115 30495 11221 30534
rect 11149 30461 11187 30495
rect 11115 30422 11221 30461
rect 11567 30680 11605 30714
rect 11533 30641 11639 30680
rect 11567 30607 11605 30641
rect 11533 30568 11639 30607
rect 11567 30534 11605 30568
rect 11533 30495 11639 30534
rect 11567 30461 11605 30495
rect 11533 30422 11639 30461
rect 11985 30680 12023 30714
rect 11951 30641 12057 30680
rect 11985 30607 12023 30641
rect 11951 30568 12057 30607
rect 11985 30534 12023 30568
rect 11951 30495 12057 30534
rect 11985 30461 12023 30495
rect 11951 30422 12057 30461
rect 12403 30680 12441 30714
rect 12369 30641 12475 30680
rect 12403 30607 12441 30641
rect 12369 30568 12475 30607
rect 12403 30534 12441 30568
rect 12369 30495 12475 30534
rect 12403 30461 12441 30495
rect 12369 30422 12475 30461
rect 12821 30680 12859 30714
rect 12787 30641 12893 30680
rect 12821 30607 12859 30641
rect 12787 30568 12893 30607
rect 12821 30534 12859 30568
rect 12787 30495 12893 30534
rect 12821 30461 12859 30495
rect 12787 30422 12893 30461
rect 13239 30680 13277 30714
rect 13205 30641 13311 30680
rect 13239 30607 13277 30641
rect 13205 30568 13311 30607
rect 13239 30534 13277 30568
rect 13205 30495 13311 30534
rect 13239 30461 13277 30495
rect 13205 30422 13311 30461
rect 3593 29368 3695 29380
rect 4429 29368 4531 29380
rect 5265 29368 5367 29380
rect 6101 29368 6203 29380
rect 6937 29368 7039 29380
rect 7773 29368 7875 29380
rect 8609 29368 8711 29380
rect 9445 29368 9547 29380
rect 10281 29368 10383 29380
rect 11117 29368 11219 29380
rect 11953 29368 12055 29380
rect 12789 29368 12891 29380
rect 2253 29325 2274 29359
rect 2219 29287 2274 29325
rect 2253 29253 2274 29287
rect 2219 29215 2274 29253
rect 2253 29181 2274 29215
rect 2219 29143 2274 29181
rect 2253 29109 2274 29143
rect 2219 29089 2274 29109
rect 2376 29089 2444 29157
rect 2673 29320 3507 29324
rect 2673 29286 2674 29320
rect 2708 29286 2750 29320
rect 2784 29286 2826 29320
rect 2860 29290 3507 29320
rect 3541 29290 3576 29324
rect 3610 29290 3645 29324
rect 3679 29290 3714 29324
rect 3748 29290 3783 29324
rect 3817 29290 3852 29324
rect 3886 29290 3921 29324
rect 3955 29290 3990 29324
rect 4024 29290 4059 29324
rect 4093 29290 4128 29324
rect 4162 29290 4197 29324
rect 4231 29290 4266 29324
rect 4300 29290 4335 29324
rect 4369 29290 4404 29324
rect 4438 29290 4473 29324
rect 4507 29290 4542 29324
rect 4576 29290 4611 29324
rect 4645 29290 4680 29324
rect 4714 29290 4749 29324
rect 4783 29290 4818 29324
rect 4852 29290 4887 29324
rect 4921 29290 4956 29324
rect 4990 29290 5025 29324
rect 5059 29290 5094 29324
rect 5128 29290 5163 29324
rect 5197 29290 5232 29324
rect 5266 29290 5301 29324
rect 5335 29290 5370 29324
rect 5404 29290 5439 29324
rect 5473 29290 5508 29324
rect 5542 29290 5577 29324
rect 5611 29290 5646 29324
rect 5680 29290 5715 29324
rect 5749 29290 5784 29324
rect 5818 29290 5853 29324
rect 5887 29290 5922 29324
rect 5956 29290 5991 29324
rect 6025 29290 6060 29324
rect 6094 29290 6129 29324
rect 6163 29290 6198 29324
rect 6232 29290 6267 29324
rect 6301 29290 6336 29324
rect 6370 29290 6405 29324
rect 6439 29290 6474 29324
rect 6508 29290 6543 29324
rect 6577 29290 6612 29324
rect 6646 29290 6681 29324
rect 6715 29290 6750 29324
rect 6784 29290 6819 29324
rect 6853 29290 6888 29324
rect 6922 29290 6957 29324
rect 6991 29290 7026 29324
rect 7060 29290 7095 29324
rect 7129 29290 7163 29324
rect 7197 29290 7231 29324
rect 7265 29290 7299 29324
rect 7333 29290 7367 29324
rect 7401 29290 7435 29324
rect 7469 29290 7503 29324
rect 7537 29290 7571 29324
rect 7605 29290 7639 29324
rect 7673 29290 7707 29324
rect 7741 29290 7775 29324
rect 7809 29290 7843 29324
rect 7877 29290 7911 29324
rect 7945 29290 7979 29324
rect 8013 29290 8047 29324
rect 8081 29290 8115 29324
rect 8149 29290 8183 29324
rect 8217 29290 8251 29324
rect 8285 29290 8319 29324
rect 8353 29290 8387 29324
rect 8421 29290 8455 29324
rect 8489 29290 8523 29324
rect 8557 29290 8591 29324
rect 8625 29290 8659 29324
rect 8693 29290 8727 29324
rect 8761 29290 8795 29324
rect 8829 29290 8863 29324
rect 8897 29290 8931 29324
rect 8965 29290 8999 29324
rect 9033 29290 9067 29324
rect 9101 29290 9135 29324
rect 9169 29290 9203 29324
rect 9237 29290 9271 29324
rect 9305 29290 9339 29324
rect 9373 29290 9407 29324
rect 9441 29290 9475 29324
rect 9509 29290 9543 29324
rect 9577 29290 9611 29324
rect 9645 29290 9679 29324
rect 9713 29290 9747 29324
rect 9781 29290 9815 29324
rect 9849 29290 9883 29324
rect 9917 29290 9951 29324
rect 9985 29290 10019 29324
rect 10053 29290 10087 29324
rect 10121 29290 10155 29324
rect 10189 29290 10223 29324
rect 10257 29290 10291 29324
rect 10325 29290 10359 29324
rect 10393 29290 10427 29324
rect 10461 29290 10495 29324
rect 10529 29290 10563 29324
rect 10597 29290 10631 29324
rect 10665 29290 10699 29324
rect 10733 29290 10767 29324
rect 10801 29290 10835 29324
rect 10869 29290 10903 29324
rect 10937 29290 10971 29324
rect 11005 29290 11039 29324
rect 11073 29290 11107 29324
rect 11141 29290 11175 29324
rect 11209 29290 11243 29324
rect 11277 29290 11311 29324
rect 11345 29290 11379 29324
rect 11413 29290 11447 29324
rect 11481 29290 11515 29324
rect 11549 29290 11583 29324
rect 11617 29290 11651 29324
rect 11685 29290 11719 29324
rect 11753 29290 11787 29324
rect 11821 29290 11855 29324
rect 11889 29290 11923 29324
rect 11957 29290 11991 29324
rect 12025 29290 12059 29324
rect 12093 29290 12127 29324
rect 12161 29290 12195 29324
rect 12229 29290 12263 29324
rect 12297 29290 12331 29324
rect 12365 29290 12399 29324
rect 12433 29290 12467 29324
rect 12501 29290 12535 29324
rect 12569 29290 12603 29324
rect 12637 29290 12671 29324
rect 12705 29290 12739 29324
rect 12773 29290 12807 29324
rect 12841 29290 12875 29324
rect 12909 29290 12943 29324
rect 12977 29290 13118 29324
rect 2860 29286 13118 29290
rect 2673 29239 13118 29286
rect 2673 29205 2674 29239
rect 2708 29205 2750 29239
rect 2784 29205 2826 29239
rect 2860 29205 13118 29239
rect 2673 29157 13118 29205
rect 2673 29123 2674 29157
rect 2708 29123 2750 29157
rect 2784 29123 2826 29157
rect 2860 29124 13118 29157
rect 2860 29123 2861 29124
rect 2219 29071 2444 29089
rect 2253 29055 2325 29071
rect 2253 29037 2274 29055
rect 2219 29021 2274 29037
rect 2308 29037 2325 29055
rect 2359 29063 2444 29071
rect 2359 29037 2410 29063
rect 2308 29021 2410 29037
rect 2219 28999 2410 29021
rect 2253 28965 2325 28999
rect 2359 28995 2410 28999
rect 4144 29029 4178 29063
rect 4212 29029 4298 29063
rect 4144 28995 4298 29029
rect 2219 28927 2342 28965
rect 4144 28961 4196 28995
rect 4076 28927 4196 28961
rect 2253 28893 2325 28927
rect 4076 28893 4128 28927
rect 4681 28854 13118 29124
rect 4681 28820 5179 28854
rect 5213 28820 5248 28854
rect 5282 28820 5317 28854
rect 5351 28820 5386 28854
rect 5420 28820 5455 28854
rect 5489 28820 5524 28854
rect 5558 28820 5593 28854
rect 5627 28820 5662 28854
rect 5696 28820 5731 28854
rect 5765 28820 5800 28854
rect 5834 28820 5869 28854
rect 5903 28820 5938 28854
rect 5972 28820 6007 28854
rect 6041 28820 6075 28854
rect 6109 28820 6143 28854
rect 6177 28820 6211 28854
rect 6245 28820 6279 28854
rect 6313 28820 6347 28854
rect 6381 28820 6415 28854
rect 6449 28820 6483 28854
rect 6517 28820 6551 28854
rect 6585 28820 6619 28854
rect 6653 28820 6687 28854
rect 6721 28820 6755 28854
rect 6789 28820 6823 28854
rect 6857 28820 6891 28854
rect 6925 28820 6959 28854
rect 6993 28820 7027 28854
rect 7061 28820 7095 28854
rect 7129 28820 7163 28854
rect 7197 28820 7231 28854
rect 7265 28820 7299 28854
rect 7333 28820 7367 28854
rect 7401 28820 7435 28854
rect 7469 28820 7503 28854
rect 7537 28820 7571 28854
rect 7605 28820 7639 28854
rect 7673 28820 7707 28854
rect 7741 28820 7775 28854
rect 7809 28820 7843 28854
rect 7877 28820 7911 28854
rect 7945 28820 7979 28854
rect 8013 28820 8047 28854
rect 8081 28820 8115 28854
rect 8149 28820 8183 28854
rect 8217 28820 8251 28854
rect 8285 28820 8319 28854
rect 8353 28820 8387 28854
rect 8421 28820 8455 28854
rect 8489 28820 8523 28854
rect 8557 28820 8591 28854
rect 8625 28820 8659 28854
rect 8693 28820 8727 28854
rect 8761 28820 8795 28854
rect 8829 28820 8863 28854
rect 8897 28820 8931 28854
rect 8965 28820 8999 28854
rect 9033 28820 9067 28854
rect 9101 28820 9135 28854
rect 9169 28820 9203 28854
rect 9237 28820 9271 28854
rect 9305 28820 9339 28854
rect 9373 28820 9407 28854
rect 9441 28820 9475 28854
rect 9509 28820 9543 28854
rect 9577 28820 9611 28854
rect 9645 28820 9679 28854
rect 9713 28820 9747 28854
rect 9781 28820 9815 28854
rect 9849 28820 9883 28854
rect 9917 28820 9951 28854
rect 9985 28820 10019 28854
rect 10053 28820 10087 28854
rect 10121 28820 10155 28854
rect 10189 28820 10223 28854
rect 10257 28820 10291 28854
rect 10325 28820 10359 28854
rect 10393 28820 10427 28854
rect 10461 28820 10495 28854
rect 10529 28820 10563 28854
rect 10597 28820 10631 28854
rect 10665 28820 10699 28854
rect 10733 28820 10767 28854
rect 10801 28820 10835 28854
rect 10869 28820 10903 28854
rect 10937 28820 10971 28854
rect 11005 28820 11039 28854
rect 11073 28820 11107 28854
rect 11141 28820 11175 28854
rect 11209 28820 11243 28854
rect 11277 28820 11311 28854
rect 11345 28820 11379 28854
rect 11413 28820 11447 28854
rect 11481 28820 11515 28854
rect 11549 28820 11583 28854
rect 11617 28820 11651 28854
rect 11685 28820 11719 28854
rect 11753 28820 11787 28854
rect 11821 28820 11855 28854
rect 11889 28820 11923 28854
rect 11957 28820 11991 28854
rect 12025 28820 12059 28854
rect 12093 28820 12127 28854
rect 12161 28820 12195 28854
rect 12229 28820 12263 28854
rect 12297 28820 12331 28854
rect 12365 28820 12399 28854
rect 12433 28820 12467 28854
rect 12501 28820 12535 28854
rect 12569 28820 12603 28854
rect 12637 28820 12671 28854
rect 12705 28820 12739 28854
rect 12773 28820 12807 28854
rect 12841 28820 12875 28854
rect 12909 28820 12943 28854
rect 12977 28820 13118 28854
rect 5265 28714 5367 28726
rect 6101 28714 6203 28726
rect 6937 28714 7039 28726
rect 7773 28714 7875 28726
rect 8609 28714 8711 28726
rect 9445 28714 9547 28726
rect 10281 28714 10383 28726
rect 11117 28714 11219 28726
rect 11953 28714 12055 28726
rect 12789 28714 12891 28726
rect 4879 28680 4917 28714
rect 4845 28641 4951 28680
rect 4879 28607 4917 28641
rect 4845 28568 4951 28607
rect 4879 28534 4917 28568
rect 4845 28495 4951 28534
rect 4879 28461 4917 28495
rect 4845 28422 4951 28461
rect 5297 28680 5335 28714
rect 5263 28641 5369 28680
rect 5297 28607 5335 28641
rect 5263 28568 5369 28607
rect 5297 28534 5335 28568
rect 5263 28495 5369 28534
rect 5297 28461 5335 28495
rect 5263 28422 5369 28461
rect 5715 28680 5753 28714
rect 5681 28641 5787 28680
rect 5715 28607 5753 28641
rect 5681 28568 5787 28607
rect 5715 28534 5753 28568
rect 5681 28495 5787 28534
rect 5715 28461 5753 28495
rect 5681 28422 5787 28461
rect 6133 28680 6171 28714
rect 6099 28641 6205 28680
rect 6133 28607 6171 28641
rect 6099 28568 6205 28607
rect 6133 28534 6171 28568
rect 6099 28495 6205 28534
rect 6133 28461 6171 28495
rect 6099 28422 6205 28461
rect 6551 28680 6589 28714
rect 6517 28641 6623 28680
rect 6551 28607 6589 28641
rect 6517 28568 6623 28607
rect 6551 28534 6589 28568
rect 6517 28495 6623 28534
rect 6551 28461 6589 28495
rect 6517 28422 6623 28461
rect 6969 28680 7007 28714
rect 6935 28641 7041 28680
rect 6969 28607 7007 28641
rect 6935 28568 7041 28607
rect 6969 28534 7007 28568
rect 6935 28495 7041 28534
rect 6969 28461 7007 28495
rect 6935 28422 7041 28461
rect 7387 28680 7425 28714
rect 7353 28641 7459 28680
rect 7387 28607 7425 28641
rect 7353 28568 7459 28607
rect 7387 28534 7425 28568
rect 7353 28495 7459 28534
rect 7387 28461 7425 28495
rect 7353 28422 7459 28461
rect 7805 28680 7843 28714
rect 7771 28641 7877 28680
rect 7805 28607 7843 28641
rect 7771 28568 7877 28607
rect 7805 28534 7843 28568
rect 7771 28495 7877 28534
rect 7805 28461 7843 28495
rect 7771 28422 7877 28461
rect 8223 28680 8261 28714
rect 8189 28641 8295 28680
rect 8223 28607 8261 28641
rect 8189 28568 8295 28607
rect 8223 28534 8261 28568
rect 8189 28495 8295 28534
rect 8223 28461 8261 28495
rect 8189 28422 8295 28461
rect 8641 28680 8679 28714
rect 8607 28641 8713 28680
rect 8641 28607 8679 28641
rect 8607 28568 8713 28607
rect 8641 28534 8679 28568
rect 8607 28495 8713 28534
rect 8641 28461 8679 28495
rect 8607 28422 8713 28461
rect 9059 28680 9097 28714
rect 9025 28641 9131 28680
rect 9059 28607 9097 28641
rect 9025 28568 9131 28607
rect 9059 28534 9097 28568
rect 9025 28495 9131 28534
rect 9059 28461 9097 28495
rect 9025 28422 9131 28461
rect 9477 28680 9515 28714
rect 9443 28641 9549 28680
rect 9477 28607 9515 28641
rect 9443 28568 9549 28607
rect 9477 28534 9515 28568
rect 9443 28495 9549 28534
rect 9477 28461 9515 28495
rect 9443 28422 9549 28461
rect 9895 28680 9933 28714
rect 9861 28641 9967 28680
rect 9895 28607 9933 28641
rect 9861 28568 9967 28607
rect 9895 28534 9933 28568
rect 9861 28495 9967 28534
rect 9895 28461 9933 28495
rect 9861 28422 9967 28461
rect 10313 28680 10351 28714
rect 10279 28641 10385 28680
rect 10313 28607 10351 28641
rect 10279 28568 10385 28607
rect 10313 28534 10351 28568
rect 10279 28495 10385 28534
rect 10313 28461 10351 28495
rect 10279 28422 10385 28461
rect 10731 28680 10769 28714
rect 10697 28641 10803 28680
rect 10731 28607 10769 28641
rect 10697 28568 10803 28607
rect 10731 28534 10769 28568
rect 10697 28495 10803 28534
rect 10731 28461 10769 28495
rect 10697 28422 10803 28461
rect 11149 28680 11187 28714
rect 11115 28641 11221 28680
rect 11149 28607 11187 28641
rect 11115 28568 11221 28607
rect 11149 28534 11187 28568
rect 11115 28495 11221 28534
rect 11149 28461 11187 28495
rect 11115 28422 11221 28461
rect 11567 28680 11605 28714
rect 11533 28641 11639 28680
rect 11567 28607 11605 28641
rect 11533 28568 11639 28607
rect 11567 28534 11605 28568
rect 11533 28495 11639 28534
rect 11567 28461 11605 28495
rect 11533 28422 11639 28461
rect 11985 28680 12023 28714
rect 11951 28641 12057 28680
rect 11985 28607 12023 28641
rect 11951 28568 12057 28607
rect 11985 28534 12023 28568
rect 11951 28495 12057 28534
rect 11985 28461 12023 28495
rect 11951 28422 12057 28461
rect 12403 28680 12441 28714
rect 12369 28641 12475 28680
rect 12403 28607 12441 28641
rect 12369 28568 12475 28607
rect 12403 28534 12441 28568
rect 12369 28495 12475 28534
rect 12403 28461 12441 28495
rect 12369 28422 12475 28461
rect 12821 28680 12859 28714
rect 12787 28641 12893 28680
rect 12821 28607 12859 28641
rect 12787 28568 12893 28607
rect 12821 28534 12859 28568
rect 12787 28495 12893 28534
rect 12821 28461 12859 28495
rect 12787 28422 12893 28461
rect 13239 28680 13277 28714
rect 13205 28641 13311 28680
rect 13239 28607 13277 28641
rect 13205 28568 13311 28607
rect 13239 28534 13277 28568
rect 13205 28495 13311 28534
rect 13239 28461 13277 28495
rect 13205 28422 13311 28461
rect 5265 27368 5367 27380
rect 6101 27368 6203 27380
rect 6937 27368 7039 27380
rect 7773 27368 7875 27380
rect 8609 27368 8711 27380
rect 9445 27368 9547 27380
rect 10281 27368 10383 27380
rect 11117 27368 11219 27380
rect 11953 27368 12055 27380
rect 12789 27368 12891 27380
rect 4338 27321 5179 27324
rect 4338 27287 4339 27321
rect 4373 27287 4415 27321
rect 4449 27287 4491 27321
rect 4525 27290 5179 27321
rect 5213 27290 5248 27324
rect 5282 27290 5317 27324
rect 5351 27290 5386 27324
rect 5420 27290 5455 27324
rect 5489 27290 5524 27324
rect 5558 27290 5593 27324
rect 5627 27290 5662 27324
rect 5696 27290 5731 27324
rect 5765 27290 5800 27324
rect 5834 27290 5869 27324
rect 5903 27290 5938 27324
rect 5972 27290 6007 27324
rect 6041 27290 6075 27324
rect 6109 27290 6143 27324
rect 6177 27290 6211 27324
rect 6245 27290 6279 27324
rect 6313 27290 6347 27324
rect 6381 27290 6415 27324
rect 6449 27290 6483 27324
rect 6517 27290 6551 27324
rect 6585 27290 6619 27324
rect 6653 27290 6687 27324
rect 6721 27290 6755 27324
rect 6789 27290 6823 27324
rect 6857 27290 6891 27324
rect 6925 27290 6959 27324
rect 6993 27290 7027 27324
rect 7061 27290 7095 27324
rect 7129 27290 7163 27324
rect 7197 27290 7231 27324
rect 7265 27290 7299 27324
rect 7333 27290 7367 27324
rect 7401 27290 7435 27324
rect 7469 27290 7503 27324
rect 7537 27290 7571 27324
rect 7605 27290 7639 27324
rect 7673 27290 7707 27324
rect 7741 27290 7775 27324
rect 7809 27290 7843 27324
rect 7877 27290 7911 27324
rect 7945 27290 7979 27324
rect 8013 27290 8047 27324
rect 8081 27290 8115 27324
rect 8149 27290 8183 27324
rect 8217 27290 8251 27324
rect 8285 27290 8319 27324
rect 8353 27290 8387 27324
rect 8421 27290 8455 27324
rect 8489 27290 8523 27324
rect 8557 27290 8591 27324
rect 8625 27290 8659 27324
rect 8693 27290 8727 27324
rect 8761 27290 8795 27324
rect 8829 27290 8863 27324
rect 8897 27290 8931 27324
rect 8965 27290 8999 27324
rect 9033 27290 9067 27324
rect 9101 27290 9135 27324
rect 9169 27290 9203 27324
rect 9237 27290 9271 27324
rect 9305 27290 9339 27324
rect 9373 27290 9407 27324
rect 9441 27290 9475 27324
rect 9509 27290 9543 27324
rect 9577 27290 9611 27324
rect 9645 27290 9679 27324
rect 9713 27290 9747 27324
rect 9781 27290 9815 27324
rect 9849 27290 9883 27324
rect 9917 27290 9951 27324
rect 9985 27290 10019 27324
rect 10053 27290 10087 27324
rect 10121 27290 10155 27324
rect 10189 27290 10223 27324
rect 10257 27290 10291 27324
rect 10325 27290 10359 27324
rect 10393 27290 10427 27324
rect 10461 27290 10495 27324
rect 10529 27290 10563 27324
rect 10597 27290 10631 27324
rect 10665 27290 10699 27324
rect 10733 27290 10767 27324
rect 10801 27290 10835 27324
rect 10869 27290 10903 27324
rect 10937 27290 10971 27324
rect 11005 27290 11039 27324
rect 11073 27290 11107 27324
rect 11141 27290 11175 27324
rect 11209 27290 11243 27324
rect 11277 27290 11311 27324
rect 11345 27290 11379 27324
rect 11413 27290 11447 27324
rect 11481 27290 11515 27324
rect 11549 27290 11583 27324
rect 11617 27290 11651 27324
rect 11685 27290 11719 27324
rect 11753 27290 11787 27324
rect 11821 27290 11855 27324
rect 11889 27290 11923 27324
rect 11957 27290 11991 27324
rect 12025 27290 12059 27324
rect 12093 27290 12127 27324
rect 12161 27290 12195 27324
rect 12229 27290 12263 27324
rect 12297 27290 12331 27324
rect 12365 27290 12399 27324
rect 12433 27290 12467 27324
rect 12501 27290 12535 27324
rect 12569 27290 12603 27324
rect 12637 27290 12671 27324
rect 12705 27290 12739 27324
rect 12773 27290 12807 27324
rect 12841 27290 12875 27324
rect 12909 27290 12943 27324
rect 12977 27290 13118 27324
rect 4525 27287 13118 27290
rect 4338 27244 13118 27287
rect 4338 27210 4339 27244
rect 4373 27210 4415 27244
rect 4449 27210 4491 27244
rect 4525 27210 13118 27244
rect 4338 27167 13118 27210
rect 4338 27133 4339 27167
rect 4373 27133 4415 27167
rect 4449 27133 4491 27167
rect 4525 27133 13118 27167
rect 4338 27089 13118 27133
rect 4338 27055 4339 27089
rect 4373 27055 4415 27089
rect 4449 27055 4491 27089
rect 4525 27055 13118 27089
rect 4338 27011 13118 27055
rect 4338 26977 4339 27011
rect 4373 26977 4415 27011
rect 4449 26977 4491 27011
rect 4525 26977 13118 27011
rect 4338 26933 13118 26977
rect 4338 26899 4339 26933
rect 4373 26899 4415 26933
rect 4449 26899 4491 26933
rect 4525 26899 13118 26933
rect 4338 26855 13118 26899
rect 4338 26821 4339 26855
rect 4373 26821 4415 26855
rect 4449 26821 4491 26855
rect 4525 26854 13118 26855
rect 4525 26821 5179 26854
rect 4338 26820 5179 26821
rect 5213 26820 5248 26854
rect 5282 26820 5317 26854
rect 5351 26820 5386 26854
rect 5420 26820 5455 26854
rect 5489 26820 5524 26854
rect 5558 26820 5593 26854
rect 5627 26820 5662 26854
rect 5696 26820 5731 26854
rect 5765 26820 5800 26854
rect 5834 26820 5869 26854
rect 5903 26820 5938 26854
rect 5972 26820 6007 26854
rect 6041 26820 6075 26854
rect 6109 26820 6143 26854
rect 6177 26820 6211 26854
rect 6245 26820 6279 26854
rect 6313 26820 6347 26854
rect 6381 26820 6415 26854
rect 6449 26820 6483 26854
rect 6517 26820 6551 26854
rect 6585 26820 6619 26854
rect 6653 26820 6687 26854
rect 6721 26820 6755 26854
rect 6789 26820 6823 26854
rect 6857 26820 6891 26854
rect 6925 26820 6959 26854
rect 6993 26820 7027 26854
rect 7061 26820 7095 26854
rect 7129 26820 7163 26854
rect 7197 26820 7231 26854
rect 7265 26820 7299 26854
rect 7333 26820 7367 26854
rect 7401 26820 7435 26854
rect 7469 26820 7503 26854
rect 7537 26820 7571 26854
rect 7605 26820 7639 26854
rect 7673 26820 7707 26854
rect 7741 26820 7775 26854
rect 7809 26820 7843 26854
rect 7877 26820 7911 26854
rect 7945 26820 7979 26854
rect 8013 26820 8047 26854
rect 8081 26820 8115 26854
rect 8149 26820 8183 26854
rect 8217 26820 8251 26854
rect 8285 26820 8319 26854
rect 8353 26820 8387 26854
rect 8421 26820 8455 26854
rect 8489 26820 8523 26854
rect 8557 26820 8591 26854
rect 8625 26820 8659 26854
rect 8693 26820 8727 26854
rect 8761 26820 8795 26854
rect 8829 26820 8863 26854
rect 8897 26820 8931 26854
rect 8965 26820 8999 26854
rect 9033 26820 9067 26854
rect 9101 26820 9135 26854
rect 9169 26820 9203 26854
rect 9237 26820 9271 26854
rect 9305 26820 9339 26854
rect 9373 26820 9407 26854
rect 9441 26820 9475 26854
rect 9509 26820 9543 26854
rect 9577 26820 9611 26854
rect 9645 26820 9679 26854
rect 9713 26820 9747 26854
rect 9781 26820 9815 26854
rect 9849 26820 9883 26854
rect 9917 26820 9951 26854
rect 9985 26820 10019 26854
rect 10053 26820 10087 26854
rect 10121 26820 10155 26854
rect 10189 26820 10223 26854
rect 10257 26820 10291 26854
rect 10325 26820 10359 26854
rect 10393 26820 10427 26854
rect 10461 26820 10495 26854
rect 10529 26820 10563 26854
rect 10597 26820 10631 26854
rect 10665 26820 10699 26854
rect 10733 26820 10767 26854
rect 10801 26820 10835 26854
rect 10869 26820 10903 26854
rect 10937 26820 10971 26854
rect 11005 26820 11039 26854
rect 11073 26820 11107 26854
rect 11141 26820 11175 26854
rect 11209 26820 11243 26854
rect 11277 26820 11311 26854
rect 11345 26820 11379 26854
rect 11413 26820 11447 26854
rect 11481 26820 11515 26854
rect 11549 26820 11583 26854
rect 11617 26820 11651 26854
rect 11685 26820 11719 26854
rect 11753 26820 11787 26854
rect 11821 26820 11855 26854
rect 11889 26820 11923 26854
rect 11957 26820 11991 26854
rect 12025 26820 12059 26854
rect 12093 26820 12127 26854
rect 12161 26820 12195 26854
rect 12229 26820 12263 26854
rect 12297 26820 12331 26854
rect 12365 26820 12399 26854
rect 12433 26820 12467 26854
rect 12501 26820 12535 26854
rect 12569 26820 12603 26854
rect 12637 26820 12671 26854
rect 12705 26820 12739 26854
rect 12773 26820 12807 26854
rect 12841 26820 12875 26854
rect 12909 26820 12943 26854
rect 12977 26820 13118 26854
rect 4879 26718 4917 26752
rect 4845 26677 4951 26718
rect 4879 26643 4917 26677
rect 4845 26602 4951 26643
rect 4879 26568 4917 26602
rect 4845 26527 4951 26568
rect 4879 26493 4917 26527
rect 4845 26452 4951 26493
rect 4879 26418 4917 26452
rect 4845 26377 4951 26418
rect 4879 26343 4917 26377
rect 4845 26302 4951 26343
rect 4879 26268 4917 26302
rect 4845 26227 4951 26268
rect 4879 26193 4917 26227
rect 4845 26152 4951 26193
rect 4879 26118 4917 26152
rect 4845 26077 4951 26118
rect 4879 26043 4917 26077
rect 4845 26002 4951 26043
rect 4879 25968 4917 26002
rect 4845 25928 4951 25968
rect 4879 25894 4917 25928
rect 4845 25854 4951 25894
rect 4879 25820 4917 25854
rect 4845 25780 4951 25820
rect 4879 25746 4917 25780
rect 5297 26709 5335 26743
rect 5263 26668 5369 26709
rect 5297 26634 5335 26668
rect 5263 26594 5369 26634
rect 5297 26560 5335 26594
rect 5263 26520 5369 26560
rect 5297 26486 5335 26520
rect 5263 26446 5369 26486
rect 5297 26412 5335 26446
rect 5263 26372 5369 26412
rect 5297 26338 5335 26372
rect 5263 26298 5369 26338
rect 5297 26264 5335 26298
rect 5263 26224 5369 26264
rect 5297 26190 5335 26224
rect 5263 26150 5369 26190
rect 5297 26116 5335 26150
rect 5263 26076 5369 26116
rect 5297 26042 5335 26076
rect 5263 26002 5369 26042
rect 5297 25968 5335 26002
rect 5263 25928 5369 25968
rect 5297 25894 5335 25928
rect 5263 25854 5369 25894
rect 5297 25820 5335 25854
rect 5263 25780 5369 25820
rect 5297 25746 5335 25780
rect 5715 26718 5753 26752
rect 5681 26679 5787 26718
rect 5715 26645 5753 26679
rect 5681 26606 5787 26645
rect 5715 26572 5753 26606
rect 5681 26533 5787 26572
rect 5715 26499 5753 26533
rect 5681 26460 5787 26499
rect 5715 26426 5753 26460
rect 5681 26387 5787 26426
rect 5715 26353 5753 26387
rect 5681 26314 5787 26353
rect 5715 26280 5753 26314
rect 5681 26241 5787 26280
rect 5715 26207 5753 26241
rect 5681 26168 5787 26207
rect 5715 26134 5753 26168
rect 5681 26095 5787 26134
rect 5715 26061 5753 26095
rect 5681 26022 5787 26061
rect 6133 26709 6171 26743
rect 6099 26668 6205 26709
rect 6133 26634 6171 26668
rect 6099 26594 6205 26634
rect 6133 26560 6171 26594
rect 6099 26520 6205 26560
rect 6133 26486 6171 26520
rect 6099 26446 6205 26486
rect 6133 26412 6171 26446
rect 6099 26372 6205 26412
rect 6133 26338 6171 26372
rect 6099 26298 6205 26338
rect 6133 26264 6171 26298
rect 6099 26224 6205 26264
rect 6133 26190 6171 26224
rect 6099 26150 6205 26190
rect 6133 26116 6171 26150
rect 6099 26076 6205 26116
rect 6133 26042 6171 26076
rect 6099 26002 6205 26042
rect 6133 25968 6171 26002
rect 6099 25928 6205 25968
rect 6133 25894 6171 25928
rect 6099 25854 6205 25894
rect 6133 25820 6171 25854
rect 6099 25780 6205 25820
rect 6133 25746 6171 25780
rect 6551 26717 6589 26751
rect 6517 26676 6623 26717
rect 6551 26642 6589 26676
rect 6517 26601 6623 26642
rect 6551 26567 6589 26601
rect 6517 26526 6623 26567
rect 6551 26492 6589 26526
rect 6517 26451 6623 26492
rect 6551 26417 6589 26451
rect 6517 26376 6623 26417
rect 6551 26342 6589 26376
rect 6517 26301 6623 26342
rect 6551 26267 6589 26301
rect 6517 26226 6623 26267
rect 6551 26192 6589 26226
rect 6517 26151 6623 26192
rect 6551 26117 6589 26151
rect 6517 26076 6623 26117
rect 6551 26042 6589 26076
rect 6517 26002 6623 26042
rect 6551 25968 6589 26002
rect 6517 25928 6623 25968
rect 6551 25894 6589 25928
rect 6517 25854 6623 25894
rect 6551 25820 6589 25854
rect 6517 25780 6623 25820
rect 6551 25746 6589 25780
rect 6969 26734 7007 26768
rect 7805 26751 7843 26785
rect 8641 26751 8679 26785
rect 9477 26751 9515 26785
rect 10313 26751 10351 26785
rect 11149 26751 11187 26785
rect 11985 26751 12023 26785
rect 12821 26751 12859 26785
rect 6935 26692 7041 26734
rect 6969 26658 7007 26692
rect 6935 26616 7041 26658
rect 6969 26582 7007 26616
rect 6935 26540 7041 26582
rect 6969 26506 7007 26540
rect 6935 26464 7041 26506
rect 6969 26430 7007 26464
rect 6935 26388 7041 26430
rect 6969 26354 7007 26388
rect 6935 26312 7041 26354
rect 6969 26278 7007 26312
rect 6935 26236 7041 26278
rect 6969 26202 7007 26236
rect 6935 26160 7041 26202
rect 6969 26126 7007 26160
rect 6935 26084 7041 26126
rect 6969 26050 7007 26084
rect 6935 26008 7041 26050
rect 6969 25974 7007 26008
rect 6935 25932 7041 25974
rect 6969 25898 7007 25932
rect 6935 25856 7041 25898
rect 6969 25822 7007 25856
rect 6935 25780 7041 25822
rect 6969 25746 7007 25780
rect 7387 26717 7425 26751
rect 7353 26676 7459 26717
rect 7387 26642 7425 26676
rect 7353 26601 7459 26642
rect 7387 26567 7425 26601
rect 7353 26526 7459 26567
rect 7387 26492 7425 26526
rect 7353 26451 7459 26492
rect 7387 26417 7425 26451
rect 7353 26376 7459 26417
rect 7387 26342 7425 26376
rect 7353 26301 7459 26342
rect 7387 26267 7425 26301
rect 7353 26226 7459 26267
rect 7387 26192 7425 26226
rect 7353 26151 7459 26192
rect 7387 26117 7425 26151
rect 7353 26076 7459 26117
rect 7387 26042 7425 26076
rect 7353 26002 7459 26042
rect 7387 25968 7425 26002
rect 7353 25928 7459 25968
rect 7387 25894 7425 25928
rect 7353 25854 7459 25894
rect 7387 25820 7425 25854
rect 7353 25780 7459 25820
rect 7387 25746 7425 25780
rect 7771 26707 7877 26751
rect 7805 26673 7843 26707
rect 7771 26629 7877 26673
rect 7805 26595 7843 26629
rect 7771 26551 7877 26595
rect 7805 26517 7843 26551
rect 7771 26473 7877 26517
rect 7805 26439 7843 26473
rect 7771 26396 7877 26439
rect 7805 26362 7843 26396
rect 7771 26319 7877 26362
rect 7805 26285 7843 26319
rect 7771 26242 7877 26285
rect 7805 26208 7843 26242
rect 7771 26165 7877 26208
rect 7805 26131 7843 26165
rect 7771 26088 7877 26131
rect 7805 26054 7843 26088
rect 7771 26011 7877 26054
rect 7805 25977 7843 26011
rect 7771 25934 7877 25977
rect 7805 25900 7843 25934
rect 7771 25857 7877 25900
rect 7805 25823 7843 25857
rect 7771 25780 7877 25823
rect 7805 25746 7843 25780
rect 8223 26717 8261 26751
rect 8189 26676 8295 26717
rect 8223 26642 8261 26676
rect 8189 26601 8295 26642
rect 8223 26567 8261 26601
rect 8189 26526 8295 26567
rect 8223 26492 8261 26526
rect 8189 26451 8295 26492
rect 8223 26417 8261 26451
rect 8189 26376 8295 26417
rect 8223 26342 8261 26376
rect 8189 26301 8295 26342
rect 8223 26267 8261 26301
rect 8189 26226 8295 26267
rect 8223 26192 8261 26226
rect 8189 26151 8295 26192
rect 8223 26117 8261 26151
rect 8189 26076 8295 26117
rect 8223 26042 8261 26076
rect 8189 26002 8295 26042
rect 8223 25968 8261 26002
rect 8189 25928 8295 25968
rect 8223 25894 8261 25928
rect 8189 25854 8295 25894
rect 8223 25820 8261 25854
rect 8189 25780 8295 25820
rect 8223 25746 8261 25780
rect 8607 26707 8713 26751
rect 8641 26673 8679 26707
rect 8607 26629 8713 26673
rect 8641 26595 8679 26629
rect 8607 26551 8713 26595
rect 8641 26517 8679 26551
rect 8607 26473 8713 26517
rect 8641 26439 8679 26473
rect 8607 26396 8713 26439
rect 8641 26362 8679 26396
rect 8607 26319 8713 26362
rect 8641 26285 8679 26319
rect 8607 26242 8713 26285
rect 8641 26208 8679 26242
rect 8607 26165 8713 26208
rect 8641 26131 8679 26165
rect 8607 26088 8713 26131
rect 8641 26054 8679 26088
rect 8607 26011 8713 26054
rect 8641 25977 8679 26011
rect 8607 25934 8713 25977
rect 8641 25900 8679 25934
rect 8607 25857 8713 25900
rect 8641 25823 8679 25857
rect 8607 25780 8713 25823
rect 8641 25746 8679 25780
rect 9059 26717 9097 26751
rect 9025 26676 9131 26717
rect 9059 26642 9097 26676
rect 9025 26601 9131 26642
rect 9059 26567 9097 26601
rect 9025 26526 9131 26567
rect 9059 26492 9097 26526
rect 9025 26451 9131 26492
rect 9059 26417 9097 26451
rect 9025 26376 9131 26417
rect 9059 26342 9097 26376
rect 9025 26301 9131 26342
rect 9059 26267 9097 26301
rect 9025 26226 9131 26267
rect 9059 26192 9097 26226
rect 9025 26151 9131 26192
rect 9059 26117 9097 26151
rect 9025 26076 9131 26117
rect 9059 26042 9097 26076
rect 9025 26002 9131 26042
rect 9059 25968 9097 26002
rect 9025 25928 9131 25968
rect 9059 25894 9097 25928
rect 9025 25854 9131 25894
rect 9059 25820 9097 25854
rect 9025 25780 9131 25820
rect 9059 25746 9097 25780
rect 9443 26707 9549 26751
rect 9477 26673 9515 26707
rect 9443 26629 9549 26673
rect 9477 26595 9515 26629
rect 9443 26551 9549 26595
rect 9477 26517 9515 26551
rect 9443 26473 9549 26517
rect 9477 26439 9515 26473
rect 9443 26396 9549 26439
rect 9477 26362 9515 26396
rect 9443 26319 9549 26362
rect 9477 26285 9515 26319
rect 9443 26242 9549 26285
rect 9477 26208 9515 26242
rect 9443 26165 9549 26208
rect 9477 26131 9515 26165
rect 9443 26088 9549 26131
rect 9477 26054 9515 26088
rect 9443 26011 9549 26054
rect 9477 25977 9515 26011
rect 9443 25934 9549 25977
rect 9477 25900 9515 25934
rect 9443 25857 9549 25900
rect 9477 25823 9515 25857
rect 9443 25780 9549 25823
rect 9477 25746 9515 25780
rect 9895 26717 9933 26751
rect 9861 26676 9967 26717
rect 9895 26642 9933 26676
rect 9861 26601 9967 26642
rect 9895 26567 9933 26601
rect 9861 26526 9967 26567
rect 9895 26492 9933 26526
rect 9861 26451 9967 26492
rect 9895 26417 9933 26451
rect 9861 26376 9967 26417
rect 9895 26342 9933 26376
rect 9861 26301 9967 26342
rect 9895 26267 9933 26301
rect 9861 26226 9967 26267
rect 9895 26192 9933 26226
rect 9861 26151 9967 26192
rect 9895 26117 9933 26151
rect 9861 26076 9967 26117
rect 9895 26042 9933 26076
rect 9861 26002 9967 26042
rect 9895 25968 9933 26002
rect 9861 25928 9967 25968
rect 9895 25894 9933 25928
rect 9861 25854 9967 25894
rect 9895 25820 9933 25854
rect 9861 25780 9967 25820
rect 9895 25746 9933 25780
rect 10279 26707 10385 26751
rect 10313 26673 10351 26707
rect 10279 26629 10385 26673
rect 10313 26595 10351 26629
rect 10279 26551 10385 26595
rect 10313 26517 10351 26551
rect 10279 26473 10385 26517
rect 10313 26439 10351 26473
rect 10279 26396 10385 26439
rect 10313 26362 10351 26396
rect 10279 26319 10385 26362
rect 10313 26285 10351 26319
rect 10279 26242 10385 26285
rect 10313 26208 10351 26242
rect 10279 26165 10385 26208
rect 10313 26131 10351 26165
rect 10279 26088 10385 26131
rect 10313 26054 10351 26088
rect 10279 26011 10385 26054
rect 10313 25977 10351 26011
rect 10279 25934 10385 25977
rect 10313 25900 10351 25934
rect 10279 25857 10385 25900
rect 10313 25823 10351 25857
rect 10279 25780 10385 25823
rect 10313 25746 10351 25780
rect 10731 26717 10769 26751
rect 10697 26676 10803 26717
rect 10731 26642 10769 26676
rect 10697 26601 10803 26642
rect 10731 26567 10769 26601
rect 10697 26526 10803 26567
rect 10731 26492 10769 26526
rect 10697 26451 10803 26492
rect 10731 26417 10769 26451
rect 10697 26376 10803 26417
rect 10731 26342 10769 26376
rect 10697 26301 10803 26342
rect 10731 26267 10769 26301
rect 10697 26226 10803 26267
rect 10731 26192 10769 26226
rect 10697 26151 10803 26192
rect 10731 26117 10769 26151
rect 10697 26076 10803 26117
rect 10731 26042 10769 26076
rect 10697 26002 10803 26042
rect 10731 25968 10769 26002
rect 10697 25928 10803 25968
rect 10731 25894 10769 25928
rect 10697 25854 10803 25894
rect 10731 25820 10769 25854
rect 10697 25780 10803 25820
rect 10731 25746 10769 25780
rect 11115 26707 11221 26751
rect 11149 26673 11187 26707
rect 11115 26629 11221 26673
rect 11149 26595 11187 26629
rect 11115 26551 11221 26595
rect 11149 26517 11187 26551
rect 11115 26473 11221 26517
rect 11149 26439 11187 26473
rect 11115 26396 11221 26439
rect 11149 26362 11187 26396
rect 11115 26319 11221 26362
rect 11149 26285 11187 26319
rect 11115 26242 11221 26285
rect 11149 26208 11187 26242
rect 11115 26165 11221 26208
rect 11149 26131 11187 26165
rect 11115 26088 11221 26131
rect 11149 26054 11187 26088
rect 11115 26011 11221 26054
rect 11149 25977 11187 26011
rect 11115 25934 11221 25977
rect 11149 25900 11187 25934
rect 11115 25857 11221 25900
rect 11149 25823 11187 25857
rect 11115 25780 11221 25823
rect 11149 25746 11187 25780
rect 11567 26717 11605 26751
rect 11533 26676 11639 26717
rect 11567 26642 11605 26676
rect 11533 26601 11639 26642
rect 11567 26567 11605 26601
rect 11533 26526 11639 26567
rect 11567 26492 11605 26526
rect 11533 26451 11639 26492
rect 11567 26417 11605 26451
rect 11533 26376 11639 26417
rect 11567 26342 11605 26376
rect 11533 26301 11639 26342
rect 11567 26267 11605 26301
rect 11533 26226 11639 26267
rect 11567 26192 11605 26226
rect 11533 26151 11639 26192
rect 11567 26117 11605 26151
rect 11533 26076 11639 26117
rect 11567 26042 11605 26076
rect 11533 26002 11639 26042
rect 11567 25968 11605 26002
rect 11533 25928 11639 25968
rect 11567 25894 11605 25928
rect 11533 25854 11639 25894
rect 11567 25820 11605 25854
rect 11533 25780 11639 25820
rect 11567 25746 11605 25780
rect 11951 26707 12057 26751
rect 11985 26673 12023 26707
rect 11951 26629 12057 26673
rect 11985 26595 12023 26629
rect 11951 26551 12057 26595
rect 11985 26517 12023 26551
rect 11951 26473 12057 26517
rect 11985 26439 12023 26473
rect 11951 26396 12057 26439
rect 11985 26362 12023 26396
rect 11951 26319 12057 26362
rect 11985 26285 12023 26319
rect 11951 26242 12057 26285
rect 11985 26208 12023 26242
rect 11951 26165 12057 26208
rect 11985 26131 12023 26165
rect 11951 26088 12057 26131
rect 11985 26054 12023 26088
rect 11951 26011 12057 26054
rect 11985 25977 12023 26011
rect 11951 25934 12057 25977
rect 11985 25900 12023 25934
rect 11951 25857 12057 25900
rect 11985 25823 12023 25857
rect 11951 25780 12057 25823
rect 11985 25746 12023 25780
rect 12403 26717 12441 26751
rect 12369 26676 12475 26717
rect 12403 26642 12441 26676
rect 12369 26601 12475 26642
rect 12403 26567 12441 26601
rect 12369 26526 12475 26567
rect 12403 26492 12441 26526
rect 12369 26451 12475 26492
rect 12403 26417 12441 26451
rect 12369 26376 12475 26417
rect 12403 26342 12441 26376
rect 12369 26301 12475 26342
rect 12403 26267 12441 26301
rect 12369 26226 12475 26267
rect 12403 26192 12441 26226
rect 12369 26151 12475 26192
rect 12403 26117 12441 26151
rect 12369 26076 12475 26117
rect 12403 26042 12441 26076
rect 12369 26002 12475 26042
rect 12403 25968 12441 26002
rect 12369 25928 12475 25968
rect 12403 25894 12441 25928
rect 12369 25854 12475 25894
rect 12403 25820 12441 25854
rect 12369 25780 12475 25820
rect 12403 25746 12441 25780
rect 12787 26707 12893 26751
rect 12821 26673 12859 26707
rect 12787 26629 12893 26673
rect 12821 26595 12859 26629
rect 12787 26551 12893 26595
rect 12821 26517 12859 26551
rect 12787 26473 12893 26517
rect 12821 26439 12859 26473
rect 12787 26396 12893 26439
rect 12821 26362 12859 26396
rect 12787 26319 12893 26362
rect 12821 26285 12859 26319
rect 12787 26242 12893 26285
rect 12821 26208 12859 26242
rect 12787 26165 12893 26208
rect 12821 26131 12859 26165
rect 12787 26088 12893 26131
rect 12821 26054 12859 26088
rect 12787 26011 12893 26054
rect 12821 25977 12859 26011
rect 12787 25934 12893 25977
rect 12821 25900 12859 25934
rect 12787 25857 12893 25900
rect 12821 25823 12859 25857
rect 12787 25780 12893 25823
rect 12821 25746 12859 25780
rect 13239 26717 13277 26751
rect 13205 26676 13311 26717
rect 13239 26642 13277 26676
rect 13205 26601 13311 26642
rect 13239 26567 13277 26601
rect 13205 26526 13311 26567
rect 13239 26492 13277 26526
rect 13205 26451 13311 26492
rect 13239 26417 13277 26451
rect 13205 26376 13311 26417
rect 13239 26342 13277 26376
rect 13205 26301 13311 26342
rect 13239 26267 13277 26301
rect 13205 26226 13311 26267
rect 13239 26192 13277 26226
rect 13205 26151 13311 26192
rect 13239 26117 13277 26151
rect 13205 26076 13311 26117
rect 13239 26042 13277 26076
rect 13205 26002 13311 26042
rect 13239 25968 13277 26002
rect 13205 25928 13311 25968
rect 13239 25894 13277 25928
rect 13205 25854 13311 25894
rect 13239 25820 13277 25854
rect 13205 25780 13311 25820
rect 13239 25746 13277 25780
rect 4332 25670 5179 25703
rect 4332 25636 4344 25670
rect 4378 25636 4486 25670
rect 4520 25669 5179 25670
rect 5213 25669 5248 25703
rect 5282 25669 5317 25703
rect 5351 25669 5386 25703
rect 5420 25669 5455 25703
rect 5489 25669 5524 25703
rect 5558 25669 5593 25703
rect 5627 25669 5662 25703
rect 5696 25669 5731 25703
rect 5765 25669 5800 25703
rect 5834 25669 5869 25703
rect 5903 25669 5938 25703
rect 5972 25669 6007 25703
rect 6041 25669 6075 25703
rect 6109 25669 6143 25703
rect 6177 25669 6211 25703
rect 6245 25669 6279 25703
rect 6313 25669 6347 25703
rect 6381 25669 6415 25703
rect 6449 25669 6483 25703
rect 6517 25669 6551 25703
rect 6585 25669 6619 25703
rect 6653 25669 6687 25703
rect 6721 25669 6755 25703
rect 6789 25669 6823 25703
rect 6857 25669 6891 25703
rect 6925 25669 6959 25703
rect 6993 25669 7027 25703
rect 7061 25669 7095 25703
rect 7129 25669 7163 25703
rect 7197 25669 7231 25703
rect 7265 25669 7299 25703
rect 7333 25669 7367 25703
rect 7401 25669 7435 25703
rect 7469 25669 7503 25703
rect 7537 25669 7571 25703
rect 7605 25669 7639 25703
rect 7673 25669 7707 25703
rect 7741 25669 7775 25703
rect 7809 25669 7843 25703
rect 7877 25669 7911 25703
rect 7945 25669 7979 25703
rect 8013 25669 8047 25703
rect 8081 25669 8115 25703
rect 8149 25669 8183 25703
rect 8217 25669 8251 25703
rect 8285 25669 8319 25703
rect 8353 25669 8387 25703
rect 8421 25669 8455 25703
rect 8489 25669 8523 25703
rect 8557 25669 8591 25703
rect 8625 25669 8659 25703
rect 8693 25669 8727 25703
rect 8761 25669 8795 25703
rect 8829 25669 8863 25703
rect 8897 25669 8931 25703
rect 8965 25669 8999 25703
rect 9033 25669 9067 25703
rect 9101 25669 9135 25703
rect 9169 25669 9203 25703
rect 9237 25669 9271 25703
rect 9305 25669 9339 25703
rect 9373 25669 9407 25703
rect 9441 25669 9475 25703
rect 9509 25669 9543 25703
rect 9577 25669 9611 25703
rect 9645 25669 9679 25703
rect 9713 25669 9747 25703
rect 9781 25669 9815 25703
rect 9849 25669 9883 25703
rect 9917 25669 9951 25703
rect 9985 25669 10019 25703
rect 10053 25669 10087 25703
rect 10121 25669 10155 25703
rect 10189 25669 10223 25703
rect 10257 25669 10291 25703
rect 10325 25669 10359 25703
rect 10393 25669 10427 25703
rect 10461 25669 10495 25703
rect 10529 25669 10563 25703
rect 10597 25669 10631 25703
rect 10665 25669 10699 25703
rect 10733 25669 10767 25703
rect 10801 25669 10835 25703
rect 10869 25669 10903 25703
rect 10937 25669 10971 25703
rect 11005 25669 11039 25703
rect 11073 25669 11107 25703
rect 11141 25669 11175 25703
rect 11209 25669 11243 25703
rect 11277 25669 11311 25703
rect 11345 25669 11379 25703
rect 11413 25669 11447 25703
rect 11481 25669 11515 25703
rect 11549 25669 11583 25703
rect 11617 25669 11651 25703
rect 11685 25669 11719 25703
rect 11753 25669 11787 25703
rect 11821 25669 11855 25703
rect 11889 25669 11923 25703
rect 11957 25669 11991 25703
rect 12025 25669 12059 25703
rect 12093 25669 12127 25703
rect 12161 25669 12195 25703
rect 12229 25669 12263 25703
rect 12297 25669 12331 25703
rect 12365 25669 12399 25703
rect 12433 25669 12467 25703
rect 12501 25669 12535 25703
rect 12569 25669 12603 25703
rect 12637 25669 12671 25703
rect 12705 25669 12739 25703
rect 12773 25669 12807 25703
rect 12841 25669 12875 25703
rect 12909 25669 12943 25703
rect 12977 25669 13118 25703
rect 4520 25636 13118 25669
rect 4332 25602 13118 25636
rect 4761 25025 4809 25149
rect 4727 24986 4809 25025
rect 4761 24952 4809 24986
rect 4727 24914 4809 24952
rect 4761 24880 4809 24914
rect 4727 24842 4809 24880
rect 4761 24808 4809 24842
rect 4727 24770 4809 24808
rect 4761 24736 4809 24770
rect 4727 24698 4809 24736
rect 4761 24664 4809 24698
rect 4727 24626 4809 24664
rect 4761 24592 4809 24626
rect 4727 24554 4809 24592
rect 4761 24520 4809 24554
rect 4727 24482 4809 24520
rect 4761 24448 4809 24482
rect 4727 24410 4809 24448
rect 4761 24376 4809 24410
rect 4727 24338 4809 24376
rect 4761 24304 4809 24338
rect 4727 24266 4809 24304
rect 4761 24232 4809 24266
rect 4727 24194 4809 24232
rect 4761 24160 4809 24194
rect 4727 24122 4809 24160
rect 4761 24088 4809 24122
rect 4727 24050 4809 24088
rect 4761 23791 4809 24050
rect 5073 24895 5107 24938
rect 5073 24818 5107 24861
rect 5073 24741 5107 24784
rect 5073 24664 5107 24707
rect 5073 24587 5107 24630
rect 5073 24510 5107 24553
rect 5073 24433 5107 24476
rect 5073 24356 5107 24399
rect 5073 24279 5107 24322
rect 5073 24202 5107 24245
rect 5073 24126 5107 24168
rect 5073 24050 5107 24092
rect 6719 24895 6753 24938
rect 6719 24818 6753 24861
rect 6719 24741 6753 24784
rect 6719 24664 6753 24707
rect 6719 24587 6753 24630
rect 6719 24510 6753 24553
rect 6719 24433 6753 24476
rect 6719 24356 6753 24399
rect 6719 24279 6753 24322
rect 6719 24202 6753 24245
rect 6719 24126 6753 24168
rect 6719 24050 6753 24092
rect 8374 24895 8408 24938
rect 8374 24818 8408 24861
rect 8374 24741 8408 24784
rect 8374 24664 8408 24707
rect 8374 24587 8408 24630
rect 8374 24510 8408 24553
rect 8374 24433 8408 24476
rect 8374 24356 8408 24399
rect 8374 24279 8408 24322
rect 8374 24202 8408 24245
rect 8374 24126 8408 24168
rect 8374 24050 8408 24092
rect 10030 24895 10064 24938
rect 10030 24818 10064 24861
rect 10030 24741 10064 24784
rect 10030 24664 10064 24707
rect 10030 24587 10064 24630
rect 10030 24510 10064 24553
rect 10030 24433 10064 24476
rect 10030 24356 10064 24399
rect 10030 24279 10064 24322
rect 10030 24202 10064 24245
rect 10030 24126 10064 24168
rect 10030 24050 10064 24092
rect 11686 24895 11720 24938
rect 11686 24818 11720 24861
rect 11686 24741 11720 24784
rect 11686 24664 11720 24707
rect 11686 24587 11720 24630
rect 11686 24510 11720 24553
rect 11686 24433 11720 24476
rect 11686 24356 11720 24399
rect 11686 24279 11720 24322
rect 11686 24202 11720 24245
rect 11686 24126 11720 24168
rect 11686 24050 11720 24092
rect 13342 24895 13376 24938
rect 13342 24818 13376 24861
rect 13342 24741 13376 24784
rect 13342 24664 13376 24707
rect 13342 24587 13376 24630
rect 13342 24510 13376 24553
rect 13342 24433 13376 24476
rect 13342 24356 13376 24399
rect 13342 24279 13376 24322
rect 13342 24202 13376 24245
rect 13342 24126 13376 24168
rect 13342 24050 13376 24092
rect 4934 23663 4954 23697
rect 4988 23663 5022 23697
rect 5056 23663 5081 23697
rect 5124 23663 5154 23697
rect 5192 23663 5226 23697
rect 5261 23663 5294 23697
rect 5334 23663 5362 23697
rect 5407 23663 5430 23697
rect 5480 23663 5498 23697
rect 5553 23663 5566 23697
rect 5626 23663 5634 23697
rect 5699 23663 5702 23697
rect 5736 23663 5737 23697
rect 5804 23663 5809 23697
rect 5872 23663 5881 23697
rect 5940 23663 5953 23697
rect 6008 23663 6025 23697
rect 6076 23663 6097 23697
rect 6144 23663 6169 23697
rect 6212 23663 6241 23697
rect 6280 23663 6313 23697
rect 6348 23663 6382 23697
rect 6419 23663 6450 23697
rect 6491 23663 6518 23697
rect 6563 23663 6586 23697
rect 6635 23663 6654 23697
rect 6707 23663 6722 23697
rect 6779 23663 6790 23697
rect 6851 23663 6858 23697
rect 6923 23663 6926 23697
rect 6960 23663 6961 23697
rect 7028 23663 7033 23697
rect 7096 23663 7105 23697
rect 7164 23663 7177 23697
rect 7232 23663 7249 23697
rect 7300 23663 7321 23697
rect 7368 23663 7393 23697
rect 7436 23663 7465 23697
rect 7504 23663 7537 23697
rect 7572 23663 7606 23697
rect 7643 23663 7674 23697
rect 7715 23663 7742 23697
rect 7787 23663 7810 23697
rect 7859 23663 7878 23697
rect 7931 23663 7946 23697
rect 8003 23663 8014 23697
rect 8075 23663 8082 23697
rect 8147 23663 8150 23697
rect 8184 23663 8185 23697
rect 8252 23663 8257 23697
rect 8320 23663 8329 23697
rect 8388 23663 8401 23697
rect 8456 23663 8473 23697
rect 8524 23663 8545 23697
rect 8592 23663 8617 23697
rect 8660 23663 8689 23697
rect 8728 23663 8761 23697
rect 8796 23663 8830 23697
rect 8867 23663 8898 23697
rect 8939 23663 8966 23697
rect 9011 23663 9034 23697
rect 9083 23663 9102 23697
rect 9155 23663 9170 23697
rect 9227 23663 9238 23697
rect 9299 23663 9306 23697
rect 9371 23663 9374 23697
rect 9408 23663 9409 23697
rect 9476 23663 9481 23697
rect 9544 23663 9553 23697
rect 9612 23663 9625 23697
rect 9680 23663 9697 23697
rect 9748 23663 9769 23697
rect 9816 23663 9841 23697
rect 9884 23663 9913 23697
rect 9952 23663 9985 23697
rect 10020 23663 10054 23697
rect 10091 23663 10122 23697
rect 10163 23663 10190 23697
rect 10235 23663 10258 23697
rect 10307 23663 10326 23697
rect 10379 23663 10394 23697
rect 10451 23663 10462 23697
rect 10523 23663 10530 23697
rect 10595 23663 10598 23697
rect 10632 23663 10633 23697
rect 10700 23663 10705 23697
rect 10768 23663 10777 23697
rect 10836 23663 10849 23697
rect 10904 23663 10921 23697
rect 10972 23663 10993 23697
rect 11040 23663 11065 23697
rect 11108 23663 11137 23697
rect 11176 23663 11209 23697
rect 11244 23663 11278 23697
rect 11315 23663 11346 23697
rect 11387 23663 11414 23697
rect 11459 23663 11482 23697
rect 11531 23663 11550 23697
rect 11603 23663 11618 23697
rect 11675 23663 11686 23697
rect 11747 23663 11754 23697
rect 11819 23663 11822 23697
rect 11856 23663 11857 23697
rect 11924 23663 11929 23697
rect 11992 23663 12001 23697
rect 12060 23663 12073 23697
rect 12128 23663 12145 23697
rect 12196 23663 12217 23697
rect 12264 23663 12289 23697
rect 12332 23663 12361 23697
rect 12400 23663 12433 23697
rect 12468 23663 12502 23697
rect 12539 23663 12570 23697
rect 12611 23663 12638 23697
rect 12683 23663 12706 23697
rect 12755 23663 12774 23697
rect 12827 23663 12842 23697
rect 12899 23663 12910 23697
rect 12971 23663 12978 23697
rect 13043 23663 13046 23697
rect 13080 23663 13081 23697
rect 13148 23663 13153 23697
rect 13216 23663 13225 23697
rect 13284 23663 13297 23697
rect 4298 23554 4335 23588
rect 4369 23554 4403 23588
rect 4437 23554 4471 23588
rect 4505 23554 4539 23588
rect 4573 23554 4607 23588
rect 4641 23554 4675 23588
rect 4709 23554 4743 23588
rect 4777 23554 4811 23588
rect 4845 23554 4879 23588
rect 4913 23554 4947 23588
rect 4981 23554 5015 23588
rect 5049 23554 5083 23588
rect 5117 23554 5151 23588
rect 5185 23554 5219 23588
rect 5253 23554 5287 23588
rect 5321 23554 5355 23588
rect 5389 23554 5423 23588
rect 5457 23554 5491 23588
rect 5525 23554 5559 23588
rect 5593 23554 5627 23588
rect 5661 23554 5695 23588
rect 5729 23554 5763 23588
rect 5797 23554 5831 23588
rect 5865 23554 5899 23588
rect 5933 23554 5967 23588
rect 6001 23554 6035 23588
rect 6069 23554 6103 23588
rect 6137 23554 6171 23588
rect 6205 23554 6239 23588
rect 6273 23554 6307 23588
rect 6341 23554 6375 23588
rect 6409 23554 6443 23588
rect 6477 23554 6511 23588
rect 6545 23554 6579 23588
rect 6613 23554 6647 23588
rect 6681 23554 6715 23588
rect 6749 23554 6783 23588
rect 6817 23554 6851 23588
rect 6885 23554 6919 23588
rect 6953 23554 6987 23588
rect 7021 23554 7055 23588
rect 7089 23554 7123 23588
rect 7157 23554 7191 23588
rect 7225 23554 7259 23588
rect 7293 23554 7327 23588
rect 7361 23554 7395 23588
rect 7429 23554 7463 23588
rect 7497 23554 7531 23588
rect 7565 23554 7599 23588
rect 7633 23554 7667 23588
rect 7701 23554 7735 23588
rect 7769 23554 7803 23588
rect 7837 23554 7871 23588
rect 7905 23554 7939 23588
rect 7973 23554 8007 23588
rect 8041 23554 8075 23588
rect 8109 23554 8143 23588
rect 8177 23554 8211 23588
rect 8245 23554 8279 23588
rect 8313 23554 8347 23588
rect 8381 23554 8415 23588
rect 8449 23554 8483 23588
rect 8517 23554 8551 23588
rect 8585 23554 8619 23588
rect 8653 23554 8687 23588
rect 8721 23554 8755 23588
rect 8789 23554 8823 23588
rect 8857 23554 8891 23588
rect 8925 23554 8959 23588
rect 8993 23554 9027 23588
rect 9061 23554 9095 23588
rect 9129 23554 9163 23588
rect 9197 23554 9231 23588
rect 9265 23554 9299 23588
rect 9333 23554 9367 23588
rect 9401 23554 9435 23588
rect 9469 23554 9503 23588
rect 9537 23554 9571 23588
rect 9605 23554 9639 23588
rect 9673 23554 9707 23588
rect 9741 23554 9775 23588
rect 9809 23554 9843 23588
rect 9877 23554 9911 23588
rect 9945 23554 9979 23588
rect 10013 23554 10047 23588
rect 10081 23554 10115 23588
rect 10149 23554 10183 23588
rect 10217 23554 10251 23588
rect 10285 23554 10319 23588
rect 10353 23554 10387 23588
rect 10421 23554 10455 23588
rect 10489 23554 10523 23588
rect 10557 23554 10591 23588
rect 10625 23554 10659 23588
rect 10693 23554 10727 23588
rect 10761 23554 10795 23588
rect 10829 23554 10863 23588
rect 10897 23554 10931 23588
rect 10965 23554 10999 23588
rect 11033 23554 11067 23588
rect 11101 23554 11135 23588
rect 11169 23554 11203 23588
rect 11237 23554 11271 23588
rect 11305 23554 11339 23588
rect 11373 23554 11407 23588
rect 11441 23554 11475 23588
rect 11509 23554 11543 23588
rect 11577 23554 11611 23588
rect 11645 23554 11679 23588
rect 11713 23554 11747 23588
rect 11781 23554 11815 23588
rect 11849 23554 11883 23588
rect 11917 23554 11951 23588
rect 11985 23554 12019 23588
rect 12053 23554 12087 23588
rect 12121 23554 12155 23588
rect 12189 23554 12223 23588
rect 12257 23554 12291 23588
rect 12325 23554 12359 23588
rect 12393 23554 12427 23588
rect 12461 23554 12495 23588
rect 12529 23554 12563 23588
rect 12597 23554 12631 23588
rect 12665 23554 12699 23588
rect 12733 23554 12767 23588
rect 12801 23554 12835 23588
rect 12869 23554 12903 23588
rect 12937 23554 12971 23588
rect 13005 23554 13039 23588
rect 13073 23554 13107 23588
rect 13141 23554 13175 23588
rect 13209 23554 13243 23588
rect 13277 23554 13311 23588
rect 13345 23554 13379 23588
rect 13413 23554 13447 23588
rect 13481 23554 13515 23588
rect 4934 23428 4954 23462
rect 4988 23428 5022 23462
rect 5056 23428 5081 23462
rect 5124 23428 5154 23462
rect 5192 23428 5226 23462
rect 5261 23428 5294 23462
rect 5334 23428 5362 23462
rect 5407 23428 5430 23462
rect 5480 23428 5498 23462
rect 5553 23428 5566 23462
rect 5626 23428 5634 23462
rect 5699 23428 5702 23462
rect 5736 23428 5737 23462
rect 5804 23428 5809 23462
rect 5872 23428 5881 23462
rect 5940 23428 5953 23462
rect 6008 23428 6025 23462
rect 6076 23428 6097 23462
rect 6144 23428 6169 23462
rect 6212 23428 6241 23462
rect 6280 23428 6313 23462
rect 6348 23428 6382 23462
rect 6419 23428 6450 23462
rect 6491 23428 6518 23462
rect 6563 23428 6586 23462
rect 6635 23428 6654 23462
rect 6707 23428 6722 23462
rect 6779 23428 6790 23462
rect 6851 23428 6858 23462
rect 6923 23428 6926 23462
rect 6960 23428 6961 23462
rect 7028 23428 7033 23462
rect 7096 23428 7105 23462
rect 7164 23428 7177 23462
rect 7232 23428 7249 23462
rect 7300 23428 7321 23462
rect 7368 23428 7393 23462
rect 7436 23428 7465 23462
rect 7504 23428 7537 23462
rect 7572 23428 7606 23462
rect 7643 23428 7674 23462
rect 7715 23428 7742 23462
rect 7787 23428 7810 23462
rect 7859 23428 7878 23462
rect 7931 23428 7946 23462
rect 8003 23428 8014 23462
rect 8075 23428 8082 23462
rect 8147 23428 8150 23462
rect 8184 23428 8185 23462
rect 8252 23428 8257 23462
rect 8320 23428 8329 23462
rect 8388 23428 8401 23462
rect 8456 23428 8473 23462
rect 8524 23428 8545 23462
rect 8592 23428 8617 23462
rect 8660 23428 8689 23462
rect 8728 23428 8761 23462
rect 8796 23428 8830 23462
rect 8867 23428 8898 23462
rect 8939 23428 8966 23462
rect 9011 23428 9034 23462
rect 9083 23428 9102 23462
rect 9155 23428 9170 23462
rect 9227 23428 9238 23462
rect 9299 23428 9306 23462
rect 9371 23428 9374 23462
rect 9408 23428 9409 23462
rect 9476 23428 9481 23462
rect 9544 23428 9553 23462
rect 9612 23428 9625 23462
rect 9680 23428 9697 23462
rect 9748 23428 9769 23462
rect 9816 23428 9841 23462
rect 9884 23428 9913 23462
rect 9952 23428 9985 23462
rect 10020 23428 10054 23462
rect 10091 23428 10122 23462
rect 10163 23428 10190 23462
rect 10235 23428 10258 23462
rect 10307 23428 10326 23462
rect 10379 23428 10394 23462
rect 10451 23428 10462 23462
rect 10523 23428 10530 23462
rect 10595 23428 10598 23462
rect 10632 23428 10633 23462
rect 10700 23428 10705 23462
rect 10768 23428 10777 23462
rect 10836 23428 10849 23462
rect 10904 23428 10921 23462
rect 10972 23428 10993 23462
rect 11040 23428 11065 23462
rect 11108 23428 11137 23462
rect 11176 23428 11209 23462
rect 11244 23428 11278 23462
rect 11315 23428 11346 23462
rect 11387 23428 11414 23462
rect 11459 23428 11482 23462
rect 11531 23428 11550 23462
rect 11603 23428 11618 23462
rect 11675 23428 11686 23462
rect 11747 23428 11754 23462
rect 11819 23428 11822 23462
rect 11856 23428 11857 23462
rect 11924 23428 11929 23462
rect 11992 23428 12001 23462
rect 12060 23428 12073 23462
rect 12128 23428 12145 23462
rect 12196 23428 12217 23462
rect 12264 23428 12289 23462
rect 12332 23428 12361 23462
rect 12400 23428 12433 23462
rect 12468 23428 12502 23462
rect 12539 23428 12570 23462
rect 12611 23428 12638 23462
rect 12683 23428 12706 23462
rect 12755 23428 12774 23462
rect 12827 23428 12842 23462
rect 12899 23428 12910 23462
rect 12971 23428 12978 23462
rect 13043 23428 13046 23462
rect 13080 23428 13081 23462
rect 13148 23428 13153 23462
rect 13216 23428 13225 23462
rect 13284 23428 13297 23462
rect 4761 23076 4809 23334
rect 4727 23037 4809 23076
rect 4761 23003 4809 23037
rect 4727 22964 4809 23003
rect 4761 22930 4809 22964
rect 4727 22891 4809 22930
rect 4761 22857 4809 22891
rect 4727 22818 4809 22857
rect 4761 22784 4809 22818
rect 4727 22745 4809 22784
rect 4761 22711 4809 22745
rect 4727 22672 4809 22711
rect 4761 22638 4809 22672
rect 4727 22599 4809 22638
rect 4761 22565 4809 22599
rect 4727 22526 4809 22565
rect 4761 22492 4809 22526
rect 4727 22453 4809 22492
rect 4761 22419 4809 22453
rect 4727 22380 4809 22419
rect 4761 22346 4809 22380
rect 4727 22306 4809 22346
rect 4761 22272 4809 22306
rect 4727 22232 4809 22272
rect 4761 22198 4809 22232
rect 4727 22158 4809 22198
rect 4761 22124 4809 22158
rect 4727 22084 4809 22124
rect 5073 22993 5107 23032
rect 5073 22920 5107 22959
rect 5073 22847 5107 22886
rect 5073 22774 5107 22813
rect 5073 22701 5107 22740
rect 5073 22628 5107 22667
rect 5073 22556 5107 22594
rect 5073 22484 5107 22522
rect 5073 22412 5107 22450
rect 5073 22340 5107 22378
rect 5073 22268 5107 22306
rect 5073 22196 5107 22234
rect 5073 22124 5107 22162
rect 6718 22976 6752 23020
rect 6718 22898 6752 22942
rect 6718 22820 6752 22864
rect 6718 22742 6752 22786
rect 6718 22664 6752 22708
rect 6718 22586 6752 22630
rect 6718 22509 6752 22552
rect 6718 22432 6752 22475
rect 6718 22355 6752 22398
rect 6718 22278 6752 22321
rect 6718 22201 6752 22244
rect 6718 22124 6752 22167
rect 8374 22976 8408 23020
rect 8374 22898 8408 22942
rect 8374 22820 8408 22864
rect 8374 22742 8408 22786
rect 8374 22664 8408 22708
rect 8374 22586 8408 22630
rect 8374 22509 8408 22552
rect 8374 22432 8408 22475
rect 8374 22355 8408 22398
rect 8374 22278 8408 22321
rect 8374 22201 8408 22244
rect 8374 22124 8408 22167
rect 10030 22976 10064 23020
rect 10030 22898 10064 22942
rect 10030 22820 10064 22864
rect 10030 22742 10064 22786
rect 10030 22664 10064 22708
rect 10030 22586 10064 22630
rect 10030 22509 10064 22552
rect 10030 22432 10064 22475
rect 10030 22355 10064 22398
rect 10030 22278 10064 22321
rect 10030 22201 10064 22244
rect 10030 22124 10064 22167
rect 11686 22976 11720 23020
rect 11686 22898 11720 22942
rect 11686 22820 11720 22864
rect 11686 22742 11720 22786
rect 11686 22664 11720 22708
rect 11686 22586 11720 22630
rect 11686 22509 11720 22552
rect 11686 22432 11720 22475
rect 11686 22355 11720 22398
rect 11686 22278 11720 22321
rect 11686 22201 11720 22244
rect 11686 22124 11720 22167
rect 13342 22976 13376 23020
rect 13342 22898 13376 22942
rect 13342 22820 13376 22864
rect 13342 22742 13376 22786
rect 13342 22664 13376 22708
rect 13342 22586 13376 22630
rect 13342 22509 13376 22552
rect 13342 22432 13376 22475
rect 13342 22355 13376 22398
rect 13342 22278 13376 22321
rect 13342 22201 13376 22244
rect 13342 22124 13376 22167
rect 13617 22178 13699 22217
rect 13627 22144 13665 22178
rect 13617 22105 13699 22144
rect 4761 22050 4809 22084
rect 4727 22010 4809 22050
rect 4761 21976 4809 22010
rect 13627 22071 13665 22105
rect 13617 22032 13699 22071
rect 13627 21998 13665 22032
rect 13617 21959 13699 21998
rect 13627 21925 13665 21959
rect 4298 21855 4335 21889
rect 4369 21855 4403 21889
rect 4437 21855 4471 21889
rect 4505 21855 4539 21889
rect 4573 21855 4607 21889
rect 4641 21855 4675 21889
rect 4709 21855 4743 21889
rect 4777 21855 4811 21889
rect 4845 21855 4879 21889
rect 4913 21855 4947 21889
rect 4981 21855 5015 21889
rect 5049 21855 5083 21889
rect 5117 21855 5151 21889
rect 5185 21855 5219 21889
rect 5253 21855 5287 21889
rect 5321 21855 5355 21889
rect 5389 21855 5423 21889
rect 5457 21855 5491 21889
rect 5525 21855 5559 21889
rect 5593 21855 5627 21889
rect 5661 21855 5695 21889
rect 5729 21855 5763 21889
rect 5797 21855 5831 21889
rect 5865 21855 5899 21889
rect 5933 21855 5967 21889
rect 6001 21855 6035 21889
rect 6069 21855 6103 21889
rect 6137 21855 6171 21889
rect 6205 21855 6239 21889
rect 6273 21855 6307 21889
rect 6341 21855 6375 21889
rect 6409 21855 6443 21889
rect 6477 21855 6511 21889
rect 6545 21855 6579 21889
rect 6613 21855 6647 21889
rect 6681 21855 6715 21889
rect 6749 21855 6783 21889
rect 6817 21855 6851 21889
rect 6885 21855 6919 21889
rect 6953 21855 6987 21889
rect 7021 21855 7055 21889
rect 7089 21855 7123 21889
rect 7157 21855 7191 21889
rect 7225 21855 7259 21889
rect 7293 21855 7327 21889
rect 7361 21855 7395 21889
rect 7429 21855 7463 21889
rect 7497 21855 7531 21889
rect 7565 21855 7599 21889
rect 7633 21855 7667 21889
rect 7701 21855 7735 21889
rect 7769 21855 7803 21889
rect 7837 21855 7871 21889
rect 7905 21855 7939 21889
rect 7973 21855 8007 21889
rect 8041 21855 8075 21889
rect 8109 21855 8143 21889
rect 8177 21855 8211 21889
rect 8245 21855 8279 21889
rect 8313 21855 8347 21889
rect 8381 21855 8415 21889
rect 8449 21855 8483 21889
rect 8517 21855 8551 21889
rect 8585 21855 8619 21889
rect 8653 21855 8687 21889
rect 8721 21855 8755 21889
rect 8789 21855 8823 21889
rect 8857 21855 8891 21889
rect 8925 21855 8959 21889
rect 8993 21855 9027 21889
rect 9061 21855 9095 21889
rect 9129 21855 9163 21889
rect 9197 21855 9231 21889
rect 9265 21855 9299 21889
rect 9333 21855 9367 21889
rect 9401 21855 9435 21889
rect 9469 21855 9503 21889
rect 9537 21855 9571 21889
rect 9605 21855 9639 21889
rect 9673 21855 9707 21889
rect 9741 21855 9775 21889
rect 9809 21855 9843 21889
rect 9877 21855 9911 21889
rect 9945 21855 9979 21889
rect 10013 21855 10047 21889
rect 10081 21855 10115 21889
rect 10149 21855 10183 21889
rect 10217 21855 10251 21889
rect 10285 21855 10319 21889
rect 10353 21855 10387 21889
rect 10421 21855 10455 21889
rect 10489 21855 10523 21889
rect 10557 21855 10591 21889
rect 10625 21855 10659 21889
rect 10693 21855 10727 21889
rect 10761 21855 10795 21889
rect 10829 21855 10863 21889
rect 10897 21855 10931 21889
rect 10965 21855 10999 21889
rect 11033 21855 11067 21889
rect 11101 21855 11135 21889
rect 11169 21855 11203 21889
rect 11237 21855 11271 21889
rect 11305 21855 11339 21889
rect 11373 21855 11407 21889
rect 11441 21855 11475 21889
rect 11509 21855 11543 21889
rect 11577 21855 11611 21889
rect 11645 21855 11679 21889
rect 11713 21855 11747 21889
rect 11781 21855 11815 21889
rect 11849 21855 11883 21889
rect 11917 21855 11951 21889
rect 11985 21855 12019 21889
rect 12053 21855 12087 21889
rect 12121 21855 12155 21889
rect 12189 21855 12223 21889
rect 12257 21855 12291 21889
rect 12325 21855 12359 21889
rect 12393 21855 12427 21889
rect 12461 21855 12495 21889
rect 12529 21855 12563 21889
rect 12597 21855 12631 21889
rect 12665 21855 12699 21889
rect 12733 21855 12767 21889
rect 12801 21855 12835 21889
rect 12869 21855 12903 21889
rect 12937 21855 12971 21889
rect 13005 21855 13039 21889
rect 13073 21855 13107 21889
rect 13141 21855 13175 21889
rect 13209 21855 13243 21889
rect 13277 21855 13311 21889
rect 13345 21855 13379 21889
rect 13413 21855 13447 21889
rect 13481 21855 13515 21889
rect 13617 21886 13699 21925
rect 13627 21852 13665 21886
rect 13617 21813 13699 21852
rect 13627 21779 13665 21813
rect 4934 21729 4954 21763
rect 4988 21729 5022 21763
rect 5056 21729 5079 21763
rect 5124 21729 5152 21763
rect 5192 21729 5225 21763
rect 5260 21729 5294 21763
rect 5332 21729 5362 21763
rect 5405 21729 5430 21763
rect 5478 21729 5498 21763
rect 5551 21729 5566 21763
rect 5624 21729 5634 21763
rect 5697 21729 5702 21763
rect 5804 21729 5809 21763
rect 5872 21729 5881 21763
rect 5940 21729 5953 21763
rect 6008 21729 6025 21763
rect 6076 21729 6097 21763
rect 6144 21729 6169 21763
rect 6212 21729 6241 21763
rect 6280 21729 6313 21763
rect 6348 21729 6382 21763
rect 6419 21729 6450 21763
rect 6491 21729 6518 21763
rect 6563 21729 6586 21763
rect 6635 21729 6654 21763
rect 6707 21729 6722 21763
rect 6779 21729 6790 21763
rect 6851 21729 6858 21763
rect 6923 21729 6926 21763
rect 6960 21729 6961 21763
rect 7028 21729 7033 21763
rect 7096 21729 7105 21763
rect 7164 21729 7177 21763
rect 7232 21729 7249 21763
rect 7300 21729 7321 21763
rect 7368 21729 7393 21763
rect 7436 21729 7465 21763
rect 7504 21729 7537 21763
rect 7572 21729 7606 21763
rect 7643 21729 7674 21763
rect 7715 21729 7742 21763
rect 7787 21729 7810 21763
rect 7859 21729 7878 21763
rect 7931 21729 7946 21763
rect 8003 21729 8014 21763
rect 8075 21729 8082 21763
rect 8147 21729 8150 21763
rect 8184 21729 8185 21763
rect 8252 21729 8257 21763
rect 8320 21729 8329 21763
rect 8388 21729 8401 21763
rect 8456 21729 8473 21763
rect 8524 21729 8545 21763
rect 8592 21729 8617 21763
rect 8660 21729 8689 21763
rect 8728 21729 8761 21763
rect 8796 21729 8830 21763
rect 8867 21729 8898 21763
rect 8939 21729 8966 21763
rect 9011 21729 9034 21763
rect 9083 21729 9102 21763
rect 9155 21729 9170 21763
rect 9227 21729 9238 21763
rect 9299 21729 9306 21763
rect 9371 21729 9374 21763
rect 9408 21729 9409 21763
rect 9476 21729 9481 21763
rect 9544 21729 9553 21763
rect 9612 21729 9625 21763
rect 9680 21729 9697 21763
rect 9748 21729 9769 21763
rect 9816 21729 9841 21763
rect 9884 21729 9913 21763
rect 9952 21729 9985 21763
rect 10020 21729 10054 21763
rect 10091 21729 10122 21763
rect 10163 21729 10190 21763
rect 10235 21729 10258 21763
rect 10307 21729 10326 21763
rect 10379 21729 10394 21763
rect 10451 21729 10462 21763
rect 10523 21729 10530 21763
rect 10595 21729 10598 21763
rect 10632 21729 10633 21763
rect 10700 21729 10705 21763
rect 10768 21729 10777 21763
rect 10836 21729 10849 21763
rect 10904 21729 10921 21763
rect 10972 21729 10993 21763
rect 11040 21729 11065 21763
rect 11108 21729 11137 21763
rect 11176 21729 11209 21763
rect 11244 21729 11278 21763
rect 11315 21729 11346 21763
rect 11387 21729 11414 21763
rect 11459 21729 11482 21763
rect 11531 21729 11550 21763
rect 11603 21729 11618 21763
rect 11675 21729 11686 21763
rect 11747 21729 11754 21763
rect 11819 21729 11822 21763
rect 11856 21729 11857 21763
rect 11924 21729 11929 21763
rect 11992 21729 12001 21763
rect 12060 21729 12073 21763
rect 12128 21729 12145 21763
rect 12196 21729 12217 21763
rect 12264 21729 12289 21763
rect 12332 21729 12361 21763
rect 12400 21729 12433 21763
rect 12468 21729 12502 21763
rect 12539 21729 12570 21763
rect 12611 21729 12638 21763
rect 12683 21729 12706 21763
rect 12755 21729 12774 21763
rect 12827 21729 12842 21763
rect 12899 21729 12910 21763
rect 12971 21729 12978 21763
rect 13043 21729 13046 21763
rect 13080 21729 13081 21763
rect 13148 21729 13153 21763
rect 13216 21729 13225 21763
rect 13284 21729 13297 21763
rect 13617 21740 13699 21779
rect 13627 21706 13665 21740
rect 13617 21667 13699 21706
rect 4761 21601 4809 21635
rect 4727 21561 4809 21601
rect 4761 21527 4809 21561
rect 4727 21487 4809 21527
rect 4761 21453 4809 21487
rect 4727 21413 4809 21453
rect 4761 21379 4809 21413
rect 4727 21339 4809 21379
rect 4761 21305 4809 21339
rect 4727 21265 4809 21305
rect 4761 21231 4809 21265
rect 13627 21633 13665 21667
rect 13617 21594 13699 21633
rect 13627 21560 13665 21594
rect 13617 21521 13699 21560
rect 13627 21487 13665 21521
rect 13617 21448 13699 21487
rect 13627 21414 13665 21448
rect 13617 21375 13699 21414
rect 13627 21341 13665 21375
rect 13617 21302 13699 21341
rect 13627 21268 13665 21302
rect 4727 21191 4809 21231
rect 4761 21157 4809 21191
rect 4727 21117 4809 21157
rect 4761 21083 4809 21117
rect 4727 21043 4809 21083
rect 4761 21009 4809 21043
rect 4727 20969 4809 21009
rect 4761 20935 4809 20969
rect 4727 20895 4809 20935
rect 4761 20861 4809 20895
rect 4727 20822 4809 20861
rect 4761 20788 4809 20822
rect 4727 20749 4809 20788
rect 4761 20715 4809 20749
rect 4727 20676 4809 20715
rect 4761 20642 4809 20676
rect 4727 20603 4809 20642
rect 4761 20569 4809 20603
rect 4727 20530 4809 20569
rect 4761 20496 4809 20530
rect 4727 20457 4809 20496
rect 4761 20423 4809 20457
rect 4727 20384 4809 20423
rect 4761 20350 4809 20384
rect 4727 20311 4809 20350
rect 4761 20277 4809 20311
rect 5073 21178 5107 21217
rect 5073 21105 5107 21144
rect 5073 21032 5107 21071
rect 5073 20959 5107 20998
rect 5073 20887 5107 20925
rect 5073 20815 5107 20853
rect 5073 20743 5107 20781
rect 5073 20671 5107 20709
rect 5073 20599 5107 20637
rect 5073 20527 5107 20565
rect 5073 20455 5107 20493
rect 5073 20383 5107 20421
rect 5073 20311 5107 20349
rect 6718 21178 6752 21217
rect 6718 21105 6752 21144
rect 6718 21032 6752 21071
rect 6718 20959 6752 20998
rect 6718 20887 6752 20925
rect 6718 20815 6752 20853
rect 6718 20743 6752 20781
rect 6718 20671 6752 20709
rect 6718 20599 6752 20637
rect 6718 20527 6752 20565
rect 6718 20455 6752 20493
rect 6718 20383 6752 20421
rect 6718 20311 6752 20349
rect 8374 21178 8408 21217
rect 8374 21105 8408 21144
rect 8374 21032 8408 21071
rect 8374 20959 8408 20998
rect 8374 20887 8408 20925
rect 8374 20815 8408 20853
rect 8374 20743 8408 20781
rect 8374 20671 8408 20709
rect 8374 20599 8408 20637
rect 8374 20527 8408 20565
rect 8374 20455 8408 20493
rect 8374 20383 8408 20421
rect 8374 20311 8408 20349
rect 10030 21178 10064 21217
rect 10030 21105 10064 21144
rect 10030 21032 10064 21071
rect 10030 20959 10064 20998
rect 10030 20887 10064 20925
rect 10030 20815 10064 20853
rect 10030 20743 10064 20781
rect 10030 20671 10064 20709
rect 10030 20599 10064 20637
rect 10030 20527 10064 20565
rect 10030 20455 10064 20493
rect 10030 20383 10064 20421
rect 10030 20311 10064 20349
rect 11686 21178 11720 21217
rect 11686 21105 11720 21144
rect 11686 21032 11720 21071
rect 11686 20959 11720 20998
rect 11686 20887 11720 20925
rect 11686 20815 11720 20853
rect 11686 20743 11720 20781
rect 11686 20671 11720 20709
rect 11686 20599 11720 20637
rect 11686 20527 11720 20565
rect 11686 20455 11720 20493
rect 11686 20383 11720 20421
rect 11686 20311 11720 20349
rect 13342 21178 13376 21217
rect 13342 21105 13376 21144
rect 13342 21032 13376 21071
rect 13342 20959 13376 20998
rect 13342 20887 13376 20925
rect 13342 20815 13376 20853
rect 13342 20743 13376 20781
rect 13342 20671 13376 20709
rect 13342 20599 13376 20637
rect 13342 20527 13376 20565
rect 13342 20455 13376 20493
rect 13342 20383 13376 20421
rect 13342 20311 13376 20349
rect 13617 21229 13699 21268
rect 13627 21195 13665 21229
rect 13617 21156 13699 21195
rect 13627 21122 13665 21156
rect 13617 21083 13699 21122
rect 13627 21049 13665 21083
rect 13617 21010 13699 21049
rect 13627 20976 13665 21010
rect 13617 20937 13699 20976
rect 13627 20903 13665 20937
rect 13617 20864 13699 20903
rect 13627 20830 13665 20864
rect 13617 20791 13699 20830
rect 13627 20757 13665 20791
rect 13617 20718 13699 20757
rect 13627 20684 13665 20718
rect 13617 20645 13699 20684
rect 13627 20611 13665 20645
rect 13617 20572 13699 20611
rect 13627 20538 13665 20572
rect 13617 20531 13699 20538
rect 13515 20499 13699 20531
rect 13515 20496 13521 20499
rect 13555 20496 13593 20499
rect 13555 20465 13583 20496
rect 13627 20465 13665 20499
rect 13549 20462 13583 20465
rect 13617 20462 13699 20465
rect 13515 20427 13699 20462
rect 13549 20426 13583 20427
rect 13617 20426 13699 20427
rect 13555 20393 13583 20426
rect 13515 20392 13521 20393
rect 13555 20392 13593 20393
rect 13627 20392 13665 20426
rect 13515 20358 13699 20392
rect 13549 20353 13583 20358
rect 13617 20353 13699 20358
rect 13555 20324 13583 20353
rect 13515 20319 13521 20324
rect 13555 20319 13593 20324
rect 13627 20319 13665 20353
rect 13515 20289 13699 20319
rect 13549 20280 13583 20289
rect 13617 20280 13699 20289
rect 4128 20207 4298 20257
rect 13555 20255 13583 20280
rect 13515 20246 13521 20255
rect 13555 20246 13593 20255
rect 13627 20246 13665 20280
rect 13515 20207 13699 20246
rect 4128 20173 4152 20207
rect 4186 20173 4221 20207
rect 4255 20173 4290 20207
rect 4324 20173 4359 20207
rect 4393 20173 4428 20207
rect 4462 20173 4497 20207
rect 4531 20173 4566 20207
rect 4600 20173 4635 20207
rect 4669 20173 4704 20207
rect 4738 20173 4773 20207
rect 4807 20173 4842 20207
rect 4876 20173 4911 20207
rect 4945 20173 4980 20207
rect 5014 20173 5049 20207
rect 5083 20173 5118 20207
rect 5152 20173 5187 20207
rect 5221 20173 5256 20207
rect 5290 20173 5325 20207
rect 5359 20173 5394 20207
rect 5428 20173 5463 20207
rect 5497 20173 5532 20207
rect 5566 20173 5601 20207
rect 5635 20173 5670 20207
rect 5704 20173 5739 20207
rect 5773 20173 5807 20207
rect 5841 20173 5875 20207
rect 5909 20173 5943 20207
rect 5977 20173 6011 20207
rect 6045 20173 6079 20207
rect 6113 20173 6147 20207
rect 6181 20173 6215 20207
rect 6249 20173 6283 20207
rect 6317 20173 6351 20207
rect 6385 20173 6419 20207
rect 6453 20173 6487 20207
rect 6521 20173 6555 20207
rect 6589 20173 6623 20207
rect 6657 20173 6691 20207
rect 6725 20173 6759 20207
rect 6793 20173 6827 20207
rect 6861 20173 6895 20207
rect 6929 20173 6963 20207
rect 6997 20173 7031 20207
rect 7065 20173 7099 20207
rect 7133 20173 7167 20207
rect 7201 20173 7235 20207
rect 7269 20173 7303 20207
rect 7337 20173 7371 20207
rect 7405 20173 7439 20207
rect 7473 20173 7507 20207
rect 7541 20173 7575 20207
rect 7609 20173 7643 20207
rect 7677 20173 7711 20207
rect 7745 20173 7779 20207
rect 7813 20173 7847 20207
rect 7881 20173 7915 20207
rect 7949 20173 7983 20207
rect 8017 20173 8051 20207
rect 8085 20173 8119 20207
rect 8153 20173 8187 20207
rect 8221 20173 8255 20207
rect 8289 20173 8323 20207
rect 8357 20173 8391 20207
rect 8425 20173 8459 20207
rect 8493 20173 8527 20207
rect 8561 20173 8595 20207
rect 8629 20173 8663 20207
rect 8697 20173 8731 20207
rect 8765 20173 8799 20207
rect 8833 20173 8867 20207
rect 8901 20173 8935 20207
rect 8969 20173 9003 20207
rect 9037 20173 9071 20207
rect 9105 20173 9139 20207
rect 9173 20173 9207 20207
rect 9241 20173 9275 20207
rect 9309 20173 9343 20207
rect 9377 20173 9411 20207
rect 9445 20173 9479 20207
rect 9513 20173 9547 20207
rect 9581 20173 9615 20207
rect 9649 20173 9683 20207
rect 9717 20173 9751 20207
rect 9785 20173 9819 20207
rect 9853 20173 9887 20207
rect 9921 20173 9955 20207
rect 9989 20173 10023 20207
rect 10057 20173 10091 20207
rect 10125 20173 10159 20207
rect 10193 20173 10227 20207
rect 10261 20173 10295 20207
rect 10329 20173 10363 20207
rect 10397 20173 10431 20207
rect 10465 20173 10499 20207
rect 10533 20173 10567 20207
rect 10601 20173 10635 20207
rect 10669 20173 10703 20207
rect 10737 20173 10771 20207
rect 10805 20173 10839 20207
rect 10873 20173 10907 20207
rect 10941 20173 10975 20207
rect 11009 20173 11043 20207
rect 11077 20173 11111 20207
rect 11145 20173 11179 20207
rect 11213 20173 11247 20207
rect 11281 20173 11315 20207
rect 11349 20173 11383 20207
rect 11417 20173 11451 20207
rect 11485 20173 11519 20207
rect 11553 20173 11587 20207
rect 11621 20173 11655 20207
rect 11689 20173 11723 20207
rect 11757 20173 11791 20207
rect 11825 20173 11859 20207
rect 11893 20173 11927 20207
rect 11961 20173 11995 20207
rect 12029 20173 12063 20207
rect 12097 20173 12131 20207
rect 12165 20173 12199 20207
rect 12233 20173 12267 20207
rect 12301 20173 12335 20207
rect 12369 20173 12403 20207
rect 12437 20173 12471 20207
rect 12505 20173 12539 20207
rect 12573 20173 12607 20207
rect 12641 20173 12675 20207
rect 12709 20173 12743 20207
rect 12777 20173 12811 20207
rect 12845 20173 12879 20207
rect 12913 20173 12947 20207
rect 12981 20173 13015 20207
rect 13049 20173 13083 20207
rect 13117 20173 13151 20207
rect 13185 20173 13219 20207
rect 13253 20173 13287 20207
rect 13321 20173 13355 20207
rect 13389 20173 13423 20207
rect 13457 20173 13491 20207
rect 13555 20173 13559 20207
rect 13627 20173 13665 20207
rect 13838 26581 13840 26620
rect 13942 26581 13944 26620
rect 13838 26508 13840 26547
rect 13942 26508 13944 26547
rect 13838 26435 13840 26474
rect 13942 26435 13944 26474
rect 13838 26362 13840 26401
rect 13942 26362 13944 26401
rect 13838 26289 13840 26328
rect 13942 26289 13944 26328
rect 13838 26216 13840 26255
rect 13942 26216 13944 26255
rect 13838 26143 13840 26182
rect 13942 26143 13944 26182
rect 13838 26070 13840 26109
rect 13942 26070 13944 26109
rect 13838 25997 13840 26036
rect 13942 25997 13944 26036
rect 13838 25924 13840 25963
rect 13942 25924 13944 25963
rect 13838 25851 13840 25890
rect 13942 25851 13944 25890
rect 13838 25778 13840 25817
rect 13942 25778 13944 25817
rect 13838 25705 13840 25744
rect 13942 25705 13944 25744
rect 13838 25632 13840 25671
rect 13942 25632 13944 25671
rect 13838 25559 13840 25598
rect 13942 25559 13944 25598
rect 13838 25486 13840 25525
rect 13942 25486 13944 25525
rect 13838 25413 13840 25452
rect 13942 25413 13944 25452
rect 13838 25340 13840 25379
rect 13942 25340 13944 25379
rect 13838 25267 13840 25306
rect 13942 25267 13944 25306
rect 13838 25194 13840 25233
rect 13942 25194 13944 25233
rect 13838 25121 13840 25160
rect 13942 25121 13944 25160
rect 13838 25048 13840 25087
rect 13942 25048 13944 25087
rect 13838 24975 13840 25014
rect 13942 24975 13944 25014
rect 13838 24902 13840 24941
rect 13942 24902 13944 24941
rect 13838 24829 13840 24868
rect 13942 24829 13944 24868
rect 13838 24756 13840 24795
rect 13942 24756 13944 24795
rect 13838 24683 13840 24722
rect 13942 24683 13944 24722
rect 13838 24610 13840 24649
rect 13942 24610 13944 24649
rect 13838 24537 13840 24576
rect 13942 24537 13944 24576
rect 13838 24464 13840 24503
rect 13942 24464 13944 24503
rect 13838 24391 13840 24430
rect 13942 24391 13944 24430
rect 13838 24318 13840 24357
rect 13942 24318 13944 24357
rect 13838 24245 13840 24284
rect 13942 24245 13944 24284
rect 13838 24172 13840 24211
rect 13942 24172 13944 24211
rect 13838 24099 13840 24138
rect 13942 24099 13944 24138
rect 13838 24026 13840 24065
rect 13942 24026 13944 24065
rect 13838 23953 13840 23992
rect 13942 23953 13944 23992
rect 13838 23880 13840 23919
rect 13942 23880 13944 23919
rect 13838 23807 13840 23846
rect 13942 23807 13944 23846
rect 13838 23734 13840 23773
rect 13942 23734 13944 23773
rect 13838 23661 13840 23700
rect 13942 23661 13944 23700
rect 13838 23588 13840 23627
rect 13942 23588 13944 23627
rect 13838 23515 13840 23554
rect 13942 23515 13944 23554
rect 13838 23442 13840 23481
rect 13942 23442 13944 23481
rect 13838 23369 13840 23408
rect 13942 23369 13944 23408
rect 13838 23296 13840 23335
rect 13942 23296 13944 23335
rect 13838 23223 13840 23262
rect 13942 23223 13944 23262
rect 13838 23150 13840 23189
rect 13942 23150 13944 23189
rect 13838 23077 13840 23116
rect 13942 23077 13944 23116
rect 13838 23004 13840 23043
rect 13942 23004 13944 23043
rect 13838 22931 13840 22970
rect 13942 22931 13944 22970
rect 13838 22858 13840 22897
rect 13942 22858 13944 22897
rect 13838 22785 13840 22824
rect 13942 22785 13944 22824
rect 13838 22712 13840 22751
rect 13942 22712 13944 22751
rect 13838 22639 13840 22678
rect 13942 22639 13944 22678
rect 13838 22566 13840 22605
rect 13942 22566 13944 22605
rect 13838 22493 13840 22532
rect 13942 22493 13944 22532
rect 13838 22420 13840 22459
rect 13942 22420 13944 22459
rect 13838 22347 13840 22386
rect 13942 22347 13944 22386
rect 13838 22274 13840 22313
rect 13942 22274 13944 22313
rect 13838 22201 13840 22240
rect 13942 22201 13944 22240
rect 13838 22128 13840 22167
rect 13942 22128 13944 22167
rect 13838 22055 13840 22094
rect 13942 22055 13944 22094
rect 13838 21982 13840 22021
rect 13942 21982 13944 22021
rect 13838 21909 13840 21948
rect 13942 21909 13944 21948
rect 13838 21836 13840 21875
rect 13942 21836 13944 21875
rect 13838 21763 13840 21802
rect 13942 21763 13944 21802
rect 13838 21690 13840 21729
rect 13942 21690 13944 21729
rect 13838 21617 13840 21656
rect 13942 21617 13944 21656
rect 13838 21544 13840 21583
rect 13942 21544 13944 21583
rect 13838 21471 13840 21510
rect 13942 21471 13944 21510
rect 13838 21329 13840 21437
rect 13942 21329 13944 21437
rect 1837 19443 1943 19477
rect 2049 19443 2056 19477
rect 1837 19403 1946 19443
rect 2048 19403 2056 19443
rect 1837 19369 1943 19403
rect 2049 19369 2056 19403
rect 1837 19329 1946 19369
rect 2048 19329 2056 19369
rect 1837 19295 1943 19329
rect 2049 19295 2056 19329
rect 1837 19255 1946 19295
rect 2048 19255 2056 19295
rect 1837 19221 1943 19255
rect 2049 19221 2056 19255
rect 1837 19181 1946 19221
rect 2048 19181 2056 19221
rect 1837 19147 1943 19181
rect 2049 19147 2056 19181
rect 1837 19107 1946 19147
rect 2048 19107 2056 19147
rect 1837 19073 1943 19107
rect 2049 19073 2056 19107
rect 1837 19033 1946 19073
rect 2048 19033 2056 19073
rect 1837 18999 1943 19033
rect 2049 18999 2056 19033
rect 1837 18959 1946 18999
rect 2048 18959 2056 18999
rect 1837 18925 1943 18959
rect 2049 18925 2056 18959
rect 1837 18884 1946 18925
rect 2048 18884 2056 18925
rect 1837 18850 1943 18884
rect 2049 18850 2056 18884
rect 1837 18809 1946 18850
rect 2048 18809 2056 18850
rect 1837 18775 1943 18809
rect 2049 18775 2056 18809
rect 1837 18734 1946 18775
rect 2048 18734 2056 18775
rect 1837 18700 1943 18734
rect 2049 18700 2056 18734
rect 1837 18659 1946 18700
rect 2048 18659 2056 18700
rect 1837 18625 1943 18659
rect 2049 18625 2056 18659
rect 1837 18584 1946 18625
rect 2048 18584 2056 18625
rect 1837 18550 1943 18584
rect 2049 18550 2056 18584
rect 1837 18509 1946 18550
rect 2048 18509 2056 18550
rect 1837 18475 1943 18509
rect 2049 18475 2056 18509
rect 1837 18434 1946 18475
rect 2048 18434 2056 18475
rect 1837 18400 1943 18434
rect 2049 18400 2056 18434
rect 1837 18359 1946 18400
rect 2048 18359 2056 18400
rect 1837 18325 1943 18359
rect 2049 18325 2056 18359
rect 1837 18284 1946 18325
rect 2048 18284 2056 18325
rect 1837 18250 1943 18284
rect 2049 18250 2056 18284
rect 1837 18209 1946 18250
rect 2048 18209 2056 18250
rect 1837 18175 1943 18209
rect 2049 18175 2056 18209
rect 1837 18134 1946 18175
rect 2048 18134 2056 18175
rect 1837 18100 1943 18134
rect 2049 18100 2056 18134
rect 1837 18059 1946 18100
rect 2048 18059 2056 18100
rect 1837 18025 1943 18059
rect 2049 18025 2056 18059
rect 1837 17984 1946 18025
rect 2048 17984 2056 18025
rect 1837 17950 1943 17984
rect 2049 17950 2056 17984
rect 1837 17909 1946 17950
rect 2048 17909 2056 17950
rect 1837 17875 1943 17909
rect 2049 17875 2056 17909
rect 1837 16100 1946 17875
rect 2048 16630 2056 17875
rect 4314 19985 4382 20019
rect 4416 19985 4450 20019
rect 4484 19985 4518 20019
rect 4552 19985 4586 20019
rect 4620 19985 4654 20019
rect 4688 19985 4722 20019
rect 4756 19985 4790 20019
rect 4824 19985 4858 20019
rect 4892 19985 4926 20019
rect 4960 19985 4994 20019
rect 5028 19985 5062 20019
rect 5096 19985 5130 20019
rect 5164 19985 5198 20019
rect 5232 19985 5266 20019
rect 5300 19985 5334 20019
rect 5368 19985 5402 20019
rect 5436 19985 5470 20019
rect 5504 19985 5538 20019
rect 5572 19985 5606 20019
rect 5640 19985 5674 20019
rect 5708 19985 5742 20019
rect 5776 19985 5810 20019
rect 5844 19985 5878 20019
rect 5912 19985 5946 20019
rect 5980 19985 6014 20019
rect 6048 19985 6082 20019
rect 6116 19985 6150 20019
rect 6184 19985 6218 20019
rect 6252 19985 6286 20019
rect 6320 19985 6354 20019
rect 6388 19985 6422 20019
rect 6456 19985 6490 20019
rect 6524 19985 6558 20019
rect 6592 19985 6626 20019
rect 6660 19985 6694 20019
rect 6728 19985 6762 20019
rect 6796 19985 6830 20019
rect 6864 19985 6898 20019
rect 6932 19985 6966 20019
rect 7000 19985 7034 20019
rect 7068 19985 7102 20019
rect 7136 19985 7170 20019
rect 7204 19985 7238 20019
rect 7272 19985 7306 20019
rect 7340 19985 7374 20019
rect 7408 19985 7442 20019
rect 7476 19985 7510 20019
rect 7544 19985 7578 20019
rect 7612 19985 7646 20019
rect 7680 19985 7714 20019
rect 7748 19985 7782 20019
rect 7816 19985 7850 20019
rect 7884 19985 7918 20019
rect 7952 19985 7986 20019
rect 8020 19985 8054 20019
rect 8088 19985 8122 20019
rect 8156 19985 8190 20019
rect 8224 19985 8258 20019
rect 8292 19985 8326 20019
rect 8360 19985 8394 20019
rect 8428 19985 8462 20019
rect 8496 19985 8530 20019
rect 8564 19985 8598 20019
rect 8632 19985 8666 20019
rect 8700 19985 8734 20019
rect 8768 19985 8802 20019
rect 8836 19985 8870 20019
rect 8904 19985 8938 20019
rect 8972 19985 9006 20019
rect 9040 19985 9074 20019
rect 9108 19985 9142 20019
rect 9176 19985 9210 20019
rect 9244 19985 9278 20019
rect 9312 19985 9346 20019
rect 9380 19985 9414 20019
rect 9448 19985 9482 20019
rect 9516 19985 9550 20019
rect 9584 19985 9618 20019
rect 9652 19985 9686 20019
rect 9720 19985 9754 20019
rect 9788 19985 9822 20019
rect 9856 19985 9890 20019
rect 9924 19985 9958 20019
rect 9992 19985 10026 20019
rect 10060 19985 10094 20019
rect 10128 19985 10162 20019
rect 10196 19985 10230 20019
rect 10264 19985 10298 20019
rect 10332 19985 10366 20019
rect 10400 19985 10434 20019
rect 10468 19985 10502 20019
rect 10536 19985 10570 20019
rect 10604 19985 10638 20019
rect 10672 19985 10706 20019
rect 10740 19985 10774 20019
rect 10808 19985 10842 20019
rect 10876 19985 10910 20019
rect 10944 19985 10978 20019
rect 11012 19985 11046 20019
rect 11080 19985 11114 20019
rect 11148 19985 11182 20019
rect 11216 19985 11250 20019
rect 11284 19985 11318 20019
rect 11352 19985 11386 20019
rect 11420 19985 11454 20019
rect 11488 19985 11522 20019
rect 11556 19985 11590 20019
rect 11624 19985 11658 20019
rect 11692 19985 11726 20019
rect 11760 19985 11794 20019
rect 11828 19985 11862 20019
rect 11896 19985 11930 20019
rect 11964 19985 11998 20019
rect 12032 19985 12066 20019
rect 12100 19985 12134 20019
rect 12168 19985 12202 20019
rect 12236 19985 12270 20019
rect 12304 19985 12338 20019
rect 12372 19985 12406 20019
rect 12440 19985 12474 20019
rect 12508 19985 12542 20019
rect 12576 19985 12610 20019
rect 12644 19985 12678 20019
rect 12712 19985 12746 20019
rect 12780 19985 12814 20019
rect 12848 19985 12882 20019
rect 12916 19985 12950 20019
rect 12984 19985 13018 20019
rect 13052 19985 13086 20019
rect 13120 19985 13154 20019
rect 13188 19985 13222 20019
rect 13256 19985 13290 20019
rect 13324 19985 13358 20019
rect 13392 19985 13426 20019
rect 13460 19985 13494 20019
rect 13528 19985 13562 20019
rect 13596 19985 13630 20019
rect 13664 19985 13838 20019
rect 4314 19894 4348 19985
rect 4314 19826 4348 19860
rect 4314 19758 4348 19792
rect 4314 19690 4348 19724
rect 4314 19622 4348 19656
rect 4314 19554 4348 19588
rect 4554 19798 4578 19832
rect 4612 19798 4647 19832
rect 4681 19798 4716 19832
rect 4750 19798 4785 19832
rect 4819 19798 4854 19832
rect 4888 19798 4923 19832
rect 4957 19798 4992 19832
rect 5026 19798 5061 19832
rect 5095 19798 5130 19832
rect 5164 19798 5199 19832
rect 5233 19798 5268 19832
rect 5302 19798 5337 19832
rect 5371 19798 5406 19832
rect 5440 19798 5475 19832
rect 5509 19798 5544 19832
rect 5578 19798 5613 19832
rect 5647 19798 5682 19832
rect 5716 19798 5750 19832
rect 5784 19798 5818 19832
rect 5852 19798 5886 19832
rect 5920 19798 5954 19832
rect 5988 19798 6022 19832
rect 6056 19798 6090 19832
rect 6124 19798 6158 19832
rect 6192 19798 6226 19832
rect 6260 19798 6294 19832
rect 6328 19798 6362 19832
rect 6396 19798 6430 19832
rect 6464 19798 6498 19832
rect 6532 19798 6566 19832
rect 6600 19798 6634 19832
rect 6668 19798 6702 19832
rect 6736 19798 6770 19832
rect 6804 19798 6838 19832
rect 6872 19798 6906 19832
rect 6940 19798 6974 19832
rect 7008 19798 7042 19832
rect 7076 19798 7110 19832
rect 7144 19798 7178 19832
rect 7212 19798 7246 19832
rect 7280 19798 7314 19832
rect 7348 19798 7382 19832
rect 7416 19798 7450 19832
rect 7484 19798 7518 19832
rect 7552 19798 7586 19832
rect 7620 19798 7654 19832
rect 7688 19798 7722 19832
rect 7756 19798 7790 19832
rect 7824 19798 7858 19832
rect 7892 19798 7926 19832
rect 7960 19798 7994 19832
rect 8028 19798 8062 19832
rect 8096 19798 8130 19832
rect 8164 19798 8198 19832
rect 8232 19798 8266 19832
rect 8300 19798 8334 19832
rect 8368 19798 8402 19832
rect 8436 19798 8470 19832
rect 8504 19798 8538 19832
rect 8572 19798 8606 19832
rect 8640 19798 8674 19832
rect 8708 19798 8742 19832
rect 8776 19798 8810 19832
rect 8844 19798 8878 19832
rect 8912 19798 8946 19832
rect 8980 19798 9014 19832
rect 9048 19798 9082 19832
rect 9116 19798 9150 19832
rect 9184 19798 9218 19832
rect 9252 19798 9286 19832
rect 9320 19798 9354 19832
rect 9388 19798 9422 19832
rect 9456 19798 9490 19832
rect 9524 19798 9558 19832
rect 9592 19798 9626 19832
rect 9660 19798 9694 19832
rect 9728 19798 9762 19832
rect 9796 19798 9830 19832
rect 9864 19798 9898 19832
rect 9932 19798 9966 19832
rect 10000 19798 10034 19832
rect 10068 19798 10102 19832
rect 10136 19798 10170 19832
rect 10204 19798 10238 19832
rect 10272 19798 10306 19832
rect 10340 19798 10374 19832
rect 10408 19798 10442 19832
rect 10476 19798 10510 19832
rect 10544 19798 10578 19832
rect 10612 19798 10646 19832
rect 10680 19798 10714 19832
rect 10748 19798 10782 19832
rect 10816 19798 10850 19832
rect 10884 19798 10918 19832
rect 10952 19798 10986 19832
rect 11020 19798 11054 19832
rect 11088 19798 11122 19832
rect 11156 19798 11190 19832
rect 11224 19798 11258 19832
rect 11292 19798 11326 19832
rect 11360 19798 11394 19832
rect 11428 19798 11462 19832
rect 11496 19798 11530 19832
rect 11564 19798 11598 19832
rect 11632 19798 11666 19832
rect 11700 19798 11734 19832
rect 11768 19798 11802 19832
rect 11836 19798 11870 19832
rect 11904 19798 11938 19832
rect 11972 19798 12006 19832
rect 12040 19798 12074 19832
rect 12108 19798 12142 19832
rect 12176 19798 12210 19832
rect 12244 19798 12278 19832
rect 12312 19798 12346 19832
rect 12380 19798 12414 19832
rect 12448 19798 12482 19832
rect 12516 19798 12550 19832
rect 12584 19798 12618 19832
rect 12652 19798 12686 19832
rect 12720 19798 12754 19832
rect 12788 19798 12822 19832
rect 12856 19798 12890 19832
rect 12924 19798 12958 19832
rect 12992 19798 13026 19832
rect 13060 19798 13094 19832
rect 13128 19798 13162 19832
rect 13196 19798 13230 19832
rect 13264 19798 13298 19832
rect 13332 19798 13366 19832
rect 13400 19798 13434 19832
rect 13468 19798 13502 19832
rect 13536 19798 13570 19832
rect 13604 19798 13628 19832
rect 4554 19764 4656 19798
rect 13458 19745 13628 19798
rect 4977 19708 4996 19742
rect 5045 19708 5069 19742
rect 5113 19708 5142 19742
rect 5181 19708 5215 19742
rect 5249 19708 5283 19742
rect 5322 19708 5351 19742
rect 5395 19708 5419 19742
rect 5468 19708 5487 19742
rect 5541 19708 5555 19742
rect 5614 19708 5623 19742
rect 5687 19708 5691 19742
rect 5725 19708 5726 19742
rect 5793 19708 5799 19742
rect 5861 19708 5872 19742
rect 5929 19708 5945 19742
rect 5997 19708 6017 19742
rect 6065 19708 6089 19742
rect 6133 19708 6161 19742
rect 6201 19708 6233 19742
rect 6269 19708 6303 19742
rect 6339 19708 6371 19742
rect 6411 19708 6439 19742
rect 6483 19708 6507 19742
rect 6555 19708 6575 19742
rect 6627 19708 6643 19742
rect 6699 19708 6711 19742
rect 6771 19708 6779 19742
rect 6843 19708 6847 19742
rect 6949 19708 6953 19742
rect 7017 19708 7025 19742
rect 7085 19708 7097 19742
rect 7153 19708 7169 19742
rect 7221 19708 7241 19742
rect 7289 19708 7313 19742
rect 7357 19708 7385 19742
rect 7425 19708 7457 19742
rect 7493 19708 7527 19742
rect 7563 19708 7595 19742
rect 7635 19708 7663 19742
rect 7707 19708 7731 19742
rect 7779 19708 7799 19742
rect 7851 19708 7867 19742
rect 7923 19708 7935 19742
rect 7995 19708 8003 19742
rect 8067 19708 8071 19742
rect 8173 19708 8177 19742
rect 8241 19708 8249 19742
rect 8309 19708 8321 19742
rect 8377 19708 8393 19742
rect 8445 19708 8465 19742
rect 8513 19708 8537 19742
rect 8581 19708 8609 19742
rect 8649 19708 8681 19742
rect 8717 19708 8751 19742
rect 8787 19708 8819 19742
rect 8859 19708 8887 19742
rect 8931 19708 8955 19742
rect 9003 19708 9023 19742
rect 9075 19708 9091 19742
rect 9147 19708 9159 19742
rect 9219 19708 9227 19742
rect 9291 19708 9295 19742
rect 9397 19708 9401 19742
rect 9465 19708 9473 19742
rect 9533 19708 9545 19742
rect 9601 19708 9617 19742
rect 9669 19708 9689 19742
rect 9737 19708 9761 19742
rect 9805 19708 9833 19742
rect 9873 19708 9905 19742
rect 9941 19708 9975 19742
rect 10011 19708 10043 19742
rect 10083 19708 10111 19742
rect 10155 19708 10179 19742
rect 10227 19708 10247 19742
rect 10299 19708 10315 19742
rect 10371 19708 10383 19742
rect 10443 19708 10451 19742
rect 10515 19708 10519 19742
rect 10621 19708 10625 19742
rect 10689 19708 10697 19742
rect 10757 19708 10769 19742
rect 10825 19708 10841 19742
rect 10893 19708 10913 19742
rect 10961 19708 10985 19742
rect 11029 19708 11057 19742
rect 11097 19708 11129 19742
rect 11165 19708 11199 19742
rect 11235 19708 11267 19742
rect 11307 19708 11335 19742
rect 11379 19708 11403 19742
rect 11451 19708 11471 19742
rect 11523 19708 11539 19742
rect 11595 19708 11607 19742
rect 11667 19708 11675 19742
rect 11739 19708 11743 19742
rect 11845 19708 11849 19742
rect 11913 19708 11921 19742
rect 11981 19708 11993 19742
rect 12049 19708 12065 19742
rect 12117 19708 12137 19742
rect 12185 19708 12209 19742
rect 12253 19708 12281 19742
rect 12321 19708 12353 19742
rect 12389 19708 12423 19742
rect 12459 19708 12491 19742
rect 12531 19708 12559 19742
rect 12603 19708 12627 19742
rect 12675 19708 12695 19742
rect 12747 19708 12763 19742
rect 12819 19708 12831 19742
rect 12891 19708 12899 19742
rect 12963 19708 12967 19742
rect 13001 19708 13035 19742
rect 13069 19708 13103 19742
rect 13137 19708 13171 19742
rect 13205 19708 13239 19742
rect 13273 19708 13331 19742
rect 13458 19701 13490 19745
rect 13596 19701 13628 19745
rect 4314 19486 4348 19520
rect 4314 19418 4348 19452
rect 4314 19350 4348 19384
rect 4314 19282 4348 19316
rect 4314 19214 4348 19248
rect 4314 19146 4348 19180
rect 4314 19078 4348 19112
rect 4314 19010 4348 19044
rect 4314 18942 4348 18976
rect 4314 18874 4348 18908
rect 4314 18806 4348 18840
rect 4314 18738 4348 18772
rect 4314 18670 4348 18704
rect 4314 18602 4348 18636
rect 4314 18534 4348 18568
rect 4314 18466 4348 18500
rect 4314 18398 4348 18432
rect 4314 18330 4348 18364
rect 4314 18262 4348 18296
rect 4314 18194 4348 18228
rect 4314 18126 4348 18160
rect 4314 18058 4348 18092
rect 4314 17990 4348 18024
rect 4314 17922 4348 17956
rect 4314 17854 4348 17888
rect 4314 17786 4348 17820
rect 4314 17718 4348 17752
rect 4314 17650 4348 17684
rect 4314 17582 4348 17616
rect 4314 17514 4348 17548
rect 4314 17446 4348 17480
rect 4314 17378 4348 17412
rect 4314 17310 4348 17344
rect 4314 17242 4348 17276
rect 4314 17174 4348 17208
rect 4314 17106 4348 17140
rect 4314 17038 4348 17072
rect 4314 16970 4348 17004
rect 2218 16883 2258 16917
rect 2292 16883 2332 16917
rect 2184 16798 2366 16883
rect 2218 16764 2258 16798
rect 2292 16764 2332 16798
rect 3933 16883 3973 16917
rect 4007 16883 4047 16917
rect 3899 16798 4081 16883
rect 3933 16764 3973 16798
rect 4007 16764 4047 16798
rect 4314 16902 4348 16936
rect 4314 16834 4348 16868
rect 4314 16766 4348 16800
rect 4314 16698 4348 16732
rect 4314 16630 4348 16664
rect 2048 16596 2208 16630
rect 2242 16596 2276 16630
rect 2310 16596 2344 16630
rect 2378 16596 2412 16630
rect 2446 16596 2480 16630
rect 2514 16596 2548 16630
rect 2582 16596 2616 16630
rect 2650 16596 2684 16630
rect 2718 16596 2752 16630
rect 2786 16596 2820 16630
rect 2854 16596 2888 16630
rect 2922 16596 2956 16630
rect 2990 16596 3024 16630
rect 3058 16596 3092 16630
rect 3126 16596 3160 16630
rect 3194 16596 3228 16630
rect 3262 16596 3296 16630
rect 3330 16596 3364 16630
rect 3398 16596 3432 16630
rect 3466 16596 3500 16630
rect 3534 16596 3568 16630
rect 3602 16596 3636 16630
rect 3670 16596 3704 16630
rect 3738 16596 3772 16630
rect 3806 16596 3840 16630
rect 3874 16596 3908 16630
rect 3942 16596 3976 16630
rect 4010 16596 4044 16630
rect 4078 16596 4112 16630
rect 4146 16596 4180 16630
rect 4214 16596 4348 16630
rect 4520 19544 4554 19578
rect 4486 19505 4554 19544
rect 4520 19471 4554 19505
rect 4486 19432 4554 19471
rect 4520 19398 4554 19432
rect 4486 19359 4554 19398
rect 4520 19325 4554 19359
rect 4486 19286 4554 19325
rect 4520 19252 4554 19286
rect 4486 19213 4554 19252
rect 4520 19179 4554 19213
rect 4486 19140 4554 19179
rect 4520 19106 4554 19140
rect 4486 19067 4554 19106
rect 4520 19033 4554 19067
rect 4486 18994 4554 19033
rect 4520 18960 4554 18994
rect 4486 18921 4554 18960
rect 4520 18887 4554 18921
rect 4486 18848 4554 18887
rect 4520 18814 4554 18848
rect 4486 18775 4554 18814
rect 4520 18741 4554 18775
rect 4486 18702 4554 18741
rect 4520 18668 4554 18702
rect 4486 18629 4554 18668
rect 4520 18595 4554 18629
rect 4486 18556 4554 18595
rect 4520 18522 4554 18556
rect 4486 18483 4554 18522
rect 4520 18449 4554 18483
rect 4486 18410 4554 18449
rect 4520 18376 4554 18410
rect 4486 18337 4554 18376
rect 4520 18303 4554 18337
rect 4486 18264 4554 18303
rect 4520 18230 4554 18264
rect 4771 19580 4809 19614
rect 4737 19540 4843 19580
rect 4771 19506 4809 19540
rect 4737 19466 4843 19506
rect 4771 19432 4809 19466
rect 4737 19392 4843 19432
rect 4771 19358 4809 19392
rect 13342 19498 13376 19540
rect 13342 19422 13376 19464
rect 4737 19318 4843 19358
rect 4771 19284 4809 19318
rect 4737 19244 4843 19284
rect 4771 19210 4809 19244
rect 4737 19170 4843 19210
rect 4771 19136 4809 19170
rect 4737 19096 4843 19136
rect 4771 19062 4809 19096
rect 4737 19022 4843 19062
rect 4771 18988 4809 19022
rect 4737 18948 4843 18988
rect 4771 18914 4809 18948
rect 4737 18874 4843 18914
rect 4771 18840 4809 18874
rect 4737 18801 4843 18840
rect 4771 18767 4809 18801
rect 4737 18728 4843 18767
rect 4771 18694 4809 18728
rect 4737 18655 4843 18694
rect 4771 18621 4809 18655
rect 4737 18582 4843 18621
rect 4771 18548 4809 18582
rect 4737 18509 4843 18548
rect 4771 18475 4809 18509
rect 4737 18436 4843 18475
rect 4771 18402 4809 18436
rect 4737 18363 4843 18402
rect 5062 19310 5096 19351
rect 5062 19235 5096 19276
rect 5062 19160 5096 19201
rect 5062 19086 5096 19126
rect 5062 19012 5096 19052
rect 5062 18938 5096 18978
rect 5062 18864 5096 18904
rect 5062 18790 5096 18830
rect 5062 18716 5096 18756
rect 5062 18642 5096 18682
rect 5062 18568 5096 18608
rect 5062 18494 5096 18534
rect 5062 18420 5096 18460
rect 6718 19310 6752 19351
rect 6718 19235 6752 19276
rect 6718 19160 6752 19201
rect 6718 19086 6752 19126
rect 6718 19012 6752 19052
rect 6718 18938 6752 18978
rect 6718 18864 6752 18904
rect 6718 18790 6752 18830
rect 6718 18716 6752 18756
rect 6718 18642 6752 18682
rect 6718 18568 6752 18608
rect 6718 18494 6752 18534
rect 6718 18420 6752 18460
rect 8374 19310 8408 19351
rect 8374 19235 8408 19276
rect 8374 19160 8408 19201
rect 8374 19086 8408 19126
rect 8374 19012 8408 19052
rect 8374 18938 8408 18978
rect 8374 18864 8408 18904
rect 8374 18790 8408 18830
rect 8374 18716 8408 18756
rect 8374 18642 8408 18682
rect 8374 18568 8408 18608
rect 8374 18494 8408 18534
rect 8374 18420 8408 18460
rect 10030 19310 10064 19351
rect 10030 19235 10064 19276
rect 10030 19160 10064 19201
rect 10030 19086 10064 19126
rect 10030 19012 10064 19052
rect 10030 18938 10064 18978
rect 10030 18864 10064 18904
rect 10030 18790 10064 18830
rect 10030 18716 10064 18756
rect 10030 18642 10064 18682
rect 10030 18568 10064 18608
rect 10030 18494 10064 18534
rect 10030 18420 10064 18460
rect 11686 19310 11720 19351
rect 11686 19235 11720 19276
rect 11686 19160 11720 19201
rect 11686 19086 11720 19126
rect 11686 19012 11720 19052
rect 11686 18938 11720 18978
rect 11686 18864 11720 18904
rect 11686 18790 11720 18830
rect 11686 18716 11720 18756
rect 11686 18642 11720 18682
rect 11686 18568 11720 18608
rect 11686 18494 11720 18534
rect 11686 18420 11720 18460
rect 13342 19346 13376 19388
rect 13342 19270 13376 19312
rect 13342 19194 13376 19236
rect 13342 19118 13376 19160
rect 13342 19042 13376 19084
rect 13342 18966 13376 19008
rect 13342 18890 13376 18932
rect 13342 18815 13376 18856
rect 13342 18740 13376 18781
rect 13342 18665 13376 18706
rect 13342 18590 13376 18631
rect 13342 18515 13376 18556
rect 13342 18440 13376 18481
rect 4771 18329 4809 18363
rect 4737 18290 4843 18329
rect 4771 18256 4809 18290
rect 13342 18365 13376 18406
rect 13342 18290 13376 18331
rect 4486 18191 4554 18230
rect 4520 18157 4554 18191
rect 4486 18118 4554 18157
rect 4656 18135 4754 18169
rect 4788 18135 4822 18169
rect 4856 18135 4890 18169
rect 4924 18135 4958 18169
rect 4992 18135 5026 18169
rect 5060 18135 5094 18169
rect 5128 18135 5162 18169
rect 5196 18135 5230 18169
rect 5264 18135 5298 18169
rect 5332 18135 5366 18169
rect 5400 18135 5434 18169
rect 5468 18135 5502 18169
rect 5536 18135 5570 18169
rect 5604 18135 5638 18169
rect 5672 18135 5706 18169
rect 5740 18135 5774 18169
rect 5808 18135 5842 18169
rect 5876 18135 5910 18169
rect 5944 18135 5978 18169
rect 6012 18135 6046 18169
rect 6080 18135 6114 18169
rect 6148 18135 6182 18169
rect 6216 18135 6250 18169
rect 6284 18135 6318 18169
rect 6352 18135 6386 18169
rect 6420 18135 6454 18169
rect 6488 18135 6522 18169
rect 6556 18135 6590 18169
rect 6624 18135 6658 18169
rect 6692 18135 6726 18169
rect 6760 18135 6794 18169
rect 6828 18135 6862 18169
rect 6896 18135 6930 18169
rect 6964 18135 6998 18169
rect 7032 18135 7066 18169
rect 7100 18135 7134 18169
rect 7168 18135 7202 18169
rect 7236 18135 7270 18169
rect 7304 18135 7338 18169
rect 7372 18135 7406 18169
rect 7440 18135 7474 18169
rect 7508 18135 7542 18169
rect 7576 18135 7610 18169
rect 7644 18135 7678 18169
rect 7712 18135 7746 18169
rect 7780 18135 7814 18169
rect 7848 18135 7882 18169
rect 7916 18135 7950 18169
rect 7984 18135 8018 18169
rect 8052 18135 8086 18169
rect 8120 18135 8154 18169
rect 8188 18135 8222 18169
rect 8256 18135 8290 18169
rect 8324 18135 8358 18169
rect 8392 18135 8426 18169
rect 8460 18135 8494 18169
rect 8528 18135 8562 18169
rect 8596 18135 8630 18169
rect 8664 18135 8698 18169
rect 8732 18135 8766 18169
rect 8800 18135 8834 18169
rect 8868 18135 8902 18169
rect 8936 18135 8970 18169
rect 9004 18135 9038 18169
rect 9072 18135 9106 18169
rect 9140 18135 9174 18169
rect 9208 18135 9242 18169
rect 9276 18135 9310 18169
rect 9344 18135 9378 18169
rect 9412 18135 9446 18169
rect 9480 18135 9514 18169
rect 9548 18135 9582 18169
rect 9616 18135 9650 18169
rect 9684 18135 9718 18169
rect 9752 18135 9786 18169
rect 9820 18135 9854 18169
rect 9888 18135 9922 18169
rect 9956 18135 9990 18169
rect 10024 18135 10058 18169
rect 10092 18135 10126 18169
rect 10160 18135 10194 18169
rect 10228 18135 10262 18169
rect 10296 18135 10330 18169
rect 10364 18135 10398 18169
rect 10432 18135 10466 18169
rect 10500 18135 10534 18169
rect 10568 18135 10602 18169
rect 10636 18135 10670 18169
rect 10704 18135 10738 18169
rect 10772 18135 10806 18169
rect 10840 18135 10874 18169
rect 10908 18135 10942 18169
rect 10976 18135 11010 18169
rect 11044 18135 11078 18169
rect 11112 18135 11146 18169
rect 11180 18135 11214 18169
rect 11248 18135 11282 18169
rect 11316 18135 11350 18169
rect 11384 18135 11418 18169
rect 11452 18135 11486 18169
rect 11520 18135 11554 18169
rect 11588 18135 11622 18169
rect 11656 18135 11690 18169
rect 11724 18135 11758 18169
rect 11792 18135 11826 18169
rect 11860 18135 11894 18169
rect 11928 18135 11962 18169
rect 11996 18135 12030 18169
rect 12064 18135 12098 18169
rect 12132 18135 12166 18169
rect 12200 18135 12234 18169
rect 12268 18135 12302 18169
rect 12336 18135 12370 18169
rect 12404 18135 12438 18169
rect 12472 18135 12506 18169
rect 12540 18135 12574 18169
rect 12608 18135 12642 18169
rect 12676 18135 12710 18169
rect 12744 18135 12778 18169
rect 12812 18135 12846 18169
rect 12880 18135 12914 18169
rect 12948 18135 12982 18169
rect 13016 18135 13050 18169
rect 13084 18135 13118 18169
rect 13152 18135 13186 18169
rect 13220 18135 13254 18169
rect 13288 18135 13322 18169
rect 13356 18135 13390 18169
rect 13424 18135 13458 18169
rect 4520 18084 4554 18118
rect 4486 18045 4554 18084
rect 4520 18011 4554 18045
rect 4486 17972 4554 18011
rect 4977 18009 4996 18043
rect 5045 18009 5069 18043
rect 5113 18009 5142 18043
rect 5181 18009 5215 18043
rect 5249 18009 5283 18043
rect 5322 18009 5351 18043
rect 5395 18009 5419 18043
rect 5468 18009 5487 18043
rect 5541 18009 5555 18043
rect 5614 18009 5623 18043
rect 5687 18009 5691 18043
rect 5725 18009 5726 18043
rect 5793 18009 5799 18043
rect 5861 18009 5872 18043
rect 5929 18009 5945 18043
rect 5997 18009 6017 18043
rect 6065 18009 6089 18043
rect 6133 18009 6161 18043
rect 6201 18009 6233 18043
rect 6269 18009 6303 18043
rect 6339 18009 6371 18043
rect 6411 18009 6439 18043
rect 6483 18009 6507 18043
rect 6555 18009 6575 18043
rect 6627 18009 6643 18043
rect 6699 18009 6711 18043
rect 6771 18009 6779 18043
rect 6843 18009 6847 18043
rect 6949 18009 6953 18043
rect 7017 18009 7025 18043
rect 7085 18009 7097 18043
rect 7153 18009 7169 18043
rect 7221 18009 7241 18043
rect 7289 18009 7313 18043
rect 7357 18009 7385 18043
rect 7425 18009 7457 18043
rect 7493 18009 7527 18043
rect 7563 18009 7595 18043
rect 7635 18009 7663 18043
rect 7707 18009 7731 18043
rect 7779 18009 7799 18043
rect 7851 18009 7867 18043
rect 7923 18009 7935 18043
rect 7995 18009 8003 18043
rect 8067 18009 8071 18043
rect 8173 18009 8177 18043
rect 8241 18009 8249 18043
rect 8309 18009 8321 18043
rect 8377 18009 8393 18043
rect 8445 18009 8465 18043
rect 8513 18009 8537 18043
rect 8581 18009 8609 18043
rect 8649 18009 8681 18043
rect 8717 18009 8751 18043
rect 8787 18009 8819 18043
rect 8859 18009 8887 18043
rect 8931 18009 8955 18043
rect 9003 18009 9023 18043
rect 9075 18009 9091 18043
rect 9147 18009 9159 18043
rect 9219 18009 9227 18043
rect 9291 18009 9295 18043
rect 9397 18009 9401 18043
rect 9465 18009 9473 18043
rect 9533 18009 9545 18043
rect 9601 18009 9617 18043
rect 9669 18009 9689 18043
rect 9737 18009 9761 18043
rect 9805 18009 9833 18043
rect 9873 18009 9905 18043
rect 9941 18009 9975 18043
rect 10011 18009 10043 18043
rect 10083 18009 10111 18043
rect 10155 18009 10179 18043
rect 10227 18009 10247 18043
rect 10299 18009 10315 18043
rect 10371 18009 10383 18043
rect 10443 18009 10451 18043
rect 10515 18009 10519 18043
rect 10621 18009 10625 18043
rect 10689 18009 10697 18043
rect 10757 18009 10769 18043
rect 10825 18009 10841 18043
rect 10893 18009 10913 18043
rect 10961 18009 10985 18043
rect 11029 18009 11057 18043
rect 11097 18009 11129 18043
rect 11165 18009 11199 18043
rect 11235 18009 11267 18043
rect 11307 18009 11335 18043
rect 11379 18009 11403 18043
rect 11451 18009 11471 18043
rect 11523 18009 11539 18043
rect 11595 18009 11607 18043
rect 11667 18009 11675 18043
rect 11739 18009 11743 18043
rect 11845 18009 11849 18043
rect 11913 18009 11921 18043
rect 11981 18009 11993 18043
rect 12049 18009 12065 18043
rect 12117 18009 12137 18043
rect 12185 18009 12209 18043
rect 12253 18009 12281 18043
rect 12321 18009 12353 18043
rect 12389 18009 12423 18043
rect 12459 18009 12491 18043
rect 12531 18009 12559 18043
rect 12603 18009 12627 18043
rect 12675 18009 12695 18043
rect 12747 18009 12763 18043
rect 12819 18009 12831 18043
rect 12891 18009 12899 18043
rect 12963 18009 12967 18043
rect 13001 18009 13035 18043
rect 13069 18009 13103 18043
rect 13137 18009 13171 18043
rect 13205 18009 13239 18043
rect 13273 18009 13331 18043
rect 4520 17938 4554 17972
rect 4486 17899 4554 17938
rect 4520 17865 4554 17899
rect 4486 17826 4554 17865
rect 4520 17792 4554 17826
rect 4486 17753 4554 17792
rect 4520 17719 4554 17753
rect 4486 17679 4554 17719
rect 4520 17645 4554 17679
rect 4486 17605 4554 17645
rect 4520 17571 4554 17605
rect 4486 17531 4554 17571
rect 4520 17497 4554 17531
rect 4486 17457 4554 17497
rect 4520 17423 4554 17457
rect 4486 17383 4554 17423
rect 4520 17349 4554 17383
rect 4486 17309 4554 17349
rect 4520 17275 4554 17309
rect 4486 17235 4554 17275
rect 4520 17201 4554 17235
rect 4486 17161 4554 17201
rect 4520 17127 4554 17161
rect 4486 17087 4554 17127
rect 4520 17053 4554 17087
rect 4486 17013 4554 17053
rect 4520 16979 4554 17013
rect 4486 16939 4554 16979
rect 4520 16905 4554 16939
rect 4486 16865 4554 16905
rect 4520 16831 4554 16865
rect 4486 16791 4554 16831
rect 4520 16757 4554 16791
rect 4486 16717 4554 16757
rect 4520 16683 4554 16717
rect 4486 16643 4554 16683
rect 4520 16609 4554 16643
rect 2048 16100 2056 16596
rect 4486 16569 4554 16609
rect 4520 16535 4554 16569
rect 4771 17881 4809 17915
rect 4737 17841 4843 17881
rect 4771 17807 4809 17841
rect 4737 17767 4843 17807
rect 4771 17733 4809 17767
rect 4737 17693 4843 17733
rect 4771 17659 4809 17693
rect 4737 17619 4843 17659
rect 4771 17585 4809 17619
rect 4737 17545 4843 17585
rect 4771 17511 4809 17545
rect 4737 17471 4843 17511
rect 4771 17437 4809 17471
rect 4737 17397 4843 17437
rect 4771 17363 4809 17397
rect 4737 17323 4843 17363
rect 4771 17289 4809 17323
rect 4737 17249 4843 17289
rect 4771 17215 4809 17249
rect 4737 17175 4843 17215
rect 4771 17141 4809 17175
rect 4737 17102 4843 17141
rect 4771 17068 4809 17102
rect 4737 17029 4843 17068
rect 4771 16995 4809 17029
rect 4737 16956 4843 16995
rect 4771 16922 4809 16956
rect 4737 16883 4843 16922
rect 4771 16849 4809 16883
rect 4737 16810 4843 16849
rect 4771 16776 4809 16810
rect 4737 16737 4843 16776
rect 4771 16703 4809 16737
rect 4737 16664 4843 16703
rect 4771 16630 4809 16664
rect 4737 16591 4843 16630
rect 4771 16557 4809 16591
rect 5062 17730 5096 17770
rect 5062 17656 5096 17696
rect 5062 17582 5096 17622
rect 5062 17508 5096 17548
rect 5062 17434 5096 17474
rect 5062 17360 5096 17400
rect 5062 17286 5096 17326
rect 5062 17212 5096 17252
rect 5062 17138 5096 17178
rect 5062 17064 5096 17104
rect 5062 16990 5096 17030
rect 5062 16916 5096 16956
rect 5062 16842 5096 16882
rect 5062 16767 5096 16808
rect 5062 16692 5096 16733
rect 5062 16617 5096 16658
rect 6718 17730 6752 17770
rect 6718 17656 6752 17696
rect 6718 17582 6752 17622
rect 6718 17508 6752 17548
rect 6718 17434 6752 17474
rect 6718 17360 6752 17400
rect 6718 17286 6752 17326
rect 6718 17212 6752 17252
rect 6718 17138 6752 17178
rect 6718 17064 6752 17104
rect 6718 16990 6752 17030
rect 6718 16916 6752 16956
rect 6718 16842 6752 16882
rect 6718 16767 6752 16808
rect 6718 16692 6752 16733
rect 6718 16617 6752 16658
rect 8374 17730 8408 17770
rect 8374 17656 8408 17696
rect 8374 17582 8408 17622
rect 8374 17508 8408 17548
rect 8374 17434 8408 17474
rect 8374 17360 8408 17400
rect 8374 17286 8408 17326
rect 8374 17212 8408 17252
rect 8374 17138 8408 17178
rect 8374 17064 8408 17104
rect 8374 16990 8408 17030
rect 8374 16916 8408 16956
rect 8374 16842 8408 16882
rect 8374 16767 8408 16808
rect 8374 16692 8408 16733
rect 8374 16617 8408 16658
rect 10030 17730 10064 17770
rect 10030 17656 10064 17696
rect 10030 17582 10064 17622
rect 10030 17508 10064 17548
rect 10030 17434 10064 17474
rect 10030 17360 10064 17400
rect 10030 17286 10064 17326
rect 10030 17212 10064 17252
rect 10030 17138 10064 17178
rect 10030 17064 10064 17104
rect 10030 16990 10064 17030
rect 10030 16916 10064 16956
rect 10030 16842 10064 16882
rect 10030 16767 10064 16808
rect 10030 16692 10064 16733
rect 10030 16617 10064 16658
rect 11686 17730 11720 17770
rect 11686 17656 11720 17696
rect 11686 17582 11720 17622
rect 11686 17508 11720 17548
rect 11686 17434 11720 17474
rect 11686 17360 11720 17400
rect 11686 17286 11720 17326
rect 11686 17212 11720 17252
rect 11686 17138 11720 17178
rect 11686 17064 11720 17104
rect 11686 16990 11720 17030
rect 11686 16916 11720 16956
rect 11686 16842 11720 16882
rect 11686 16767 11720 16808
rect 11686 16692 11720 16733
rect 11686 16617 11720 16658
rect 13342 17800 13376 17841
rect 13342 17725 13376 17766
rect 13342 17650 13376 17691
rect 13342 17575 13376 17616
rect 13342 17500 13376 17541
rect 13342 17425 13376 17466
rect 13342 17350 13376 17391
rect 13342 17275 13376 17316
rect 13342 17199 13376 17241
rect 13342 17123 13376 17165
rect 13342 17047 13376 17089
rect 13342 16971 13376 17013
rect 13342 16895 13376 16937
rect 13342 16819 13376 16861
rect 13342 16743 13376 16785
rect 13342 16667 13376 16709
rect 13342 16591 13376 16633
rect 4486 16495 4554 16535
rect 4520 16466 4554 16495
rect 4520 16461 4622 16466
rect 4656 16461 4754 16470
rect 4486 16436 4754 16461
rect 4788 16436 4822 16470
rect 4856 16436 4890 16470
rect 4924 16436 4958 16470
rect 4992 16436 5026 16470
rect 5060 16436 5094 16470
rect 5128 16436 5162 16470
rect 5196 16436 5230 16470
rect 5264 16436 5298 16470
rect 5332 16436 5366 16470
rect 5400 16436 5434 16470
rect 5468 16436 5502 16470
rect 5536 16436 5570 16470
rect 5604 16436 5638 16470
rect 5672 16436 5706 16470
rect 5740 16436 5774 16470
rect 5808 16436 5842 16470
rect 5876 16436 5910 16470
rect 5944 16436 5978 16470
rect 6012 16436 6046 16470
rect 6080 16436 6114 16470
rect 6148 16436 6182 16470
rect 6216 16436 6250 16470
rect 6284 16436 6318 16470
rect 6352 16436 6386 16470
rect 6420 16436 6454 16470
rect 6488 16436 6522 16470
rect 6556 16436 6590 16470
rect 6624 16436 6658 16470
rect 6692 16436 6726 16470
rect 6760 16436 6794 16470
rect 6828 16436 6862 16470
rect 6896 16436 6930 16470
rect 6964 16436 6998 16470
rect 7032 16436 7066 16470
rect 7100 16436 7134 16470
rect 7168 16436 7202 16470
rect 7236 16436 7270 16470
rect 7304 16436 7338 16470
rect 7372 16436 7406 16470
rect 7440 16436 7474 16470
rect 7508 16436 7542 16470
rect 7576 16436 7610 16470
rect 7644 16436 7678 16470
rect 7712 16436 7746 16470
rect 7780 16436 7814 16470
rect 7848 16436 7882 16470
rect 7916 16436 7950 16470
rect 7984 16436 8018 16470
rect 8052 16436 8086 16470
rect 8120 16436 8154 16470
rect 8188 16436 8222 16470
rect 8256 16436 8290 16470
rect 8324 16436 8358 16470
rect 8392 16436 8426 16470
rect 8460 16436 8494 16470
rect 8528 16436 8562 16470
rect 8596 16436 8630 16470
rect 8664 16436 8698 16470
rect 8732 16436 8766 16470
rect 8800 16436 8834 16470
rect 8868 16436 8902 16470
rect 8936 16436 8970 16470
rect 9004 16436 9038 16470
rect 9072 16436 9106 16470
rect 9140 16436 9174 16470
rect 9208 16436 9242 16470
rect 9276 16436 9310 16470
rect 9344 16436 9378 16470
rect 9412 16436 9446 16470
rect 9480 16436 9514 16470
rect 9548 16436 9582 16470
rect 9616 16436 9650 16470
rect 9684 16436 9718 16470
rect 9752 16436 9786 16470
rect 9820 16436 9854 16470
rect 9888 16436 9922 16470
rect 9956 16436 9990 16470
rect 10024 16436 10058 16470
rect 10092 16436 10126 16470
rect 10160 16436 10194 16470
rect 10228 16436 10262 16470
rect 10296 16436 10330 16470
rect 10364 16436 10398 16470
rect 10432 16436 10466 16470
rect 10500 16436 10534 16470
rect 10568 16436 10602 16470
rect 10636 16436 10670 16470
rect 10704 16436 10738 16470
rect 10772 16436 10806 16470
rect 10840 16436 10874 16470
rect 10908 16436 10942 16470
rect 10976 16436 11010 16470
rect 11044 16436 11078 16470
rect 11112 16436 11146 16470
rect 11180 16436 11214 16470
rect 11248 16436 11282 16470
rect 11316 16436 11350 16470
rect 11384 16436 11418 16470
rect 11452 16436 11486 16470
rect 11520 16436 11554 16470
rect 11588 16436 11622 16470
rect 11656 16436 11690 16470
rect 11724 16436 11758 16470
rect 11792 16436 11826 16470
rect 11860 16436 11894 16470
rect 11928 16436 11962 16470
rect 11996 16436 12030 16470
rect 12064 16436 12098 16470
rect 12132 16436 12166 16470
rect 12200 16436 12234 16470
rect 12268 16436 12302 16470
rect 12336 16436 12370 16470
rect 12404 16436 12438 16470
rect 12472 16436 12506 16470
rect 12540 16436 12574 16470
rect 12608 16436 12642 16470
rect 12676 16436 12710 16470
rect 12744 16436 12778 16470
rect 12812 16436 12846 16470
rect 12880 16436 12914 16470
rect 12948 16436 12982 16470
rect 13016 16436 13050 16470
rect 13084 16436 13118 16470
rect 13152 16436 13186 16470
rect 13220 16436 13254 16470
rect 13288 16436 13322 16470
rect 13356 16436 13390 16470
rect 13424 16436 13458 16470
rect 4486 16432 4656 16436
rect 4486 16421 4622 16432
rect 4520 16417 4622 16421
rect 1837 15922 1944 16100
rect 2050 15922 2056 16100
rect 1837 15883 1946 15922
rect 2048 15883 2056 15922
rect 1837 15849 1944 15883
rect 2050 15849 2056 15883
rect 1837 15810 1946 15849
rect 2048 15810 2056 15849
rect 1837 15776 1944 15810
rect 2050 15776 2056 15810
rect 1837 15737 1946 15776
rect 2048 15737 2056 15776
rect 1837 15703 1944 15737
rect 2050 15703 2056 15737
rect 1837 15664 1946 15703
rect 2048 15664 2056 15703
rect 1837 15630 1944 15664
rect 2050 15630 2056 15664
rect 1837 15591 1946 15630
rect 2048 15591 2056 15630
rect 1837 15557 1944 15591
rect 2050 15557 2056 15591
rect 1837 15518 1946 15557
rect 2048 15518 2056 15557
rect 1837 15484 1944 15518
rect 2050 15484 2056 15518
rect 1837 15445 1946 15484
rect 2048 15445 2056 15484
rect 1837 15411 1944 15445
rect 2050 15411 2056 15445
rect 1837 15372 1946 15411
rect 2048 15372 2056 15411
rect 1837 15338 1944 15372
rect 2050 15338 2056 15372
rect 1837 14974 1946 15338
rect 2048 14974 2056 15338
rect 1837 14940 1944 14974
rect 2050 14940 2056 14974
rect 1837 14899 1946 14940
rect 2048 14899 2056 14940
rect 1837 14865 1944 14899
rect 2050 14865 2056 14899
rect 1837 14824 1946 14865
rect 2048 14824 2056 14865
rect 1837 14790 1944 14824
rect 2050 14790 2056 14824
rect 1837 14749 1946 14790
rect 2048 14749 2056 14790
rect 1837 14715 1944 14749
rect 2050 14715 2056 14749
rect 1837 14674 1946 14715
rect 2048 14674 2056 14715
rect 1837 14640 1944 14674
rect 2050 14640 2056 14674
rect 1837 14599 1946 14640
rect 2048 14599 2056 14640
rect 1837 14565 1944 14599
rect 2050 14565 2056 14599
rect 1837 14524 1946 14565
rect 2048 14524 2056 14565
rect 1837 14490 1944 14524
rect 2050 14490 2056 14524
rect 1837 14449 1946 14490
rect 2048 14449 2056 14490
rect 1837 14415 1944 14449
rect 2050 14415 2056 14449
rect 1837 14374 1946 14415
rect 2048 14374 2056 14415
rect 1837 14340 1944 14374
rect 2050 14340 2056 14374
rect 1837 14299 1946 14340
rect 2048 14299 2056 14340
rect 1837 14265 1944 14299
rect 2050 14265 2056 14299
rect 1837 14224 1946 14265
rect 2048 14224 2056 14265
rect 1837 14190 1944 14224
rect 2050 14190 2056 14224
rect 1837 14149 1946 14190
rect 2048 14149 2056 14190
rect 1837 14115 1944 14149
rect 2050 14115 2056 14149
rect 1837 14075 1946 14115
rect 2048 14075 2056 14115
rect 1837 14041 1944 14075
rect 2050 14041 2056 14075
rect 1837 14001 1946 14041
rect 2048 14001 2056 14041
rect 1837 13967 1944 14001
rect 2050 13967 2056 14001
rect 1837 13927 1946 13967
rect 2048 13927 2056 13967
rect 1837 13893 1944 13927
rect 2050 13893 2056 13927
rect 1837 13853 1946 13893
rect 2048 13853 2056 13893
rect 1837 13819 1944 13853
rect 2050 13819 2056 13853
rect 1837 13779 1946 13819
rect 2048 13779 2056 13819
rect 1837 13745 1944 13779
rect 2050 13745 2056 13779
rect 1837 13705 1946 13745
rect 2048 13705 2056 13745
rect 1837 13671 1944 13705
rect 2050 13671 2056 13705
rect 1837 13631 1946 13671
rect 2048 13631 2056 13671
rect 1837 13597 1944 13631
rect 2050 13597 2056 13631
rect 1837 13557 1946 13597
rect 2048 13557 2056 13597
rect 1837 13523 1944 13557
rect 2050 13523 2056 13557
rect 1837 13483 1946 13523
rect 2048 13483 2056 13523
rect 1837 13449 1944 13483
rect 2050 13449 2056 13483
rect 1837 13409 1946 13449
rect 2048 13409 2056 13449
rect 1837 13375 1944 13409
rect 2050 13375 2056 13409
rect 1837 13335 1946 13375
rect 2048 13335 2056 13375
rect 1837 13301 1944 13335
rect 2050 13301 2056 13335
rect 1837 12889 1946 13301
rect 2048 12889 2056 13301
rect 1837 12855 1944 12889
rect 2050 12855 2056 12889
rect 1837 12814 1946 12855
rect 2048 12814 2056 12855
rect 1837 12780 1944 12814
rect 2050 12780 2056 12814
rect 1837 12739 1946 12780
rect 2048 12739 2056 12780
rect 1837 12705 1944 12739
rect 2050 12705 2056 12739
rect 1837 12664 1946 12705
rect 2048 12664 2056 12705
rect 1837 12630 1944 12664
rect 2050 12630 2056 12664
rect 1837 12589 1946 12630
rect 2048 12589 2056 12630
rect 1837 12555 1944 12589
rect 2050 12555 2056 12589
rect 1837 12514 1946 12555
rect 2048 12514 2056 12555
rect 1837 12480 1944 12514
rect 2050 12480 2056 12514
rect 1837 12439 1946 12480
rect 2048 12439 2056 12480
rect 1837 12405 1944 12439
rect 2050 12405 2056 12439
rect 1837 12364 1946 12405
rect 2048 12364 2056 12405
rect 1837 12330 1944 12364
rect 2050 12330 2056 12364
rect 1837 12289 1946 12330
rect 2048 12289 2056 12330
rect 1837 12255 1944 12289
rect 2050 12255 2056 12289
rect 1837 12214 1946 12255
rect 2048 12214 2056 12255
rect 1837 12180 1944 12214
rect 2050 12180 2056 12214
rect 1837 12139 1946 12180
rect 2048 12139 2056 12180
rect 1837 12105 1944 12139
rect 2050 12105 2056 12139
rect 1837 12064 1946 12105
rect 2048 12064 2056 12105
rect 1837 12030 1944 12064
rect 2050 12030 2056 12064
rect 1837 11989 1946 12030
rect 2048 11989 2056 12030
rect 1837 11955 1944 11989
rect 2050 11955 2056 11989
rect 1837 11914 1946 11955
rect 2048 11914 2056 11955
rect 1837 11880 1944 11914
rect 2050 11880 2056 11914
rect 1837 11839 1946 11880
rect 2048 11839 2056 11880
rect 1837 11805 1944 11839
rect 2050 11805 2056 11839
rect 1837 11764 1946 11805
rect 2048 11764 2056 11805
rect 1837 11730 1944 11764
rect 2050 11730 2056 11764
rect 1837 11689 1946 11730
rect 2048 11689 2056 11730
rect 1837 11655 1944 11689
rect 2050 11655 2056 11689
rect 1837 11614 1946 11655
rect 2048 11614 2056 11655
rect 1837 11580 1944 11614
rect 2050 11580 2056 11614
rect 1837 11539 1946 11580
rect 2048 11539 2056 11580
rect 1837 11505 1944 11539
rect 2050 11505 2056 11539
rect 1837 11464 1946 11505
rect 2048 11464 2056 11505
rect 1837 11430 1944 11464
rect 2050 11430 2056 11464
rect 1837 11389 1946 11430
rect 2048 11389 2056 11430
rect 1837 11355 1944 11389
rect 2050 11355 2056 11389
rect 1837 11313 1946 11355
rect 2048 11313 2056 11355
rect 1837 11279 1944 11313
rect 2050 11279 2056 11313
rect 1837 10847 1946 11279
rect 2048 10847 2056 11279
rect 1837 10813 1944 10847
rect 2050 10813 2056 10847
rect 1837 10771 1946 10813
rect 2048 10771 2056 10813
rect 1837 10737 1944 10771
rect 2050 10737 2056 10771
rect 1837 10695 1946 10737
rect 2048 10695 2056 10737
rect 1837 10661 1944 10695
rect 2050 10661 2056 10695
rect 1837 10620 1946 10661
rect 2048 10620 2056 10661
rect 1837 10586 1944 10620
rect 2050 10586 2056 10620
rect 1837 10545 1946 10586
rect 2048 10545 2056 10586
rect 1837 10511 1944 10545
rect 2050 10511 2056 10545
rect 1837 10470 1946 10511
rect 2048 10470 2056 10511
rect 1837 10436 1944 10470
rect 2050 10436 2056 10470
rect 1837 10395 1946 10436
rect 2048 10395 2056 10436
rect 1837 10361 1944 10395
rect 2050 10361 2056 10395
rect 1837 10320 1946 10361
rect 2048 10320 2056 10361
rect 1837 10286 1944 10320
rect 2050 10286 2056 10320
rect 1837 10245 1946 10286
rect 2048 10245 2056 10286
rect 1837 10211 1944 10245
rect 2050 10211 2056 10245
rect 1837 10170 1946 10211
rect 2048 10170 2056 10211
rect 1837 10136 1944 10170
rect 2050 10136 2056 10170
rect 1837 10095 1946 10136
rect 2048 10095 2056 10136
rect 1837 10061 1944 10095
rect 2050 10061 2056 10095
rect 1837 10020 1946 10061
rect 2048 10020 2056 10061
rect 1837 9986 1944 10020
rect 2050 9986 2056 10020
rect 1837 9945 1946 9986
rect 2048 9945 2056 9986
rect 1837 9911 1944 9945
rect 2050 9911 2056 9945
rect 1837 9870 1946 9911
rect 2048 9870 2056 9911
rect 1837 9836 1944 9870
rect 2050 9836 2056 9870
rect 1837 9795 1946 9836
rect 2048 9795 2056 9836
rect 1837 9761 1944 9795
rect 2050 9761 2056 9795
rect 1837 9720 1946 9761
rect 2048 9720 2056 9761
rect 1837 9686 1944 9720
rect 2050 9686 2056 9720
rect 1837 9645 1946 9686
rect 2048 9645 2056 9686
rect 1837 9611 1944 9645
rect 2050 9611 2056 9645
rect 1837 9570 1946 9611
rect 2048 9570 2056 9611
rect 1837 9536 1944 9570
rect 2050 9536 2056 9570
rect 1837 9495 1946 9536
rect 2048 9495 2056 9536
rect 1837 9461 1944 9495
rect 2050 9461 2056 9495
rect 1837 9420 1946 9461
rect 2048 9420 2056 9461
rect 1837 9386 1944 9420
rect 2050 9386 2056 9420
rect 1837 8732 1946 9386
rect 2048 8732 2056 9386
rect 2255 16383 2514 16417
rect 4588 16387 4622 16417
rect 2255 12789 2274 16383
rect 2444 16315 2514 16383
rect 4588 16315 4656 16387
rect 2595 16209 2615 16243
rect 2649 16209 2683 16243
rect 2717 16209 2751 16243
rect 2785 16209 2819 16243
rect 2853 16209 2887 16243
rect 2921 16209 2955 16243
rect 2989 16209 3023 16243
rect 3057 16209 3091 16243
rect 3125 16209 3159 16243
rect 3193 16209 3227 16243
rect 3261 16209 3295 16243
rect 3329 16209 3363 16243
rect 3397 16209 3431 16243
rect 3465 16209 3499 16243
rect 3533 16209 3567 16243
rect 3601 16209 3635 16243
rect 3669 16209 3703 16243
rect 3737 16209 3771 16243
rect 3805 16209 3839 16243
rect 3873 16209 3907 16243
rect 3941 16209 3975 16243
rect 4009 16209 4043 16243
rect 4077 16209 4111 16243
rect 4145 16209 4179 16243
rect 4213 16209 4247 16243
rect 4281 16209 4315 16243
rect 4349 16209 4383 16243
rect 4417 16209 4451 16243
rect 4485 16209 4519 16243
rect 4553 16209 4587 16243
rect 4621 16209 4655 16243
rect 4689 16209 4723 16243
rect 4757 16209 4791 16243
rect 4825 16209 4859 16243
rect 4893 16209 4923 16243
rect 4961 16209 4995 16243
rect 5030 16209 5063 16243
rect 5103 16209 5131 16243
rect 5176 16209 5199 16243
rect 5249 16209 5267 16243
rect 5322 16209 5335 16243
rect 5395 16209 5403 16243
rect 5468 16209 5471 16243
rect 5505 16209 5507 16243
rect 5573 16209 5580 16243
rect 5641 16209 5653 16243
rect 5709 16209 5726 16243
rect 5777 16209 5799 16243
rect 5845 16209 5872 16243
rect 5913 16209 5945 16243
rect 5981 16209 6015 16243
rect 6051 16209 6083 16243
rect 6123 16209 6151 16243
rect 6195 16209 6219 16243
rect 6267 16209 6287 16243
rect 6339 16209 6355 16243
rect 6411 16209 6423 16243
rect 6483 16209 6491 16243
rect 6555 16209 6559 16243
rect 6661 16209 6665 16243
rect 6729 16209 6737 16243
rect 6797 16209 6809 16243
rect 6865 16209 6881 16243
rect 6933 16209 6953 16243
rect 7001 16209 7025 16243
rect 7069 16209 7097 16243
rect 7137 16209 7169 16243
rect 7205 16209 7239 16243
rect 7275 16209 7307 16243
rect 7347 16209 7375 16243
rect 7419 16209 7443 16243
rect 7491 16209 7511 16243
rect 7563 16209 7579 16243
rect 7635 16209 7647 16243
rect 7707 16209 7715 16243
rect 7779 16209 7783 16243
rect 7885 16209 7889 16243
rect 7953 16209 7961 16243
rect 8021 16209 8033 16243
rect 8089 16209 8105 16243
rect 8157 16209 8177 16243
rect 8225 16209 8249 16243
rect 8293 16209 8321 16243
rect 8361 16209 8393 16243
rect 8429 16209 8463 16243
rect 8499 16209 8531 16243
rect 8571 16209 8599 16243
rect 8643 16209 8667 16243
rect 8715 16209 8735 16243
rect 8787 16209 8803 16243
rect 8859 16209 8871 16243
rect 8931 16209 8939 16243
rect 9003 16209 9007 16243
rect 9109 16209 9113 16243
rect 9177 16209 9185 16243
rect 9245 16209 9257 16243
rect 9313 16209 9329 16243
rect 9381 16209 9401 16243
rect 9449 16209 9473 16243
rect 9517 16209 9545 16243
rect 9585 16209 9617 16243
rect 9653 16209 9687 16243
rect 9723 16209 9755 16243
rect 9795 16209 9823 16243
rect 9867 16209 9891 16243
rect 9939 16209 9959 16243
rect 10011 16209 10027 16243
rect 10083 16209 10095 16243
rect 10155 16209 10163 16243
rect 10227 16209 10231 16243
rect 10333 16209 10337 16243
rect 10401 16209 10409 16243
rect 10469 16209 10481 16243
rect 10537 16209 10553 16243
rect 10605 16209 10625 16243
rect 10673 16209 10697 16243
rect 10741 16209 10769 16243
rect 10809 16209 10841 16243
rect 10877 16209 10911 16243
rect 10947 16209 10979 16243
rect 11019 16209 11047 16243
rect 11091 16209 11115 16243
rect 11163 16209 11183 16243
rect 11235 16209 11251 16243
rect 11307 16209 11319 16243
rect 11379 16209 11387 16243
rect 11451 16209 11455 16243
rect 11557 16209 11561 16243
rect 11625 16209 11633 16243
rect 11693 16209 11705 16243
rect 11761 16209 11777 16243
rect 11829 16209 11849 16243
rect 11897 16209 11921 16243
rect 11965 16209 11993 16243
rect 12033 16209 12065 16243
rect 12101 16209 12135 16243
rect 12171 16209 12203 16243
rect 12243 16209 12271 16243
rect 12315 16209 12339 16243
rect 12387 16209 12407 16243
rect 12459 16209 12475 16243
rect 12531 16209 12543 16243
rect 12603 16209 12611 16243
rect 12675 16209 12679 16243
rect 12781 16209 12785 16243
rect 12849 16209 12857 16243
rect 12917 16209 12929 16243
rect 12985 16209 13019 16243
rect 13053 16209 13087 16243
rect 13121 16209 13155 16243
rect 13189 16209 13223 16243
rect 13257 16209 13331 16243
rect 2550 15987 2584 16026
rect 2550 15914 2584 15953
rect 2550 15841 2584 15880
rect 2550 15768 2584 15807
rect 2550 15695 2584 15734
rect 2550 15623 2584 15661
rect 2550 15551 2584 15589
rect 2550 15479 2584 15517
rect 2550 15407 2584 15445
rect 2550 15335 2584 15373
rect 2550 15263 2584 15301
rect 2550 15191 2584 15229
rect 3406 15987 3440 16026
rect 3406 15914 3440 15953
rect 3406 15841 3440 15880
rect 3406 15768 3440 15807
rect 3406 15695 3440 15734
rect 3406 15623 3440 15661
rect 3406 15551 3440 15589
rect 3406 15479 3440 15517
rect 3406 15407 3440 15445
rect 3406 15335 3440 15373
rect 3406 15263 3440 15301
rect 3406 15191 3440 15229
rect 5062 15987 5096 16026
rect 5062 15914 5096 15953
rect 5062 15841 5096 15880
rect 5062 15768 5096 15807
rect 5062 15695 5096 15734
rect 5062 15623 5096 15661
rect 5062 15551 5096 15589
rect 5062 15479 5096 15517
rect 5062 15407 5096 15445
rect 5062 15335 5096 15373
rect 5062 15263 5096 15301
rect 5062 15191 5096 15229
rect 6718 15987 6752 16026
rect 6718 15914 6752 15953
rect 6718 15841 6752 15880
rect 6718 15768 6752 15807
rect 6718 15695 6752 15734
rect 6718 15623 6752 15661
rect 6718 15551 6752 15589
rect 6718 15479 6752 15517
rect 6718 15407 6752 15445
rect 6718 15335 6752 15373
rect 6718 15263 6752 15301
rect 6718 15191 6752 15229
rect 8374 15987 8408 16026
rect 8374 15914 8408 15953
rect 8374 15841 8408 15880
rect 8374 15768 8408 15807
rect 8374 15695 8408 15734
rect 8374 15623 8408 15661
rect 8374 15551 8408 15589
rect 8374 15479 8408 15517
rect 8374 15407 8408 15445
rect 8374 15335 8408 15373
rect 8374 15263 8408 15301
rect 8374 15191 8408 15229
rect 10030 15987 10064 16026
rect 10030 15914 10064 15953
rect 10030 15841 10064 15880
rect 10030 15768 10064 15807
rect 10030 15695 10064 15734
rect 10030 15623 10064 15661
rect 10030 15551 10064 15589
rect 10030 15479 10064 15517
rect 10030 15407 10064 15445
rect 10030 15335 10064 15373
rect 10030 15263 10064 15301
rect 10030 15191 10064 15229
rect 11686 15987 11720 16026
rect 11686 15914 11720 15953
rect 11686 15841 11720 15880
rect 11686 15768 11720 15807
rect 11686 15695 11720 15734
rect 11686 15623 11720 15661
rect 11686 15551 11720 15589
rect 11686 15479 11720 15517
rect 11686 15407 11720 15445
rect 11686 15335 11720 15373
rect 11686 15263 11720 15301
rect 11686 15191 11720 15229
rect 13342 16030 13376 16073
rect 13342 15953 13376 15996
rect 13342 15876 13376 15919
rect 13342 15799 13376 15842
rect 13342 15723 13376 15765
rect 13342 15647 13376 15689
rect 13342 15571 13376 15613
rect 13342 15495 13376 15537
rect 13342 15419 13376 15461
rect 13342 15343 13376 15385
rect 13342 15267 13376 15309
rect 13342 15191 13376 15233
rect 2713 14311 2751 14345
rect 2679 14267 2785 14311
rect 2713 14233 2751 14267
rect 2679 14189 2785 14233
rect 2713 14155 2751 14189
rect 2679 14111 2785 14155
rect 2713 14077 2751 14111
rect 2679 14033 2785 14077
rect 2713 13999 2751 14033
rect 2679 13955 2785 13999
rect 2713 13921 2751 13955
rect 2679 13877 2785 13921
rect 2713 13843 2751 13877
rect 2679 13799 2785 13843
rect 2713 13765 2751 13799
rect 2679 13722 2785 13765
rect 2713 13688 2751 13722
rect 2679 13645 2785 13688
rect 2713 13611 2751 13645
rect 2679 13568 2785 13611
rect 2713 13534 2751 13568
rect 2679 13491 2785 13534
rect 2713 13457 2751 13491
rect 2679 13414 2785 13457
rect 2713 13380 2751 13414
rect 2990 14311 3028 14345
rect 2956 14267 3062 14311
rect 2990 14233 3028 14267
rect 2956 14189 3062 14233
rect 2990 14155 3028 14189
rect 2956 14111 3062 14155
rect 2990 14077 3028 14111
rect 2956 14033 3062 14077
rect 2990 13999 3028 14033
rect 2956 13955 3062 13999
rect 2990 13921 3028 13955
rect 2956 13877 3062 13921
rect 2990 13843 3028 13877
rect 2956 13799 3062 13843
rect 2990 13765 3028 13799
rect 2956 13722 3062 13765
rect 2990 13688 3028 13722
rect 2956 13645 3062 13688
rect 2990 13611 3028 13645
rect 2956 13568 3062 13611
rect 2990 13534 3028 13568
rect 2956 13491 3062 13534
rect 2990 13457 3028 13491
rect 2956 13414 3062 13457
rect 2990 13380 3028 13414
rect 3267 14311 3305 14345
rect 3233 14267 3339 14311
rect 3267 14233 3305 14267
rect 3233 14189 3339 14233
rect 3267 14155 3305 14189
rect 3233 14111 3339 14155
rect 3267 14077 3305 14111
rect 3233 14033 3339 14077
rect 3267 13999 3305 14033
rect 3233 13955 3339 13999
rect 3267 13921 3305 13955
rect 3233 13877 3339 13921
rect 3267 13843 3305 13877
rect 3233 13799 3339 13843
rect 3267 13765 3305 13799
rect 3233 13722 3339 13765
rect 3267 13688 3305 13722
rect 3233 13645 3339 13688
rect 3267 13611 3305 13645
rect 3233 13568 3339 13611
rect 3267 13534 3305 13568
rect 3233 13491 3339 13534
rect 3267 13457 3305 13491
rect 3233 13414 3339 13457
rect 3267 13380 3305 13414
rect 3544 14311 3582 14345
rect 3510 14267 3616 14311
rect 3544 14233 3582 14267
rect 3510 14189 3616 14233
rect 3544 14155 3582 14189
rect 3510 14111 3616 14155
rect 3544 14077 3582 14111
rect 3510 14033 3616 14077
rect 3544 13999 3582 14033
rect 3510 13955 3616 13999
rect 3544 13921 3582 13955
rect 3510 13877 3616 13921
rect 3544 13843 3582 13877
rect 3510 13799 3616 13843
rect 3544 13765 3582 13799
rect 3510 13722 3616 13765
rect 3544 13688 3582 13722
rect 3510 13645 3616 13688
rect 3544 13611 3582 13645
rect 3510 13568 3616 13611
rect 3544 13534 3582 13568
rect 3510 13491 3616 13534
rect 3544 13457 3582 13491
rect 3510 13414 3616 13457
rect 3544 13380 3582 13414
rect 3821 14311 3859 14345
rect 3787 14267 3893 14311
rect 3821 14233 3859 14267
rect 3787 14189 3893 14233
rect 3821 14155 3859 14189
rect 3787 14111 3893 14155
rect 3821 14077 3859 14111
rect 3787 14033 3893 14077
rect 3821 13999 3859 14033
rect 3787 13955 3893 13999
rect 3821 13921 3859 13955
rect 3787 13877 3893 13921
rect 3821 13843 3859 13877
rect 3787 13799 3893 13843
rect 3821 13765 3859 13799
rect 3787 13722 3893 13765
rect 3821 13688 3859 13722
rect 3787 13645 3893 13688
rect 3821 13611 3859 13645
rect 3787 13568 3893 13611
rect 3821 13534 3859 13568
rect 3787 13491 3893 13534
rect 3821 13457 3859 13491
rect 3787 13414 3893 13457
rect 3821 13380 3859 13414
rect 4098 14311 4136 14345
rect 4064 14267 4170 14311
rect 4098 14233 4136 14267
rect 4064 14189 4170 14233
rect 4098 14155 4136 14189
rect 4064 14111 4170 14155
rect 4098 14077 4136 14111
rect 4064 14033 4170 14077
rect 4098 13999 4136 14033
rect 4064 13955 4170 13999
rect 4098 13921 4136 13955
rect 4064 13877 4170 13921
rect 4098 13843 4136 13877
rect 4064 13799 4170 13843
rect 4098 13765 4136 13799
rect 4064 13722 4170 13765
rect 4098 13688 4136 13722
rect 4064 13645 4170 13688
rect 4098 13611 4136 13645
rect 4064 13568 4170 13611
rect 4098 13534 4136 13568
rect 4064 13491 4170 13534
rect 4098 13457 4136 13491
rect 4064 13414 4170 13457
rect 4098 13380 4136 13414
rect 4375 14311 4413 14345
rect 4341 14267 4447 14311
rect 4375 14233 4413 14267
rect 4341 14189 4447 14233
rect 4375 14155 4413 14189
rect 4341 14111 4447 14155
rect 4375 14077 4413 14111
rect 4341 14033 4447 14077
rect 4375 13999 4413 14033
rect 4341 13955 4447 13999
rect 4375 13921 4413 13955
rect 4341 13877 4447 13921
rect 4375 13843 4413 13877
rect 4341 13799 4447 13843
rect 4375 13765 4413 13799
rect 4341 13722 4447 13765
rect 4375 13688 4413 13722
rect 4341 13645 4447 13688
rect 4375 13611 4413 13645
rect 4341 13568 4447 13611
rect 4375 13534 4413 13568
rect 4341 13491 4447 13534
rect 4375 13457 4413 13491
rect 4341 13414 4447 13457
rect 4375 13380 4413 13414
rect 4652 14311 4690 14345
rect 4618 14267 4724 14311
rect 4652 14233 4690 14267
rect 4618 14189 4724 14233
rect 4652 14155 4690 14189
rect 4618 14111 4724 14155
rect 4652 14077 4690 14111
rect 4618 14033 4724 14077
rect 4652 13999 4690 14033
rect 4618 13955 4724 13999
rect 4652 13921 4690 13955
rect 4618 13877 4724 13921
rect 4652 13843 4690 13877
rect 4618 13799 4724 13843
rect 4652 13765 4690 13799
rect 4618 13722 4724 13765
rect 4652 13688 4690 13722
rect 4618 13645 4724 13688
rect 4652 13611 4690 13645
rect 4618 13568 4724 13611
rect 4652 13534 4690 13568
rect 4618 13491 4724 13534
rect 4652 13457 4690 13491
rect 4618 13414 4724 13457
rect 4652 13380 4690 13414
rect 4929 14311 4967 14345
rect 4895 14267 5001 14311
rect 4929 14233 4967 14267
rect 4895 14189 5001 14233
rect 4929 14155 4967 14189
rect 4895 14111 5001 14155
rect 4929 14077 4967 14111
rect 4895 14033 5001 14077
rect 4929 13999 4967 14033
rect 4895 13955 5001 13999
rect 4929 13921 4967 13955
rect 4895 13877 5001 13921
rect 4929 13843 4967 13877
rect 4895 13799 5001 13843
rect 4929 13765 4967 13799
rect 4895 13722 5001 13765
rect 4929 13688 4967 13722
rect 4895 13645 5001 13688
rect 4929 13611 4967 13645
rect 4895 13568 5001 13611
rect 4929 13534 4967 13568
rect 4895 13491 5001 13534
rect 4929 13457 4967 13491
rect 4895 13414 5001 13457
rect 4929 13380 4967 13414
rect 5206 14311 5244 14345
rect 5172 14267 5278 14311
rect 5206 14233 5244 14267
rect 5172 14189 5278 14233
rect 5206 14155 5244 14189
rect 5172 14111 5278 14155
rect 5206 14077 5244 14111
rect 5172 14033 5278 14077
rect 5206 13999 5244 14033
rect 5172 13955 5278 13999
rect 5206 13921 5244 13955
rect 5172 13877 5278 13921
rect 5206 13843 5244 13877
rect 5172 13799 5278 13843
rect 5206 13765 5244 13799
rect 5172 13722 5278 13765
rect 5206 13688 5244 13722
rect 5172 13645 5278 13688
rect 5206 13611 5244 13645
rect 5172 13568 5278 13611
rect 5206 13534 5244 13568
rect 5172 13491 5278 13534
rect 5206 13457 5244 13491
rect 5172 13414 5278 13457
rect 5206 13380 5244 13414
rect 5483 14311 5521 14345
rect 5449 14267 5555 14311
rect 5483 14233 5521 14267
rect 5449 14189 5555 14233
rect 5483 14155 5521 14189
rect 5449 14111 5555 14155
rect 5483 14077 5521 14111
rect 5449 14033 5555 14077
rect 5483 13999 5521 14033
rect 5449 13955 5555 13999
rect 5483 13921 5521 13955
rect 5449 13877 5555 13921
rect 5483 13843 5521 13877
rect 5449 13799 5555 13843
rect 5483 13765 5521 13799
rect 5449 13722 5555 13765
rect 5483 13688 5521 13722
rect 5449 13645 5555 13688
rect 5483 13611 5521 13645
rect 5449 13568 5555 13611
rect 5483 13534 5521 13568
rect 5449 13491 5555 13534
rect 5483 13457 5521 13491
rect 5449 13414 5555 13457
rect 5483 13380 5521 13414
rect 5760 14311 5798 14345
rect 5726 14267 5832 14311
rect 5760 14233 5798 14267
rect 5726 14189 5832 14233
rect 5760 14155 5798 14189
rect 5726 14111 5832 14155
rect 5760 14077 5798 14111
rect 5726 14033 5832 14077
rect 5760 13999 5798 14033
rect 5726 13955 5832 13999
rect 5760 13921 5798 13955
rect 5726 13877 5832 13921
rect 5760 13843 5798 13877
rect 5726 13799 5832 13843
rect 5760 13765 5798 13799
rect 5726 13722 5832 13765
rect 5760 13688 5798 13722
rect 5726 13645 5832 13688
rect 5760 13611 5798 13645
rect 5726 13568 5832 13611
rect 5760 13534 5798 13568
rect 5726 13491 5832 13534
rect 5760 13457 5798 13491
rect 5726 13414 5832 13457
rect 5760 13380 5798 13414
rect 6037 14311 6075 14345
rect 6003 14267 6109 14311
rect 6037 14233 6075 14267
rect 6003 14189 6109 14233
rect 6037 14155 6075 14189
rect 6003 14111 6109 14155
rect 6037 14077 6075 14111
rect 6003 14033 6109 14077
rect 6037 13999 6075 14033
rect 6003 13955 6109 13999
rect 6037 13921 6075 13955
rect 6003 13877 6109 13921
rect 6037 13843 6075 13877
rect 6003 13799 6109 13843
rect 6037 13765 6075 13799
rect 6003 13722 6109 13765
rect 6037 13688 6075 13722
rect 6003 13645 6109 13688
rect 6037 13611 6075 13645
rect 6003 13568 6109 13611
rect 6037 13534 6075 13568
rect 6003 13491 6109 13534
rect 6037 13457 6075 13491
rect 6003 13414 6109 13457
rect 6037 13380 6075 13414
rect 6314 14311 6352 14345
rect 6280 14267 6386 14311
rect 6314 14233 6352 14267
rect 6280 14189 6386 14233
rect 6314 14155 6352 14189
rect 6280 14111 6386 14155
rect 6314 14077 6352 14111
rect 6280 14033 6386 14077
rect 6314 13999 6352 14033
rect 6280 13955 6386 13999
rect 6314 13921 6352 13955
rect 6280 13877 6386 13921
rect 6314 13843 6352 13877
rect 6280 13799 6386 13843
rect 6314 13765 6352 13799
rect 6280 13722 6386 13765
rect 6314 13688 6352 13722
rect 6280 13645 6386 13688
rect 6314 13611 6352 13645
rect 6280 13568 6386 13611
rect 6314 13534 6352 13568
rect 6280 13491 6386 13534
rect 6314 13457 6352 13491
rect 6280 13414 6386 13457
rect 6314 13380 6352 13414
rect 6591 14311 6629 14345
rect 6557 14267 6663 14311
rect 6591 14233 6629 14267
rect 6557 14189 6663 14233
rect 6591 14155 6629 14189
rect 6557 14111 6663 14155
rect 6591 14077 6629 14111
rect 6557 14033 6663 14077
rect 6591 13999 6629 14033
rect 6557 13955 6663 13999
rect 6591 13921 6629 13955
rect 6557 13877 6663 13921
rect 6591 13843 6629 13877
rect 6557 13799 6663 13843
rect 6591 13765 6629 13799
rect 6557 13722 6663 13765
rect 6591 13688 6629 13722
rect 6557 13645 6663 13688
rect 6591 13611 6629 13645
rect 6557 13568 6663 13611
rect 6591 13534 6629 13568
rect 6557 13491 6663 13534
rect 6591 13457 6629 13491
rect 6557 13414 6663 13457
rect 6591 13380 6629 13414
rect 6868 14311 6906 14345
rect 6834 14267 6940 14311
rect 6868 14233 6906 14267
rect 6834 14189 6940 14233
rect 6868 14155 6906 14189
rect 6834 14111 6940 14155
rect 6868 14077 6906 14111
rect 6834 14033 6940 14077
rect 6868 13999 6906 14033
rect 6834 13955 6940 13999
rect 6868 13921 6906 13955
rect 6834 13877 6940 13921
rect 6868 13843 6906 13877
rect 6834 13799 6940 13843
rect 6868 13765 6906 13799
rect 6834 13722 6940 13765
rect 6868 13688 6906 13722
rect 6834 13645 6940 13688
rect 6868 13611 6906 13645
rect 6834 13568 6940 13611
rect 6868 13534 6906 13568
rect 6834 13491 6940 13534
rect 6868 13457 6906 13491
rect 6834 13414 6940 13457
rect 6868 13380 6906 13414
rect 7145 14311 7183 14345
rect 7111 14267 7217 14311
rect 7145 14233 7183 14267
rect 7111 14189 7217 14233
rect 7145 14155 7183 14189
rect 7111 14111 7217 14155
rect 7145 14077 7183 14111
rect 7111 14033 7217 14077
rect 7145 13999 7183 14033
rect 7111 13955 7217 13999
rect 7145 13921 7183 13955
rect 7111 13877 7217 13921
rect 7145 13843 7183 13877
rect 7111 13799 7217 13843
rect 7145 13765 7183 13799
rect 7111 13722 7217 13765
rect 7145 13688 7183 13722
rect 7111 13645 7217 13688
rect 7145 13611 7183 13645
rect 7111 13568 7217 13611
rect 7145 13534 7183 13568
rect 7111 13491 7217 13534
rect 7145 13457 7183 13491
rect 7111 13414 7217 13457
rect 7145 13380 7183 13414
rect 7422 14311 7460 14345
rect 7388 14267 7494 14311
rect 7422 14233 7460 14267
rect 7388 14189 7494 14233
rect 7422 14155 7460 14189
rect 7388 14111 7494 14155
rect 7422 14077 7460 14111
rect 7388 14033 7494 14077
rect 7422 13999 7460 14033
rect 7388 13955 7494 13999
rect 7422 13921 7460 13955
rect 7388 13877 7494 13921
rect 7422 13843 7460 13877
rect 7388 13799 7494 13843
rect 7422 13765 7460 13799
rect 7388 13722 7494 13765
rect 7422 13688 7460 13722
rect 7388 13645 7494 13688
rect 7422 13611 7460 13645
rect 7388 13568 7494 13611
rect 7422 13534 7460 13568
rect 7388 13491 7494 13534
rect 7422 13457 7460 13491
rect 7388 13414 7494 13457
rect 7422 13380 7460 13414
rect 7699 14311 7737 14345
rect 7665 14267 7771 14311
rect 7699 14233 7737 14267
rect 7665 14189 7771 14233
rect 7699 14155 7737 14189
rect 7665 14111 7771 14155
rect 7699 14077 7737 14111
rect 7665 14033 7771 14077
rect 7699 13999 7737 14033
rect 7665 13955 7771 13999
rect 7699 13921 7737 13955
rect 7665 13877 7771 13921
rect 7699 13843 7737 13877
rect 7665 13799 7771 13843
rect 7699 13765 7737 13799
rect 7665 13722 7771 13765
rect 7699 13688 7737 13722
rect 7665 13645 7771 13688
rect 7699 13611 7737 13645
rect 7665 13568 7771 13611
rect 7699 13534 7737 13568
rect 7665 13491 7771 13534
rect 7699 13457 7737 13491
rect 7665 13414 7771 13457
rect 7699 13380 7737 13414
rect 7976 14311 8014 14345
rect 7942 14267 8048 14311
rect 7976 14233 8014 14267
rect 7942 14189 8048 14233
rect 7976 14155 8014 14189
rect 7942 14111 8048 14155
rect 7976 14077 8014 14111
rect 7942 14033 8048 14077
rect 7976 13999 8014 14033
rect 7942 13955 8048 13999
rect 7976 13921 8014 13955
rect 7942 13877 8048 13921
rect 7976 13843 8014 13877
rect 7942 13799 8048 13843
rect 7976 13765 8014 13799
rect 7942 13722 8048 13765
rect 7976 13688 8014 13722
rect 7942 13645 8048 13688
rect 7976 13611 8014 13645
rect 7942 13568 8048 13611
rect 7976 13534 8014 13568
rect 7942 13491 8048 13534
rect 7976 13457 8014 13491
rect 7942 13414 8048 13457
rect 7976 13380 8014 13414
rect 8253 14311 8291 14345
rect 8219 14267 8325 14311
rect 8253 14233 8291 14267
rect 8219 14189 8325 14233
rect 8253 14155 8291 14189
rect 8219 14111 8325 14155
rect 8253 14077 8291 14111
rect 8219 14033 8325 14077
rect 8253 13999 8291 14033
rect 8219 13955 8325 13999
rect 8253 13921 8291 13955
rect 8219 13877 8325 13921
rect 8253 13843 8291 13877
rect 8219 13799 8325 13843
rect 8253 13765 8291 13799
rect 8219 13722 8325 13765
rect 8253 13688 8291 13722
rect 8219 13645 8325 13688
rect 8253 13611 8291 13645
rect 8219 13568 8325 13611
rect 8253 13534 8291 13568
rect 8219 13491 8325 13534
rect 8253 13457 8291 13491
rect 8219 13414 8325 13457
rect 8253 13380 8291 13414
rect 8530 14311 8568 14345
rect 8496 14267 8602 14311
rect 8530 14233 8568 14267
rect 8496 14189 8602 14233
rect 8530 14155 8568 14189
rect 8496 14111 8602 14155
rect 8530 14077 8568 14111
rect 8496 14033 8602 14077
rect 8530 13999 8568 14033
rect 8496 13955 8602 13999
rect 8530 13921 8568 13955
rect 8496 13877 8602 13921
rect 8530 13843 8568 13877
rect 8496 13799 8602 13843
rect 8530 13765 8568 13799
rect 8496 13722 8602 13765
rect 8530 13688 8568 13722
rect 8496 13645 8602 13688
rect 8530 13611 8568 13645
rect 8496 13568 8602 13611
rect 8530 13534 8568 13568
rect 8496 13491 8602 13534
rect 8530 13457 8568 13491
rect 8496 13414 8602 13457
rect 8530 13380 8568 13414
rect 8807 14311 8845 14345
rect 8773 14267 8879 14311
rect 8807 14233 8845 14267
rect 8773 14189 8879 14233
rect 8807 14155 8845 14189
rect 8773 14111 8879 14155
rect 8807 14077 8845 14111
rect 8773 14033 8879 14077
rect 8807 13999 8845 14033
rect 8773 13955 8879 13999
rect 8807 13921 8845 13955
rect 8773 13877 8879 13921
rect 8807 13843 8845 13877
rect 8773 13799 8879 13843
rect 8807 13765 8845 13799
rect 8773 13722 8879 13765
rect 8807 13688 8845 13722
rect 8773 13645 8879 13688
rect 8807 13611 8845 13645
rect 8773 13568 8879 13611
rect 8807 13534 8845 13568
rect 8773 13491 8879 13534
rect 8807 13457 8845 13491
rect 8773 13414 8879 13457
rect 8807 13380 8845 13414
rect 9084 14311 9122 14345
rect 9050 14267 9156 14311
rect 9084 14233 9122 14267
rect 9050 14189 9156 14233
rect 9084 14155 9122 14189
rect 9050 14111 9156 14155
rect 9084 14077 9122 14111
rect 9050 14033 9156 14077
rect 9084 13999 9122 14033
rect 9050 13955 9156 13999
rect 9084 13921 9122 13955
rect 9050 13877 9156 13921
rect 9084 13843 9122 13877
rect 9050 13799 9156 13843
rect 9084 13765 9122 13799
rect 9050 13722 9156 13765
rect 9084 13688 9122 13722
rect 9050 13645 9156 13688
rect 9084 13611 9122 13645
rect 9050 13568 9156 13611
rect 9084 13534 9122 13568
rect 9050 13491 9156 13534
rect 9084 13457 9122 13491
rect 9050 13414 9156 13457
rect 9084 13380 9122 13414
rect 9361 14311 9399 14345
rect 9327 14267 9433 14311
rect 9361 14233 9399 14267
rect 9327 14189 9433 14233
rect 9361 14155 9399 14189
rect 9327 14111 9433 14155
rect 9361 14077 9399 14111
rect 9327 14033 9433 14077
rect 9361 13999 9399 14033
rect 9327 13955 9433 13999
rect 9361 13921 9399 13955
rect 9327 13877 9433 13921
rect 9361 13843 9399 13877
rect 9327 13799 9433 13843
rect 9361 13765 9399 13799
rect 9327 13722 9433 13765
rect 9361 13688 9399 13722
rect 9327 13645 9433 13688
rect 9361 13611 9399 13645
rect 9327 13568 9433 13611
rect 9361 13534 9399 13568
rect 9327 13491 9433 13534
rect 9361 13457 9399 13491
rect 9327 13414 9433 13457
rect 9361 13380 9399 13414
rect 9638 14311 9676 14345
rect 9604 14267 9710 14311
rect 9638 14233 9676 14267
rect 9604 14189 9710 14233
rect 9638 14155 9676 14189
rect 9604 14111 9710 14155
rect 9638 14077 9676 14111
rect 9604 14033 9710 14077
rect 9638 13999 9676 14033
rect 9604 13955 9710 13999
rect 9638 13921 9676 13955
rect 9604 13877 9710 13921
rect 9638 13843 9676 13877
rect 9604 13799 9710 13843
rect 9638 13765 9676 13799
rect 9604 13722 9710 13765
rect 9638 13688 9676 13722
rect 9604 13645 9710 13688
rect 9638 13611 9676 13645
rect 9604 13568 9710 13611
rect 9638 13534 9676 13568
rect 9604 13491 9710 13534
rect 9638 13457 9676 13491
rect 9604 13414 9710 13457
rect 9638 13380 9676 13414
rect 9915 14311 9953 14345
rect 9881 14267 9987 14311
rect 9915 14233 9953 14267
rect 9881 14189 9987 14233
rect 9915 14155 9953 14189
rect 9881 14111 9987 14155
rect 9915 14077 9953 14111
rect 9881 14033 9987 14077
rect 9915 13999 9953 14033
rect 9881 13955 9987 13999
rect 9915 13921 9953 13955
rect 9881 13877 9987 13921
rect 9915 13843 9953 13877
rect 9881 13799 9987 13843
rect 9915 13765 9953 13799
rect 9881 13722 9987 13765
rect 9915 13688 9953 13722
rect 9881 13645 9987 13688
rect 9915 13611 9953 13645
rect 9881 13568 9987 13611
rect 9915 13534 9953 13568
rect 9881 13491 9987 13534
rect 9915 13457 9953 13491
rect 9881 13414 9987 13457
rect 9915 13380 9953 13414
rect 10192 14311 10230 14345
rect 10158 14267 10264 14311
rect 10192 14233 10230 14267
rect 10158 14189 10264 14233
rect 10192 14155 10230 14189
rect 10158 14111 10264 14155
rect 10192 14077 10230 14111
rect 10158 14033 10264 14077
rect 10192 13999 10230 14033
rect 10158 13955 10264 13999
rect 10192 13921 10230 13955
rect 10158 13877 10264 13921
rect 10192 13843 10230 13877
rect 10158 13799 10264 13843
rect 10192 13765 10230 13799
rect 10158 13722 10264 13765
rect 10192 13688 10230 13722
rect 10158 13645 10264 13688
rect 10192 13611 10230 13645
rect 10158 13568 10264 13611
rect 10192 13534 10230 13568
rect 10158 13491 10264 13534
rect 10192 13457 10230 13491
rect 10158 13414 10264 13457
rect 10192 13380 10230 13414
rect 10469 14311 10507 14345
rect 10435 14267 10541 14311
rect 10469 14233 10507 14267
rect 10435 14189 10541 14233
rect 10469 14155 10507 14189
rect 10435 14111 10541 14155
rect 10469 14077 10507 14111
rect 10435 14033 10541 14077
rect 10469 13999 10507 14033
rect 10435 13955 10541 13999
rect 10469 13921 10507 13955
rect 10435 13877 10541 13921
rect 10469 13843 10507 13877
rect 10435 13799 10541 13843
rect 10469 13765 10507 13799
rect 10435 13722 10541 13765
rect 10469 13688 10507 13722
rect 10435 13645 10541 13688
rect 10469 13611 10507 13645
rect 10435 13568 10541 13611
rect 10469 13534 10507 13568
rect 10435 13491 10541 13534
rect 10469 13457 10507 13491
rect 10435 13414 10541 13457
rect 10469 13380 10507 13414
rect 10746 14311 10784 14345
rect 10712 14267 10818 14311
rect 10746 14233 10784 14267
rect 10712 14189 10818 14233
rect 10746 14155 10784 14189
rect 10712 14111 10818 14155
rect 10746 14077 10784 14111
rect 10712 14033 10818 14077
rect 10746 13999 10784 14033
rect 10712 13955 10818 13999
rect 10746 13921 10784 13955
rect 10712 13877 10818 13921
rect 10746 13843 10784 13877
rect 10712 13799 10818 13843
rect 10746 13765 10784 13799
rect 10712 13722 10818 13765
rect 10746 13688 10784 13722
rect 10712 13645 10818 13688
rect 10746 13611 10784 13645
rect 10712 13568 10818 13611
rect 10746 13534 10784 13568
rect 10712 13491 10818 13534
rect 10746 13457 10784 13491
rect 10712 13414 10818 13457
rect 10746 13380 10784 13414
rect 11023 14311 11061 14345
rect 10989 14267 11095 14311
rect 11023 14233 11061 14267
rect 10989 14189 11095 14233
rect 11023 14155 11061 14189
rect 10989 14111 11095 14155
rect 11023 14077 11061 14111
rect 10989 14033 11095 14077
rect 11023 13999 11061 14033
rect 10989 13955 11095 13999
rect 11023 13921 11061 13955
rect 10989 13877 11095 13921
rect 11023 13843 11061 13877
rect 10989 13799 11095 13843
rect 11023 13765 11061 13799
rect 10989 13722 11095 13765
rect 11023 13688 11061 13722
rect 10989 13645 11095 13688
rect 11023 13611 11061 13645
rect 10989 13568 11095 13611
rect 11023 13534 11061 13568
rect 10989 13491 11095 13534
rect 11023 13457 11061 13491
rect 10989 13414 11095 13457
rect 11023 13380 11061 13414
rect 11300 14311 11338 14345
rect 11266 14267 11372 14311
rect 11300 14233 11338 14267
rect 11266 14189 11372 14233
rect 11300 14155 11338 14189
rect 11266 14111 11372 14155
rect 11300 14077 11338 14111
rect 11266 14033 11372 14077
rect 11300 13999 11338 14033
rect 11266 13955 11372 13999
rect 11300 13921 11338 13955
rect 11266 13877 11372 13921
rect 11300 13843 11338 13877
rect 11266 13799 11372 13843
rect 11300 13765 11338 13799
rect 11266 13722 11372 13765
rect 11300 13688 11338 13722
rect 11266 13645 11372 13688
rect 11300 13611 11338 13645
rect 11266 13568 11372 13611
rect 11300 13534 11338 13568
rect 11266 13491 11372 13534
rect 11300 13457 11338 13491
rect 11266 13414 11372 13457
rect 11300 13380 11338 13414
rect 11577 14311 11615 14345
rect 11543 14267 11649 14311
rect 11577 14233 11615 14267
rect 11543 14189 11649 14233
rect 11577 14155 11615 14189
rect 11543 14111 11649 14155
rect 11577 14077 11615 14111
rect 11543 14033 11649 14077
rect 11577 13999 11615 14033
rect 11543 13955 11649 13999
rect 11577 13921 11615 13955
rect 11543 13877 11649 13921
rect 11577 13843 11615 13877
rect 11543 13799 11649 13843
rect 11577 13765 11615 13799
rect 11543 13722 11649 13765
rect 11577 13688 11615 13722
rect 11543 13645 11649 13688
rect 11577 13611 11615 13645
rect 11543 13568 11649 13611
rect 11577 13534 11615 13568
rect 11543 13491 11649 13534
rect 11577 13457 11615 13491
rect 11543 13414 11649 13457
rect 11577 13380 11615 13414
rect 11854 14311 11892 14345
rect 11820 14267 11926 14311
rect 11854 14233 11892 14267
rect 11820 14189 11926 14233
rect 11854 14155 11892 14189
rect 11820 14111 11926 14155
rect 11854 14077 11892 14111
rect 11820 14033 11926 14077
rect 11854 13999 11892 14033
rect 11820 13955 11926 13999
rect 11854 13921 11892 13955
rect 11820 13877 11926 13921
rect 11854 13843 11892 13877
rect 11820 13799 11926 13843
rect 11854 13765 11892 13799
rect 11820 13722 11926 13765
rect 11854 13688 11892 13722
rect 11820 13645 11926 13688
rect 11854 13611 11892 13645
rect 11820 13568 11926 13611
rect 11854 13534 11892 13568
rect 11820 13491 11926 13534
rect 11854 13457 11892 13491
rect 11820 13414 11926 13457
rect 11854 13380 11892 13414
rect 12131 14311 12169 14345
rect 12097 14267 12203 14311
rect 12131 14233 12169 14267
rect 12097 14189 12203 14233
rect 12131 14155 12169 14189
rect 12097 14111 12203 14155
rect 12131 14077 12169 14111
rect 12097 14033 12203 14077
rect 12131 13999 12169 14033
rect 12097 13955 12203 13999
rect 12131 13921 12169 13955
rect 12097 13877 12203 13921
rect 12131 13843 12169 13877
rect 12097 13799 12203 13843
rect 12131 13765 12169 13799
rect 12097 13722 12203 13765
rect 12131 13688 12169 13722
rect 12097 13645 12203 13688
rect 12131 13611 12169 13645
rect 12097 13568 12203 13611
rect 12131 13534 12169 13568
rect 12097 13491 12203 13534
rect 12131 13457 12169 13491
rect 12097 13414 12203 13457
rect 12131 13380 12169 13414
rect 12408 14311 12446 14345
rect 12374 14267 12480 14311
rect 12408 14233 12446 14267
rect 12374 14189 12480 14233
rect 12408 14155 12446 14189
rect 12374 14111 12480 14155
rect 12408 14077 12446 14111
rect 12374 14033 12480 14077
rect 12408 13999 12446 14033
rect 12374 13955 12480 13999
rect 12408 13921 12446 13955
rect 12374 13877 12480 13921
rect 12408 13843 12446 13877
rect 12374 13799 12480 13843
rect 12408 13765 12446 13799
rect 12374 13722 12480 13765
rect 12408 13688 12446 13722
rect 12374 13645 12480 13688
rect 12408 13611 12446 13645
rect 12374 13568 12480 13611
rect 12408 13534 12446 13568
rect 12374 13491 12480 13534
rect 12408 13457 12446 13491
rect 12374 13414 12480 13457
rect 12408 13380 12446 13414
rect 12685 14311 12723 14345
rect 12651 14267 12757 14311
rect 12685 14233 12723 14267
rect 12651 14189 12757 14233
rect 12685 14155 12723 14189
rect 12651 14111 12757 14155
rect 12685 14077 12723 14111
rect 12651 14033 12757 14077
rect 12685 13999 12723 14033
rect 12651 13955 12757 13999
rect 12685 13921 12723 13955
rect 12651 13877 12757 13921
rect 12685 13843 12723 13877
rect 12651 13799 12757 13843
rect 12685 13765 12723 13799
rect 12651 13722 12757 13765
rect 12685 13688 12723 13722
rect 12651 13645 12757 13688
rect 12685 13611 12723 13645
rect 12651 13568 12757 13611
rect 12685 13534 12723 13568
rect 12651 13491 12757 13534
rect 12685 13457 12723 13491
rect 12651 13414 12757 13457
rect 12685 13380 12723 13414
rect 12962 14311 13000 14345
rect 12928 14267 13034 14311
rect 12962 14233 13000 14267
rect 12928 14189 13034 14233
rect 12962 14155 13000 14189
rect 12928 14111 13034 14155
rect 12962 14077 13000 14111
rect 12928 14033 13034 14077
rect 12962 13999 13000 14033
rect 12928 13955 13034 13999
rect 12962 13921 13000 13955
rect 12928 13877 13034 13921
rect 12962 13843 13000 13877
rect 12928 13799 13034 13843
rect 12962 13765 13000 13799
rect 12928 13722 13034 13765
rect 12962 13688 13000 13722
rect 12928 13645 13034 13688
rect 12962 13611 13000 13645
rect 12928 13568 13034 13611
rect 12962 13534 13000 13568
rect 12928 13491 13034 13534
rect 12962 13457 13000 13491
rect 12928 13414 13034 13457
rect 12962 13380 13000 13414
rect 13239 14311 13277 14345
rect 13205 14267 13311 14311
rect 13239 14233 13277 14267
rect 13205 14189 13311 14233
rect 13239 14155 13277 14189
rect 13205 14111 13311 14155
rect 13239 14077 13277 14111
rect 13205 14033 13311 14077
rect 13239 13999 13277 14033
rect 13205 13955 13311 13999
rect 13239 13921 13277 13955
rect 13205 13877 13311 13921
rect 13239 13843 13277 13877
rect 13205 13799 13311 13843
rect 13239 13765 13277 13799
rect 13205 13722 13311 13765
rect 13239 13688 13277 13722
rect 13205 13645 13311 13688
rect 13239 13611 13277 13645
rect 13205 13568 13311 13611
rect 13239 13534 13277 13568
rect 13205 13491 13311 13534
rect 13239 13457 13277 13491
rect 13205 13414 13311 13457
rect 13239 13380 13277 13414
rect 2958 13368 3060 13380
rect 3512 13368 3614 13380
rect 4066 13368 4168 13380
rect 4620 13368 4722 13380
rect 5174 13368 5276 13380
rect 5728 13368 5830 13380
rect 6282 13368 6384 13380
rect 6836 13368 6938 13380
rect 7390 13368 7492 13380
rect 7944 13368 8046 13380
rect 8498 13368 8600 13380
rect 9052 13368 9154 13380
rect 9606 13368 9708 13380
rect 10160 13368 10262 13380
rect 10714 13368 10816 13380
rect 11268 13368 11370 13380
rect 11822 13368 11924 13380
rect 12376 13368 12478 13380
rect 12930 13368 13032 13380
rect 2612 13290 2888 13324
rect 2922 13290 2957 13324
rect 2991 13290 3026 13324
rect 3060 13290 3095 13324
rect 3129 13290 3164 13324
rect 3198 13290 3233 13324
rect 3267 13290 3302 13324
rect 3336 13290 3371 13324
rect 3405 13290 3440 13324
rect 3474 13290 3509 13324
rect 3543 13290 3578 13324
rect 3612 13290 3647 13324
rect 3681 13290 3716 13324
rect 3750 13290 3785 13324
rect 3819 13290 3854 13324
rect 3888 13290 3923 13324
rect 3957 13290 3992 13324
rect 4026 13290 4061 13324
rect 4095 13290 4130 13324
rect 4164 13290 4199 13324
rect 4233 13290 4268 13324
rect 4302 13290 4337 13324
rect 4371 13290 4406 13324
rect 4440 13290 4475 13324
rect 4509 13290 4544 13324
rect 4578 13290 4613 13324
rect 4647 13290 4682 13324
rect 4716 13290 4751 13324
rect 4785 13290 4820 13324
rect 4854 13290 4889 13324
rect 4923 13290 4958 13324
rect 4992 13290 5027 13324
rect 5061 13290 5096 13324
rect 5130 13290 5165 13324
rect 5199 13290 5234 13324
rect 5268 13290 5303 13324
rect 5337 13290 5372 13324
rect 5406 13290 5441 13324
rect 5475 13290 5510 13324
rect 5544 13290 5579 13324
rect 5613 13290 5648 13324
rect 5682 13290 5717 13324
rect 5751 13290 5786 13324
rect 5820 13290 5855 13324
rect 5889 13290 5924 13324
rect 5958 13290 5993 13324
rect 6027 13290 6062 13324
rect 6096 13290 6131 13324
rect 6165 13290 6200 13324
rect 6234 13290 6268 13324
rect 6302 13290 6336 13324
rect 6370 13290 6404 13324
rect 6438 13290 6472 13324
rect 6506 13290 6540 13324
rect 6574 13290 6608 13324
rect 6642 13290 6676 13324
rect 6710 13290 6744 13324
rect 6778 13290 6812 13324
rect 6846 13290 6880 13324
rect 6914 13290 6948 13324
rect 6982 13290 7016 13324
rect 7050 13290 7084 13324
rect 7118 13290 7152 13324
rect 7186 13290 7220 13324
rect 7254 13290 7288 13324
rect 7322 13290 7356 13324
rect 7390 13290 7424 13324
rect 7458 13290 7492 13324
rect 7526 13290 7560 13324
rect 7594 13290 7628 13324
rect 7662 13290 7696 13324
rect 7730 13290 7764 13324
rect 7798 13290 7832 13324
rect 7866 13290 7900 13324
rect 7934 13290 7968 13324
rect 8002 13290 8036 13324
rect 8070 13290 8104 13324
rect 8138 13290 8172 13324
rect 8206 13290 8240 13324
rect 8274 13290 8308 13324
rect 8342 13290 8376 13324
rect 8410 13290 8444 13324
rect 8478 13290 8512 13324
rect 8546 13290 8580 13324
rect 8614 13290 8648 13324
rect 8682 13290 8716 13324
rect 8750 13290 8784 13324
rect 8818 13290 8852 13324
rect 8886 13290 8920 13324
rect 8954 13290 8988 13324
rect 9022 13290 9056 13324
rect 9090 13290 9124 13324
rect 9158 13290 9192 13324
rect 9226 13290 9260 13324
rect 9294 13290 9328 13324
rect 9362 13290 9396 13324
rect 9430 13290 9464 13324
rect 9498 13290 9532 13324
rect 9566 13290 9600 13324
rect 9634 13290 9668 13324
rect 9702 13290 9736 13324
rect 9770 13290 9804 13324
rect 9838 13290 9872 13324
rect 9906 13290 9940 13324
rect 9974 13290 10008 13324
rect 10042 13290 10076 13324
rect 10110 13290 10144 13324
rect 10178 13290 10212 13324
rect 10246 13290 10280 13324
rect 10314 13290 10348 13324
rect 10382 13290 10416 13324
rect 10450 13290 10484 13324
rect 10518 13290 10552 13324
rect 10586 13290 10620 13324
rect 10654 13290 10688 13324
rect 10722 13290 10756 13324
rect 10790 13290 10824 13324
rect 10858 13290 10892 13324
rect 10926 13290 10960 13324
rect 10994 13290 11028 13324
rect 11062 13290 11096 13324
rect 11130 13290 11164 13324
rect 11198 13290 11232 13324
rect 11266 13290 11300 13324
rect 11334 13290 11368 13324
rect 11402 13290 11436 13324
rect 11470 13290 11504 13324
rect 11538 13290 11572 13324
rect 11606 13290 11640 13324
rect 11674 13290 11708 13324
rect 11742 13290 11776 13324
rect 11810 13290 11844 13324
rect 11878 13290 11912 13324
rect 11946 13290 11980 13324
rect 12014 13290 12048 13324
rect 12082 13290 12116 13324
rect 12150 13290 12184 13324
rect 12218 13290 12252 13324
rect 12286 13290 12320 13324
rect 12354 13290 12388 13324
rect 12422 13290 12456 13324
rect 12490 13290 12524 13324
rect 12558 13290 12592 13324
rect 12626 13290 12660 13324
rect 12694 13290 12728 13324
rect 12762 13290 12796 13324
rect 12830 13290 12864 13324
rect 12898 13290 12932 13324
rect 12966 13290 13000 13324
rect 13034 13290 13068 13324
rect 13102 13290 13118 13324
rect 2612 13218 13118 13290
rect 2612 13184 2669 13218
rect 2703 13184 2741 13218
rect 2775 13184 13118 13218
rect 2612 13111 13118 13184
rect 2612 13077 2669 13111
rect 2703 13077 2741 13111
rect 2775 13077 13118 13111
rect 2612 13004 13118 13077
rect 2612 12970 2669 13004
rect 2703 12970 2741 13004
rect 2775 12970 13118 13004
rect 2612 12854 13118 12970
rect 2612 12820 2888 12854
rect 2922 12820 2957 12854
rect 2991 12820 3026 12854
rect 3060 12820 3095 12854
rect 3129 12820 3164 12854
rect 3198 12820 3233 12854
rect 3267 12820 3302 12854
rect 3336 12820 3371 12854
rect 3405 12820 3440 12854
rect 3474 12820 3509 12854
rect 3543 12820 3578 12854
rect 3612 12820 3647 12854
rect 3681 12820 3716 12854
rect 3750 12820 3785 12854
rect 3819 12820 3854 12854
rect 3888 12820 3923 12854
rect 3957 12820 3992 12854
rect 4026 12820 4061 12854
rect 4095 12820 4130 12854
rect 4164 12820 4199 12854
rect 4233 12820 4268 12854
rect 4302 12820 4337 12854
rect 4371 12820 4406 12854
rect 4440 12820 4475 12854
rect 4509 12820 4544 12854
rect 4578 12820 4613 12854
rect 4647 12820 4682 12854
rect 4716 12820 4751 12854
rect 4785 12820 4820 12854
rect 4854 12820 4889 12854
rect 4923 12820 4958 12854
rect 4992 12820 5027 12854
rect 5061 12820 5096 12854
rect 5130 12820 5165 12854
rect 5199 12820 5234 12854
rect 5268 12820 5303 12854
rect 5337 12820 5372 12854
rect 5406 12820 5441 12854
rect 5475 12820 5510 12854
rect 5544 12820 5579 12854
rect 5613 12820 5648 12854
rect 5682 12820 5717 12854
rect 5751 12820 5786 12854
rect 5820 12820 5855 12854
rect 5889 12820 5924 12854
rect 5958 12820 5993 12854
rect 6027 12820 6062 12854
rect 6096 12820 6131 12854
rect 6165 12820 6200 12854
rect 6234 12820 6268 12854
rect 6302 12820 6336 12854
rect 6370 12820 6404 12854
rect 6438 12820 6472 12854
rect 6506 12820 6540 12854
rect 6574 12820 6608 12854
rect 6642 12820 6676 12854
rect 6710 12820 6744 12854
rect 6778 12820 6812 12854
rect 6846 12820 6880 12854
rect 6914 12820 6948 12854
rect 6982 12820 7016 12854
rect 7050 12820 7084 12854
rect 7118 12820 7152 12854
rect 7186 12820 7220 12854
rect 7254 12820 7288 12854
rect 7322 12820 7356 12854
rect 7390 12820 7424 12854
rect 7458 12820 7492 12854
rect 7526 12820 7560 12854
rect 7594 12820 7628 12854
rect 7662 12820 7696 12854
rect 7730 12820 7764 12854
rect 7798 12820 7832 12854
rect 7866 12820 7900 12854
rect 7934 12820 7968 12854
rect 8002 12820 8036 12854
rect 8070 12820 8104 12854
rect 8138 12820 8172 12854
rect 8206 12820 8240 12854
rect 8274 12820 8308 12854
rect 8342 12820 8376 12854
rect 8410 12820 8444 12854
rect 8478 12820 8512 12854
rect 8546 12820 8580 12854
rect 8614 12820 8648 12854
rect 8682 12820 8716 12854
rect 8750 12820 8784 12854
rect 8818 12820 8852 12854
rect 8886 12820 8920 12854
rect 8954 12820 8988 12854
rect 9022 12820 9056 12854
rect 9090 12820 9124 12854
rect 9158 12820 9192 12854
rect 9226 12820 9260 12854
rect 9294 12820 9328 12854
rect 9362 12820 9396 12854
rect 9430 12820 9464 12854
rect 9498 12820 9532 12854
rect 9566 12820 9600 12854
rect 9634 12820 9668 12854
rect 9702 12820 9736 12854
rect 9770 12820 9804 12854
rect 9838 12820 9872 12854
rect 9906 12820 9940 12854
rect 9974 12820 10008 12854
rect 10042 12820 10076 12854
rect 10110 12820 10144 12854
rect 10178 12820 10212 12854
rect 10246 12820 10280 12854
rect 10314 12820 10348 12854
rect 10382 12820 10416 12854
rect 10450 12820 10484 12854
rect 10518 12820 10552 12854
rect 10586 12820 10620 12854
rect 10654 12820 10688 12854
rect 10722 12820 10756 12854
rect 10790 12820 10824 12854
rect 10858 12820 10892 12854
rect 10926 12820 10960 12854
rect 10994 12820 11028 12854
rect 11062 12820 11096 12854
rect 11130 12820 11164 12854
rect 11198 12820 11232 12854
rect 11266 12820 11300 12854
rect 11334 12820 11368 12854
rect 11402 12820 11436 12854
rect 11470 12820 11504 12854
rect 11538 12820 11572 12854
rect 11606 12820 11640 12854
rect 11674 12820 11708 12854
rect 11742 12820 11776 12854
rect 11810 12820 11844 12854
rect 11878 12820 11912 12854
rect 11946 12820 11980 12854
rect 12014 12820 12048 12854
rect 12082 12820 12116 12854
rect 12150 12820 12184 12854
rect 12218 12820 12252 12854
rect 12286 12820 12320 12854
rect 12354 12820 12388 12854
rect 12422 12820 12456 12854
rect 12490 12820 12524 12854
rect 12558 12820 12592 12854
rect 12626 12820 12660 12854
rect 12694 12820 12728 12854
rect 12762 12820 12796 12854
rect 12830 12820 12864 12854
rect 12898 12820 12932 12854
rect 12966 12820 13000 12854
rect 13034 12820 13068 12854
rect 13102 12820 13118 12854
rect 2958 12714 3060 12726
rect 3512 12714 3614 12726
rect 4066 12714 4168 12726
rect 4620 12714 4722 12726
rect 5174 12714 5276 12726
rect 5728 12714 5830 12726
rect 6282 12714 6384 12726
rect 6836 12714 6938 12726
rect 7390 12714 7492 12726
rect 7944 12714 8046 12726
rect 8498 12714 8600 12726
rect 9052 12714 9154 12726
rect 9606 12714 9708 12726
rect 10160 12714 10262 12726
rect 10714 12714 10816 12726
rect 11268 12714 11370 12726
rect 11822 12714 11924 12726
rect 12376 12714 12478 12726
rect 12930 12714 13032 12726
rect 2255 11852 2274 11891
rect 2255 11779 2274 11818
rect 2255 11706 2274 11745
rect 2255 11633 2274 11672
rect 2255 11560 2274 11599
rect 2255 11487 2274 11526
rect 2255 11414 2274 11453
rect 2713 12680 2751 12714
rect 2679 12641 2785 12680
rect 2713 12607 2751 12641
rect 2679 12568 2785 12607
rect 2713 12534 2751 12568
rect 2679 12495 2785 12534
rect 2713 12461 2751 12495
rect 2679 12422 2785 12461
rect 2990 12680 3028 12714
rect 2956 12641 3062 12680
rect 2990 12607 3028 12641
rect 2956 12568 3062 12607
rect 2990 12534 3028 12568
rect 2956 12495 3062 12534
rect 2990 12461 3028 12495
rect 2956 12422 3062 12461
rect 3267 12680 3305 12714
rect 3233 12641 3339 12680
rect 3267 12607 3305 12641
rect 3233 12568 3339 12607
rect 3267 12534 3305 12568
rect 3233 12495 3339 12534
rect 3267 12461 3305 12495
rect 3233 12422 3339 12461
rect 3544 12680 3582 12714
rect 3510 12641 3616 12680
rect 3544 12607 3582 12641
rect 3510 12568 3616 12607
rect 3544 12534 3582 12568
rect 3510 12495 3616 12534
rect 3544 12461 3582 12495
rect 3510 12422 3616 12461
rect 3821 12680 3859 12714
rect 3787 12641 3893 12680
rect 3821 12607 3859 12641
rect 3787 12568 3893 12607
rect 3821 12534 3859 12568
rect 3787 12495 3893 12534
rect 3821 12461 3859 12495
rect 3787 12422 3893 12461
rect 4098 12680 4136 12714
rect 4064 12641 4170 12680
rect 4098 12607 4136 12641
rect 4064 12568 4170 12607
rect 4098 12534 4136 12568
rect 4064 12495 4170 12534
rect 4098 12461 4136 12495
rect 4064 12422 4170 12461
rect 4375 12680 4413 12714
rect 4341 12641 4447 12680
rect 4375 12607 4413 12641
rect 4341 12568 4447 12607
rect 4375 12534 4413 12568
rect 4341 12495 4447 12534
rect 4375 12461 4413 12495
rect 4341 12422 4447 12461
rect 4652 12680 4690 12714
rect 4618 12641 4724 12680
rect 4652 12607 4690 12641
rect 4618 12568 4724 12607
rect 4652 12534 4690 12568
rect 4618 12495 4724 12534
rect 4652 12461 4690 12495
rect 4618 12422 4724 12461
rect 4929 12680 4967 12714
rect 4895 12641 5001 12680
rect 4929 12607 4967 12641
rect 4895 12568 5001 12607
rect 4929 12534 4967 12568
rect 4895 12495 5001 12534
rect 4929 12461 4967 12495
rect 4895 12422 5001 12461
rect 5206 12680 5244 12714
rect 5172 12641 5278 12680
rect 5206 12607 5244 12641
rect 5172 12568 5278 12607
rect 5206 12534 5244 12568
rect 5172 12495 5278 12534
rect 5206 12461 5244 12495
rect 5172 12422 5278 12461
rect 5483 12680 5521 12714
rect 5449 12641 5555 12680
rect 5483 12607 5521 12641
rect 5449 12568 5555 12607
rect 5483 12534 5521 12568
rect 5449 12495 5555 12534
rect 5483 12461 5521 12495
rect 5449 12422 5555 12461
rect 5760 12680 5798 12714
rect 5726 12641 5832 12680
rect 5760 12607 5798 12641
rect 5726 12568 5832 12607
rect 5760 12534 5798 12568
rect 5726 12495 5832 12534
rect 5760 12461 5798 12495
rect 5726 12422 5832 12461
rect 6037 12680 6075 12714
rect 6003 12641 6109 12680
rect 6037 12607 6075 12641
rect 6003 12568 6109 12607
rect 6037 12534 6075 12568
rect 6003 12495 6109 12534
rect 6037 12461 6075 12495
rect 6003 12422 6109 12461
rect 6314 12680 6352 12714
rect 6280 12641 6386 12680
rect 6314 12607 6352 12641
rect 6280 12568 6386 12607
rect 6314 12534 6352 12568
rect 6280 12495 6386 12534
rect 6314 12461 6352 12495
rect 6280 12422 6386 12461
rect 6591 12680 6629 12714
rect 6557 12641 6663 12680
rect 6591 12607 6629 12641
rect 6557 12568 6663 12607
rect 6591 12534 6629 12568
rect 6557 12495 6663 12534
rect 6591 12461 6629 12495
rect 6557 12422 6663 12461
rect 6868 12680 6906 12714
rect 6834 12641 6940 12680
rect 6868 12607 6906 12641
rect 6834 12568 6940 12607
rect 6868 12534 6906 12568
rect 6834 12495 6940 12534
rect 6868 12461 6906 12495
rect 6834 12422 6940 12461
rect 7145 12680 7183 12714
rect 7111 12641 7217 12680
rect 7145 12607 7183 12641
rect 7111 12568 7217 12607
rect 7145 12534 7183 12568
rect 7111 12495 7217 12534
rect 7145 12461 7183 12495
rect 7111 12422 7217 12461
rect 7422 12680 7460 12714
rect 7388 12641 7494 12680
rect 7422 12607 7460 12641
rect 7388 12568 7494 12607
rect 7422 12534 7460 12568
rect 7388 12495 7494 12534
rect 7422 12461 7460 12495
rect 7388 12422 7494 12461
rect 7699 12680 7737 12714
rect 7665 12641 7771 12680
rect 7699 12607 7737 12641
rect 7665 12568 7771 12607
rect 7699 12534 7737 12568
rect 7665 12495 7771 12534
rect 7699 12461 7737 12495
rect 7665 12422 7771 12461
rect 7976 12680 8014 12714
rect 7942 12641 8048 12680
rect 7976 12607 8014 12641
rect 7942 12568 8048 12607
rect 7976 12534 8014 12568
rect 7942 12495 8048 12534
rect 7976 12461 8014 12495
rect 7942 12422 8048 12461
rect 8253 12680 8291 12714
rect 8219 12641 8325 12680
rect 8253 12607 8291 12641
rect 8219 12568 8325 12607
rect 8253 12534 8291 12568
rect 8219 12495 8325 12534
rect 8253 12461 8291 12495
rect 8219 12422 8325 12461
rect 8530 12680 8568 12714
rect 8496 12641 8602 12680
rect 8530 12607 8568 12641
rect 8496 12568 8602 12607
rect 8530 12534 8568 12568
rect 8496 12495 8602 12534
rect 8530 12461 8568 12495
rect 8496 12422 8602 12461
rect 8807 12680 8845 12714
rect 8773 12641 8879 12680
rect 8807 12607 8845 12641
rect 8773 12568 8879 12607
rect 8807 12534 8845 12568
rect 8773 12495 8879 12534
rect 8807 12461 8845 12495
rect 8773 12422 8879 12461
rect 9084 12680 9122 12714
rect 9050 12641 9156 12680
rect 9084 12607 9122 12641
rect 9050 12568 9156 12607
rect 9084 12534 9122 12568
rect 9050 12495 9156 12534
rect 9084 12461 9122 12495
rect 9050 12422 9156 12461
rect 9361 12680 9399 12714
rect 9327 12641 9433 12680
rect 9361 12607 9399 12641
rect 9327 12568 9433 12607
rect 9361 12534 9399 12568
rect 9327 12495 9433 12534
rect 9361 12461 9399 12495
rect 9327 12422 9433 12461
rect 9638 12680 9676 12714
rect 9604 12641 9710 12680
rect 9638 12607 9676 12641
rect 9604 12568 9710 12607
rect 9638 12534 9676 12568
rect 9604 12495 9710 12534
rect 9638 12461 9676 12495
rect 9604 12422 9710 12461
rect 9915 12680 9953 12714
rect 9881 12641 9987 12680
rect 9915 12607 9953 12641
rect 9881 12568 9987 12607
rect 9915 12534 9953 12568
rect 9881 12495 9987 12534
rect 9915 12461 9953 12495
rect 9881 12422 9987 12461
rect 10192 12680 10230 12714
rect 10158 12641 10264 12680
rect 10192 12607 10230 12641
rect 10158 12568 10264 12607
rect 10192 12534 10230 12568
rect 10158 12495 10264 12534
rect 10192 12461 10230 12495
rect 10158 12422 10264 12461
rect 10469 12680 10507 12714
rect 10435 12641 10541 12680
rect 10469 12607 10507 12641
rect 10435 12568 10541 12607
rect 10469 12534 10507 12568
rect 10435 12495 10541 12534
rect 10469 12461 10507 12495
rect 10435 12422 10541 12461
rect 10746 12680 10784 12714
rect 10712 12641 10818 12680
rect 10746 12607 10784 12641
rect 10712 12568 10818 12607
rect 10746 12534 10784 12568
rect 10712 12495 10818 12534
rect 10746 12461 10784 12495
rect 10712 12422 10818 12461
rect 11023 12680 11061 12714
rect 10989 12641 11095 12680
rect 11023 12607 11061 12641
rect 10989 12568 11095 12607
rect 11023 12534 11061 12568
rect 10989 12495 11095 12534
rect 11023 12461 11061 12495
rect 10989 12422 11095 12461
rect 11300 12680 11338 12714
rect 11266 12641 11372 12680
rect 11300 12607 11338 12641
rect 11266 12568 11372 12607
rect 11300 12534 11338 12568
rect 11266 12495 11372 12534
rect 11300 12461 11338 12495
rect 11266 12422 11372 12461
rect 11577 12680 11615 12714
rect 11543 12641 11649 12680
rect 11577 12607 11615 12641
rect 11543 12568 11649 12607
rect 11577 12534 11615 12568
rect 11543 12495 11649 12534
rect 11577 12461 11615 12495
rect 11543 12422 11649 12461
rect 11854 12680 11892 12714
rect 11820 12641 11926 12680
rect 11854 12607 11892 12641
rect 11820 12568 11926 12607
rect 11854 12534 11892 12568
rect 11820 12495 11926 12534
rect 11854 12461 11892 12495
rect 11820 12422 11926 12461
rect 12131 12680 12169 12714
rect 12097 12641 12203 12680
rect 12131 12607 12169 12641
rect 12097 12568 12203 12607
rect 12131 12534 12169 12568
rect 12097 12495 12203 12534
rect 12131 12461 12169 12495
rect 12097 12422 12203 12461
rect 12408 12680 12446 12714
rect 12374 12641 12480 12680
rect 12408 12607 12446 12641
rect 12374 12568 12480 12607
rect 12408 12534 12446 12568
rect 12374 12495 12480 12534
rect 12408 12461 12446 12495
rect 12374 12422 12480 12461
rect 12685 12680 12723 12714
rect 12651 12641 12757 12680
rect 12685 12607 12723 12641
rect 12651 12568 12757 12607
rect 12685 12534 12723 12568
rect 12651 12495 12757 12534
rect 12685 12461 12723 12495
rect 12651 12422 12757 12461
rect 12962 12680 13000 12714
rect 12928 12641 13034 12680
rect 12962 12607 13000 12641
rect 12928 12568 13034 12607
rect 12962 12534 13000 12568
rect 12928 12495 13034 12534
rect 12962 12461 13000 12495
rect 12928 12422 13034 12461
rect 13239 12680 13277 12714
rect 13205 12641 13311 12680
rect 13239 12607 13277 12641
rect 13205 12568 13311 12607
rect 13239 12534 13277 12568
rect 13205 12495 13311 12534
rect 13239 12461 13277 12495
rect 13205 12422 13311 12461
rect 2255 10714 2274 11380
rect 2958 11368 3060 11380
rect 3512 11368 3614 11380
rect 4066 11368 4168 11380
rect 4620 11368 4722 11380
rect 5174 11368 5276 11380
rect 5728 11368 5830 11380
rect 6282 11368 6384 11380
rect 6836 11368 6938 11380
rect 7390 11368 7492 11380
rect 7944 11368 8046 11380
rect 8498 11368 8600 11380
rect 9052 11368 9154 11380
rect 9606 11368 9708 11380
rect 10160 11368 10262 11380
rect 10714 11368 10816 11380
rect 11268 11368 11370 11380
rect 11822 11368 11924 11380
rect 12376 11368 12478 11380
rect 12930 11368 13032 11380
rect 2638 11290 2888 11324
rect 2922 11290 2957 11324
rect 2991 11290 3026 11324
rect 3060 11290 3095 11324
rect 3129 11290 3164 11324
rect 3198 11290 3233 11324
rect 3267 11290 3302 11324
rect 3336 11290 3371 11324
rect 3405 11290 3440 11324
rect 3474 11290 3509 11324
rect 3543 11290 3578 11324
rect 3612 11290 3647 11324
rect 3681 11290 3716 11324
rect 3750 11290 3785 11324
rect 3819 11290 3854 11324
rect 3888 11290 3923 11324
rect 3957 11290 3992 11324
rect 4026 11290 4061 11324
rect 4095 11290 4130 11324
rect 4164 11290 4199 11324
rect 4233 11290 4268 11324
rect 4302 11290 4337 11324
rect 4371 11290 4406 11324
rect 4440 11290 4475 11324
rect 4509 11290 4544 11324
rect 4578 11290 4613 11324
rect 4647 11290 4682 11324
rect 4716 11290 4751 11324
rect 4785 11290 4820 11324
rect 4854 11290 4889 11324
rect 4923 11290 4958 11324
rect 4992 11290 5027 11324
rect 5061 11290 5096 11324
rect 5130 11290 5165 11324
rect 5199 11290 5234 11324
rect 5268 11290 5303 11324
rect 5337 11290 5372 11324
rect 5406 11290 5441 11324
rect 5475 11290 5510 11324
rect 5544 11290 5579 11324
rect 5613 11290 5648 11324
rect 5682 11290 5717 11324
rect 5751 11290 5786 11324
rect 5820 11290 5855 11324
rect 5889 11290 5924 11324
rect 5958 11290 5993 11324
rect 6027 11290 6062 11324
rect 6096 11290 6131 11324
rect 6165 11290 6200 11324
rect 6234 11290 6268 11324
rect 6302 11290 6336 11324
rect 6370 11290 6404 11324
rect 6438 11290 6472 11324
rect 6506 11290 6540 11324
rect 6574 11290 6608 11324
rect 6642 11290 6676 11324
rect 6710 11290 6744 11324
rect 6778 11290 6812 11324
rect 6846 11290 6880 11324
rect 6914 11290 6948 11324
rect 6982 11290 7016 11324
rect 7050 11290 7084 11324
rect 7118 11290 7152 11324
rect 7186 11290 7220 11324
rect 7254 11290 7288 11324
rect 7322 11290 7356 11324
rect 7390 11290 7424 11324
rect 7458 11290 7492 11324
rect 7526 11290 7560 11324
rect 7594 11290 7628 11324
rect 7662 11290 7696 11324
rect 7730 11290 7764 11324
rect 7798 11290 7832 11324
rect 7866 11290 7900 11324
rect 7934 11290 7968 11324
rect 8002 11290 8036 11324
rect 8070 11290 8104 11324
rect 8138 11290 8172 11324
rect 8206 11290 8240 11324
rect 8274 11290 8308 11324
rect 8342 11290 8376 11324
rect 8410 11290 8444 11324
rect 8478 11290 8512 11324
rect 8546 11290 8580 11324
rect 8614 11290 8648 11324
rect 8682 11290 8716 11324
rect 8750 11290 8784 11324
rect 8818 11290 8852 11324
rect 8886 11290 8920 11324
rect 8954 11290 8988 11324
rect 9022 11290 9056 11324
rect 9090 11290 9124 11324
rect 9158 11290 9192 11324
rect 9226 11290 9260 11324
rect 9294 11290 9328 11324
rect 9362 11290 9396 11324
rect 9430 11290 9464 11324
rect 9498 11290 9532 11324
rect 9566 11290 9600 11324
rect 9634 11290 9668 11324
rect 9702 11290 9736 11324
rect 9770 11290 9804 11324
rect 9838 11290 9872 11324
rect 9906 11290 9940 11324
rect 9974 11290 10008 11324
rect 10042 11290 10076 11324
rect 10110 11290 10144 11324
rect 10178 11290 10212 11324
rect 10246 11290 10280 11324
rect 10314 11290 10348 11324
rect 10382 11290 10416 11324
rect 10450 11290 10484 11324
rect 10518 11290 10552 11324
rect 10586 11290 10620 11324
rect 10654 11290 10688 11324
rect 10722 11290 10756 11324
rect 10790 11290 10824 11324
rect 10858 11290 10892 11324
rect 10926 11290 10960 11324
rect 10994 11290 11028 11324
rect 11062 11290 11096 11324
rect 11130 11290 11164 11324
rect 11198 11290 11232 11324
rect 11266 11290 11300 11324
rect 11334 11290 11368 11324
rect 11402 11290 11436 11324
rect 11470 11290 11504 11324
rect 11538 11290 11572 11324
rect 11606 11290 11640 11324
rect 11674 11290 11708 11324
rect 11742 11290 11776 11324
rect 11810 11290 11844 11324
rect 11878 11290 11912 11324
rect 11946 11290 11980 11324
rect 12014 11290 12048 11324
rect 12082 11290 12116 11324
rect 12150 11290 12184 11324
rect 12218 11290 12252 11324
rect 12286 11290 12320 11324
rect 12354 11290 12388 11324
rect 12422 11290 12456 11324
rect 12490 11290 12524 11324
rect 12558 11290 12592 11324
rect 12626 11290 12660 11324
rect 12694 11290 12728 11324
rect 12762 11290 12796 11324
rect 12830 11290 12864 11324
rect 12898 11290 12932 11324
rect 12966 11290 13000 11324
rect 13034 11290 13068 11324
rect 13102 11290 13118 11324
rect 2638 11194 13118 11290
rect 2672 11160 2710 11194
rect 2744 11160 13118 11194
rect 2638 11087 13118 11160
rect 2672 11053 2710 11087
rect 2744 11053 13118 11087
rect 2638 10980 13118 11053
rect 2672 10946 2710 10980
rect 2744 10946 13118 10980
rect 2638 10854 13118 10946
rect 2638 10820 2888 10854
rect 2922 10820 2957 10854
rect 2991 10820 3026 10854
rect 3060 10820 3095 10854
rect 3129 10820 3164 10854
rect 3198 10820 3233 10854
rect 3267 10820 3302 10854
rect 3336 10820 3371 10854
rect 3405 10820 3440 10854
rect 3474 10820 3509 10854
rect 3543 10820 3578 10854
rect 3612 10820 3647 10854
rect 3681 10820 3716 10854
rect 3750 10820 3785 10854
rect 3819 10820 3854 10854
rect 3888 10820 3923 10854
rect 3957 10820 3992 10854
rect 4026 10820 4061 10854
rect 4095 10820 4130 10854
rect 4164 10820 4199 10854
rect 4233 10820 4268 10854
rect 4302 10820 4337 10854
rect 4371 10820 4406 10854
rect 4440 10820 4475 10854
rect 4509 10820 4544 10854
rect 4578 10820 4613 10854
rect 4647 10820 4682 10854
rect 4716 10820 4751 10854
rect 4785 10820 4820 10854
rect 4854 10820 4889 10854
rect 4923 10820 4958 10854
rect 4992 10820 5027 10854
rect 5061 10820 5096 10854
rect 5130 10820 5165 10854
rect 5199 10820 5234 10854
rect 5268 10820 5303 10854
rect 5337 10820 5372 10854
rect 5406 10820 5441 10854
rect 5475 10820 5510 10854
rect 5544 10820 5579 10854
rect 5613 10820 5648 10854
rect 5682 10820 5717 10854
rect 5751 10820 5786 10854
rect 5820 10820 5855 10854
rect 5889 10820 5924 10854
rect 5958 10820 5993 10854
rect 6027 10820 6062 10854
rect 6096 10820 6131 10854
rect 6165 10820 6200 10854
rect 6234 10820 6268 10854
rect 6302 10820 6336 10854
rect 6370 10820 6404 10854
rect 6438 10820 6472 10854
rect 6506 10820 6540 10854
rect 6574 10820 6608 10854
rect 6642 10820 6676 10854
rect 6710 10820 6744 10854
rect 6778 10820 6812 10854
rect 6846 10820 6880 10854
rect 6914 10820 6948 10854
rect 6982 10820 7016 10854
rect 7050 10820 7084 10854
rect 7118 10820 7152 10854
rect 7186 10820 7220 10854
rect 7254 10820 7288 10854
rect 7322 10820 7356 10854
rect 7390 10820 7424 10854
rect 7458 10820 7492 10854
rect 7526 10820 7560 10854
rect 7594 10820 7628 10854
rect 7662 10820 7696 10854
rect 7730 10820 7764 10854
rect 7798 10820 7832 10854
rect 7866 10820 7900 10854
rect 7934 10820 7968 10854
rect 8002 10820 8036 10854
rect 8070 10820 8104 10854
rect 8138 10820 8172 10854
rect 8206 10820 8240 10854
rect 8274 10820 8308 10854
rect 8342 10820 8376 10854
rect 8410 10820 8444 10854
rect 8478 10820 8512 10854
rect 8546 10820 8580 10854
rect 8614 10820 8648 10854
rect 8682 10820 8716 10854
rect 8750 10820 8784 10854
rect 8818 10820 8852 10854
rect 8886 10820 8920 10854
rect 8954 10820 8988 10854
rect 9022 10820 9056 10854
rect 9090 10820 9124 10854
rect 9158 10820 9192 10854
rect 9226 10820 9260 10854
rect 9294 10820 9328 10854
rect 9362 10820 9396 10854
rect 9430 10820 9464 10854
rect 9498 10820 9532 10854
rect 9566 10820 9600 10854
rect 9634 10820 9668 10854
rect 9702 10820 9736 10854
rect 9770 10820 9804 10854
rect 9838 10820 9872 10854
rect 9906 10820 9940 10854
rect 9974 10820 10008 10854
rect 10042 10820 10076 10854
rect 10110 10820 10144 10854
rect 10178 10820 10212 10854
rect 10246 10820 10280 10854
rect 10314 10820 10348 10854
rect 10382 10820 10416 10854
rect 10450 10820 10484 10854
rect 10518 10820 10552 10854
rect 10586 10820 10620 10854
rect 10654 10820 10688 10854
rect 10722 10820 10756 10854
rect 10790 10820 10824 10854
rect 10858 10820 10892 10854
rect 10926 10820 10960 10854
rect 10994 10820 11028 10854
rect 11062 10820 11096 10854
rect 11130 10820 11164 10854
rect 11198 10820 11232 10854
rect 11266 10820 11300 10854
rect 11334 10820 11368 10854
rect 11402 10820 11436 10854
rect 11470 10820 11504 10854
rect 11538 10820 11572 10854
rect 11606 10820 11640 10854
rect 11674 10820 11708 10854
rect 11742 10820 11776 10854
rect 11810 10820 11844 10854
rect 11878 10820 11912 10854
rect 11946 10820 11980 10854
rect 12014 10820 12048 10854
rect 12082 10820 12116 10854
rect 12150 10820 12184 10854
rect 12218 10820 12252 10854
rect 12286 10820 12320 10854
rect 12354 10820 12388 10854
rect 12422 10820 12456 10854
rect 12490 10820 12524 10854
rect 12558 10820 12592 10854
rect 12626 10820 12660 10854
rect 12694 10820 12728 10854
rect 12762 10820 12796 10854
rect 12830 10820 12864 10854
rect 12898 10820 12932 10854
rect 12966 10820 13000 10854
rect 13034 10820 13068 10854
rect 13102 10820 13118 10854
rect 2958 10714 3060 10726
rect 3512 10714 3614 10726
rect 4066 10714 4168 10726
rect 4620 10714 4722 10726
rect 5174 10714 5276 10726
rect 5728 10714 5830 10726
rect 6282 10714 6384 10726
rect 6836 10714 6938 10726
rect 7390 10714 7492 10726
rect 7944 10714 8046 10726
rect 8498 10714 8600 10726
rect 9052 10714 9154 10726
rect 9606 10714 9708 10726
rect 10160 10714 10262 10726
rect 10714 10714 10816 10726
rect 11268 10714 11370 10726
rect 11822 10714 11924 10726
rect 12376 10714 12478 10726
rect 12930 10714 13032 10726
rect 2255 9561 2274 9600
rect 2255 9488 2274 9527
rect 2255 9415 2274 9454
rect 1837 7618 1944 8732
rect 2050 7618 2056 8732
rect 2713 10680 2751 10714
rect 2679 10641 2785 10680
rect 2713 10607 2751 10641
rect 2679 10568 2785 10607
rect 2713 10534 2751 10568
rect 2679 10495 2785 10534
rect 2713 10461 2751 10495
rect 2679 10422 2785 10461
rect 2990 10680 3028 10714
rect 2956 10641 3062 10680
rect 2990 10607 3028 10641
rect 2956 10568 3062 10607
rect 2990 10534 3028 10568
rect 2956 10495 3062 10534
rect 2990 10461 3028 10495
rect 2956 10422 3062 10461
rect 3267 10680 3305 10714
rect 3233 10641 3339 10680
rect 3267 10607 3305 10641
rect 3233 10568 3339 10607
rect 3267 10534 3305 10568
rect 3233 10495 3339 10534
rect 3267 10461 3305 10495
rect 3233 10422 3339 10461
rect 3544 10680 3582 10714
rect 3510 10641 3616 10680
rect 3544 10607 3582 10641
rect 3510 10568 3616 10607
rect 3544 10534 3582 10568
rect 3510 10495 3616 10534
rect 3544 10461 3582 10495
rect 3510 10422 3616 10461
rect 3821 10680 3859 10714
rect 3787 10641 3893 10680
rect 3821 10607 3859 10641
rect 3787 10568 3893 10607
rect 3821 10534 3859 10568
rect 3787 10495 3893 10534
rect 3821 10461 3859 10495
rect 3787 10422 3893 10461
rect 4098 10680 4136 10714
rect 4064 10641 4170 10680
rect 4098 10607 4136 10641
rect 4064 10568 4170 10607
rect 4098 10534 4136 10568
rect 4064 10495 4170 10534
rect 4098 10461 4136 10495
rect 4064 10422 4170 10461
rect 4375 10680 4413 10714
rect 4341 10641 4447 10680
rect 4375 10607 4413 10641
rect 4341 10568 4447 10607
rect 4375 10534 4413 10568
rect 4341 10495 4447 10534
rect 4375 10461 4413 10495
rect 4341 10422 4447 10461
rect 4652 10680 4690 10714
rect 4618 10641 4724 10680
rect 4652 10607 4690 10641
rect 4618 10568 4724 10607
rect 4652 10534 4690 10568
rect 4618 10495 4724 10534
rect 4652 10461 4690 10495
rect 4618 10422 4724 10461
rect 4929 10680 4967 10714
rect 4895 10641 5001 10680
rect 4929 10607 4967 10641
rect 4895 10568 5001 10607
rect 4929 10534 4967 10568
rect 4895 10495 5001 10534
rect 4929 10461 4967 10495
rect 4895 10422 5001 10461
rect 5206 10680 5244 10714
rect 5172 10641 5278 10680
rect 5206 10607 5244 10641
rect 5172 10568 5278 10607
rect 5206 10534 5244 10568
rect 5172 10495 5278 10534
rect 5206 10461 5244 10495
rect 5172 10422 5278 10461
rect 5483 10680 5521 10714
rect 5449 10641 5555 10680
rect 5483 10607 5521 10641
rect 5449 10568 5555 10607
rect 5483 10534 5521 10568
rect 5449 10495 5555 10534
rect 5483 10461 5521 10495
rect 5449 10422 5555 10461
rect 5760 10680 5798 10714
rect 5726 10641 5832 10680
rect 5760 10607 5798 10641
rect 5726 10568 5832 10607
rect 5760 10534 5798 10568
rect 5726 10495 5832 10534
rect 5760 10461 5798 10495
rect 5726 10422 5832 10461
rect 6037 10680 6075 10714
rect 6003 10641 6109 10680
rect 6037 10607 6075 10641
rect 6003 10568 6109 10607
rect 6037 10534 6075 10568
rect 6003 10495 6109 10534
rect 6037 10461 6075 10495
rect 6003 10422 6109 10461
rect 6314 10680 6352 10714
rect 6280 10641 6386 10680
rect 6314 10607 6352 10641
rect 6280 10568 6386 10607
rect 6314 10534 6352 10568
rect 6280 10495 6386 10534
rect 6314 10461 6352 10495
rect 6280 10422 6386 10461
rect 6591 10680 6629 10714
rect 6557 10641 6663 10680
rect 6591 10607 6629 10641
rect 6557 10568 6663 10607
rect 6591 10534 6629 10568
rect 6557 10495 6663 10534
rect 6591 10461 6629 10495
rect 6557 10422 6663 10461
rect 6868 10680 6906 10714
rect 6834 10641 6940 10680
rect 6868 10607 6906 10641
rect 6834 10568 6940 10607
rect 6868 10534 6906 10568
rect 6834 10495 6940 10534
rect 6868 10461 6906 10495
rect 6834 10422 6940 10461
rect 7145 10680 7183 10714
rect 7111 10641 7217 10680
rect 7145 10607 7183 10641
rect 7111 10568 7217 10607
rect 7145 10534 7183 10568
rect 7111 10495 7217 10534
rect 7145 10461 7183 10495
rect 7111 10422 7217 10461
rect 7422 10680 7460 10714
rect 7388 10641 7494 10680
rect 7422 10607 7460 10641
rect 7388 10568 7494 10607
rect 7422 10534 7460 10568
rect 7388 10495 7494 10534
rect 7422 10461 7460 10495
rect 7388 10422 7494 10461
rect 7699 10680 7737 10714
rect 7665 10641 7771 10680
rect 7699 10607 7737 10641
rect 7665 10568 7771 10607
rect 7699 10534 7737 10568
rect 7665 10495 7771 10534
rect 7699 10461 7737 10495
rect 7665 10422 7771 10461
rect 7976 10680 8014 10714
rect 7942 10641 8048 10680
rect 7976 10607 8014 10641
rect 7942 10568 8048 10607
rect 7976 10534 8014 10568
rect 7942 10495 8048 10534
rect 7976 10461 8014 10495
rect 7942 10422 8048 10461
rect 8253 10680 8291 10714
rect 8219 10641 8325 10680
rect 8253 10607 8291 10641
rect 8219 10568 8325 10607
rect 8253 10534 8291 10568
rect 8219 10495 8325 10534
rect 8253 10461 8291 10495
rect 8219 10422 8325 10461
rect 8530 10680 8568 10714
rect 8496 10641 8602 10680
rect 8530 10607 8568 10641
rect 8496 10568 8602 10607
rect 8530 10534 8568 10568
rect 8496 10495 8602 10534
rect 8530 10461 8568 10495
rect 8496 10422 8602 10461
rect 8807 10680 8845 10714
rect 8773 10641 8879 10680
rect 8807 10607 8845 10641
rect 8773 10568 8879 10607
rect 8807 10534 8845 10568
rect 8773 10495 8879 10534
rect 8807 10461 8845 10495
rect 8773 10422 8879 10461
rect 9084 10680 9122 10714
rect 9050 10641 9156 10680
rect 9084 10607 9122 10641
rect 9050 10568 9156 10607
rect 9084 10534 9122 10568
rect 9050 10495 9156 10534
rect 9084 10461 9122 10495
rect 9050 10422 9156 10461
rect 9361 10680 9399 10714
rect 9327 10641 9433 10680
rect 9361 10607 9399 10641
rect 9327 10568 9433 10607
rect 9361 10534 9399 10568
rect 9327 10495 9433 10534
rect 9361 10461 9399 10495
rect 9327 10422 9433 10461
rect 9638 10680 9676 10714
rect 9604 10641 9710 10680
rect 9638 10607 9676 10641
rect 9604 10568 9710 10607
rect 9638 10534 9676 10568
rect 9604 10495 9710 10534
rect 9638 10461 9676 10495
rect 9604 10422 9710 10461
rect 9915 10680 9953 10714
rect 9881 10641 9987 10680
rect 9915 10607 9953 10641
rect 9881 10568 9987 10607
rect 9915 10534 9953 10568
rect 9881 10495 9987 10534
rect 9915 10461 9953 10495
rect 9881 10422 9987 10461
rect 10192 10680 10230 10714
rect 10158 10641 10264 10680
rect 10192 10607 10230 10641
rect 10158 10568 10264 10607
rect 10192 10534 10230 10568
rect 10158 10495 10264 10534
rect 10192 10461 10230 10495
rect 10158 10422 10264 10461
rect 10469 10680 10507 10714
rect 10435 10641 10541 10680
rect 10469 10607 10507 10641
rect 10435 10568 10541 10607
rect 10469 10534 10507 10568
rect 10435 10495 10541 10534
rect 10469 10461 10507 10495
rect 10435 10422 10541 10461
rect 10746 10680 10784 10714
rect 10712 10641 10818 10680
rect 10746 10607 10784 10641
rect 10712 10568 10818 10607
rect 10746 10534 10784 10568
rect 10712 10495 10818 10534
rect 10746 10461 10784 10495
rect 10712 10422 10818 10461
rect 11023 10680 11061 10714
rect 10989 10641 11095 10680
rect 11023 10607 11061 10641
rect 10989 10568 11095 10607
rect 11023 10534 11061 10568
rect 10989 10495 11095 10534
rect 11023 10461 11061 10495
rect 10989 10422 11095 10461
rect 11300 10680 11338 10714
rect 11266 10641 11372 10680
rect 11300 10607 11338 10641
rect 11266 10568 11372 10607
rect 11300 10534 11338 10568
rect 11266 10495 11372 10534
rect 11300 10461 11338 10495
rect 11266 10422 11372 10461
rect 11577 10680 11615 10714
rect 11543 10641 11649 10680
rect 11577 10607 11615 10641
rect 11543 10568 11649 10607
rect 11577 10534 11615 10568
rect 11543 10495 11649 10534
rect 11577 10461 11615 10495
rect 11543 10422 11649 10461
rect 11854 10680 11892 10714
rect 11820 10641 11926 10680
rect 11854 10607 11892 10641
rect 11820 10568 11926 10607
rect 11854 10534 11892 10568
rect 11820 10495 11926 10534
rect 11854 10461 11892 10495
rect 11820 10422 11926 10461
rect 12131 10680 12169 10714
rect 12097 10641 12203 10680
rect 12131 10607 12169 10641
rect 12097 10568 12203 10607
rect 12131 10534 12169 10568
rect 12097 10495 12203 10534
rect 12131 10461 12169 10495
rect 12097 10422 12203 10461
rect 12408 10680 12446 10714
rect 12374 10641 12480 10680
rect 12408 10607 12446 10641
rect 12374 10568 12480 10607
rect 12408 10534 12446 10568
rect 12374 10495 12480 10534
rect 12408 10461 12446 10495
rect 12374 10422 12480 10461
rect 12685 10680 12723 10714
rect 12651 10641 12757 10680
rect 12685 10607 12723 10641
rect 12651 10568 12757 10607
rect 12685 10534 12723 10568
rect 12651 10495 12757 10534
rect 12685 10461 12723 10495
rect 12651 10422 12757 10461
rect 12962 10680 13000 10714
rect 12928 10641 13034 10680
rect 12962 10607 13000 10641
rect 12928 10568 13034 10607
rect 12962 10534 13000 10568
rect 12928 10495 13034 10534
rect 12962 10461 13000 10495
rect 12928 10422 13034 10461
rect 13239 10680 13277 10714
rect 13205 10641 13311 10680
rect 13239 10607 13277 10641
rect 13205 10568 13311 10607
rect 13239 10534 13277 10568
rect 13205 10495 13311 10534
rect 13239 10461 13277 10495
rect 13205 10422 13311 10461
rect 2958 9368 3060 9380
rect 3512 9368 3614 9380
rect 4066 9368 4168 9380
rect 4620 9368 4722 9380
rect 5174 9368 5276 9380
rect 5728 9368 5830 9380
rect 6282 9368 6384 9380
rect 6836 9368 6938 9380
rect 7390 9368 7492 9380
rect 7944 9368 8046 9380
rect 8498 9368 8600 9380
rect 9052 9368 9154 9380
rect 9606 9368 9708 9380
rect 10160 9368 10262 9380
rect 10714 9368 10816 9380
rect 11268 9368 11370 9380
rect 11822 9368 11924 9380
rect 12376 9368 12478 9380
rect 12930 9368 13032 9380
rect 2612 9290 2888 9324
rect 2922 9290 2957 9324
rect 2991 9290 3026 9324
rect 3060 9290 3095 9324
rect 3129 9290 3164 9324
rect 3198 9290 3233 9324
rect 3267 9290 3302 9324
rect 3336 9290 3371 9324
rect 3405 9290 3440 9324
rect 3474 9290 3509 9324
rect 3543 9290 3578 9324
rect 3612 9290 3647 9324
rect 3681 9290 3716 9324
rect 3750 9290 3785 9324
rect 3819 9290 3854 9324
rect 3888 9290 3923 9324
rect 3957 9290 3992 9324
rect 4026 9290 4061 9324
rect 4095 9290 4130 9324
rect 4164 9290 4199 9324
rect 4233 9290 4268 9324
rect 4302 9290 4337 9324
rect 4371 9290 4406 9324
rect 4440 9290 4475 9324
rect 4509 9290 4544 9324
rect 4578 9290 4613 9324
rect 4647 9290 4682 9324
rect 4716 9290 4751 9324
rect 4785 9290 4820 9324
rect 4854 9290 4889 9324
rect 4923 9290 4958 9324
rect 4992 9290 5027 9324
rect 5061 9290 5096 9324
rect 5130 9290 5165 9324
rect 5199 9290 5234 9324
rect 5268 9290 5303 9324
rect 5337 9290 5372 9324
rect 5406 9290 5441 9324
rect 5475 9290 5510 9324
rect 5544 9290 5579 9324
rect 5613 9290 5648 9324
rect 5682 9290 5717 9324
rect 5751 9290 5786 9324
rect 5820 9290 5855 9324
rect 5889 9290 5924 9324
rect 5958 9290 5993 9324
rect 6027 9290 6062 9324
rect 6096 9290 6131 9324
rect 6165 9290 6200 9324
rect 6234 9290 6268 9324
rect 6302 9290 6336 9324
rect 6370 9290 6404 9324
rect 6438 9290 6472 9324
rect 6506 9290 6540 9324
rect 6574 9290 6608 9324
rect 6642 9290 6676 9324
rect 6710 9290 6744 9324
rect 6778 9290 6812 9324
rect 6846 9290 6880 9324
rect 6914 9290 6948 9324
rect 6982 9290 7016 9324
rect 7050 9290 7084 9324
rect 7118 9290 7152 9324
rect 7186 9290 7220 9324
rect 7254 9290 7288 9324
rect 7322 9290 7356 9324
rect 7390 9290 7424 9324
rect 7458 9290 7492 9324
rect 7526 9290 7560 9324
rect 7594 9290 7628 9324
rect 7662 9290 7696 9324
rect 7730 9290 7764 9324
rect 7798 9290 7832 9324
rect 7866 9290 7900 9324
rect 7934 9290 7968 9324
rect 8002 9290 8036 9324
rect 8070 9290 8104 9324
rect 8138 9290 8172 9324
rect 8206 9290 8240 9324
rect 8274 9290 8308 9324
rect 8342 9290 8376 9324
rect 8410 9290 8444 9324
rect 8478 9290 8512 9324
rect 8546 9290 8580 9324
rect 8614 9290 8648 9324
rect 8682 9290 8716 9324
rect 8750 9290 8784 9324
rect 8818 9290 8852 9324
rect 8886 9290 8920 9324
rect 8954 9290 8988 9324
rect 9022 9290 9056 9324
rect 9090 9290 9124 9324
rect 9158 9290 9192 9324
rect 9226 9290 9260 9324
rect 9294 9290 9328 9324
rect 9362 9290 9396 9324
rect 9430 9290 9464 9324
rect 9498 9290 9532 9324
rect 9566 9290 9600 9324
rect 9634 9290 9668 9324
rect 9702 9290 9736 9324
rect 9770 9290 9804 9324
rect 9838 9290 9872 9324
rect 9906 9290 9940 9324
rect 9974 9290 10008 9324
rect 10042 9290 10076 9324
rect 10110 9290 10144 9324
rect 10178 9290 10212 9324
rect 10246 9290 10280 9324
rect 10314 9290 10348 9324
rect 10382 9290 10416 9324
rect 10450 9290 10484 9324
rect 10518 9290 10552 9324
rect 10586 9290 10620 9324
rect 10654 9290 10688 9324
rect 10722 9290 10756 9324
rect 10790 9290 10824 9324
rect 10858 9290 10892 9324
rect 10926 9290 10960 9324
rect 10994 9290 11028 9324
rect 11062 9290 11096 9324
rect 11130 9290 11164 9324
rect 11198 9290 11232 9324
rect 11266 9290 11300 9324
rect 11334 9290 11368 9324
rect 11402 9290 11436 9324
rect 11470 9290 11504 9324
rect 11538 9290 11572 9324
rect 11606 9290 11640 9324
rect 11674 9290 11708 9324
rect 11742 9290 11776 9324
rect 11810 9290 11844 9324
rect 11878 9290 11912 9324
rect 11946 9290 11980 9324
rect 12014 9290 12048 9324
rect 12082 9290 12116 9324
rect 12150 9290 12184 9324
rect 12218 9290 12252 9324
rect 12286 9290 12320 9324
rect 12354 9290 12388 9324
rect 12422 9290 12456 9324
rect 12490 9290 12524 9324
rect 12558 9290 12592 9324
rect 12626 9290 12660 9324
rect 12694 9290 12728 9324
rect 12762 9290 12796 9324
rect 12830 9290 12864 9324
rect 12898 9290 12932 9324
rect 12966 9290 13000 9324
rect 13034 9290 13068 9324
rect 13102 9290 13118 9324
rect 2612 9233 13118 9290
rect 2646 9199 2684 9233
rect 2718 9199 13118 9233
rect 2612 9160 13118 9199
rect 2646 9126 2684 9160
rect 2718 9126 13118 9160
rect 2612 9086 13118 9126
rect 2646 9052 2684 9086
rect 2718 9052 13118 9086
rect 2612 9012 13118 9052
rect 2646 8978 2684 9012
rect 2718 8978 13118 9012
rect 2612 8938 13118 8978
rect 2646 8904 2684 8938
rect 2718 8904 13118 8938
rect 2612 8854 13118 8904
rect 2612 8820 2888 8854
rect 2922 8820 2957 8854
rect 2991 8820 3026 8854
rect 3060 8820 3095 8854
rect 3129 8820 3164 8854
rect 3198 8820 3233 8854
rect 3267 8820 3302 8854
rect 3336 8820 3371 8854
rect 3405 8820 3440 8854
rect 3474 8820 3509 8854
rect 3543 8820 3578 8854
rect 3612 8820 3647 8854
rect 3681 8820 3716 8854
rect 3750 8820 3785 8854
rect 3819 8820 3854 8854
rect 3888 8820 3923 8854
rect 3957 8820 3992 8854
rect 4026 8820 4061 8854
rect 4095 8820 4130 8854
rect 4164 8820 4199 8854
rect 4233 8820 4268 8854
rect 4302 8820 4337 8854
rect 4371 8820 4406 8854
rect 4440 8820 4475 8854
rect 4509 8820 4544 8854
rect 4578 8820 4613 8854
rect 4647 8820 4682 8854
rect 4716 8820 4751 8854
rect 4785 8820 4820 8854
rect 4854 8820 4889 8854
rect 4923 8820 4958 8854
rect 4992 8820 5027 8854
rect 5061 8820 5096 8854
rect 5130 8820 5165 8854
rect 5199 8820 5234 8854
rect 5268 8820 5303 8854
rect 5337 8820 5372 8854
rect 5406 8820 5441 8854
rect 5475 8820 5510 8854
rect 5544 8820 5579 8854
rect 5613 8820 5648 8854
rect 5682 8820 5717 8854
rect 5751 8820 5786 8854
rect 5820 8820 5855 8854
rect 5889 8820 5924 8854
rect 5958 8820 5993 8854
rect 6027 8820 6062 8854
rect 6096 8820 6131 8854
rect 6165 8820 6200 8854
rect 6234 8820 6268 8854
rect 6302 8820 6336 8854
rect 6370 8820 6404 8854
rect 6438 8820 6472 8854
rect 6506 8820 6540 8854
rect 6574 8820 6608 8854
rect 6642 8820 6676 8854
rect 6710 8820 6744 8854
rect 6778 8820 6812 8854
rect 6846 8820 6880 8854
rect 6914 8820 6948 8854
rect 6982 8820 7016 8854
rect 7050 8820 7084 8854
rect 7118 8820 7152 8854
rect 7186 8820 7220 8854
rect 7254 8820 7288 8854
rect 7322 8820 7356 8854
rect 7390 8820 7424 8854
rect 7458 8820 7492 8854
rect 7526 8820 7560 8854
rect 7594 8820 7628 8854
rect 7662 8820 7696 8854
rect 7730 8820 7764 8854
rect 7798 8820 7832 8854
rect 7866 8820 7900 8854
rect 7934 8820 7968 8854
rect 8002 8820 8036 8854
rect 8070 8820 8104 8854
rect 8138 8820 8172 8854
rect 8206 8820 8240 8854
rect 8274 8820 8308 8854
rect 8342 8820 8376 8854
rect 8410 8820 8444 8854
rect 8478 8820 8512 8854
rect 8546 8820 8580 8854
rect 8614 8820 8648 8854
rect 8682 8820 8716 8854
rect 8750 8820 8784 8854
rect 8818 8820 8852 8854
rect 8886 8820 8920 8854
rect 8954 8820 8988 8854
rect 9022 8820 9056 8854
rect 9090 8820 9124 8854
rect 9158 8820 9192 8854
rect 9226 8820 9260 8854
rect 9294 8820 9328 8854
rect 9362 8820 9396 8854
rect 9430 8820 9464 8854
rect 9498 8820 9532 8854
rect 9566 8820 9600 8854
rect 9634 8820 9668 8854
rect 9702 8820 9736 8854
rect 9770 8820 9804 8854
rect 9838 8820 9872 8854
rect 9906 8820 9940 8854
rect 9974 8820 10008 8854
rect 10042 8820 10076 8854
rect 10110 8820 10144 8854
rect 10178 8820 10212 8854
rect 10246 8820 10280 8854
rect 10314 8820 10348 8854
rect 10382 8820 10416 8854
rect 10450 8820 10484 8854
rect 10518 8820 10552 8854
rect 10586 8820 10620 8854
rect 10654 8820 10688 8854
rect 10722 8820 10756 8854
rect 10790 8820 10824 8854
rect 10858 8820 10892 8854
rect 10926 8820 10960 8854
rect 10994 8820 11028 8854
rect 11062 8820 11096 8854
rect 11130 8820 11164 8854
rect 11198 8820 11232 8854
rect 11266 8820 11300 8854
rect 11334 8820 11368 8854
rect 11402 8820 11436 8854
rect 11470 8820 11504 8854
rect 11538 8820 11572 8854
rect 11606 8820 11640 8854
rect 11674 8820 11708 8854
rect 11742 8820 11776 8854
rect 11810 8820 11844 8854
rect 11878 8820 11912 8854
rect 11946 8820 11980 8854
rect 12014 8820 12048 8854
rect 12082 8820 12116 8854
rect 12150 8820 12184 8854
rect 12218 8820 12252 8854
rect 12286 8820 12320 8854
rect 12354 8820 12388 8854
rect 12422 8820 12456 8854
rect 12490 8820 12524 8854
rect 12558 8820 12592 8854
rect 12626 8820 12660 8854
rect 12694 8820 12728 8854
rect 12762 8820 12796 8854
rect 12830 8820 12864 8854
rect 12898 8820 12932 8854
rect 12966 8820 13000 8854
rect 13034 8820 13068 8854
rect 13102 8820 13118 8854
rect 1837 7579 1946 7618
rect 2048 7579 2056 7618
rect 1837 7545 1944 7579
rect 2050 7545 2056 7579
rect 1837 6560 1946 7545
rect 2048 6560 2056 7545
rect 2958 8714 3060 8726
rect 3512 8714 3614 8726
rect 4066 8714 4168 8726
rect 4620 8714 4722 8726
rect 5174 8714 5276 8726
rect 5728 8714 5830 8726
rect 6282 8714 6384 8726
rect 6836 8714 6938 8726
rect 7390 8714 7492 8726
rect 7944 8714 8046 8726
rect 8498 8714 8600 8726
rect 9052 8714 9154 8726
rect 9606 8714 9708 8726
rect 10160 8714 10262 8726
rect 10714 8714 10816 8726
rect 11268 8714 11370 8726
rect 11822 8714 11924 8726
rect 12376 8714 12478 8726
rect 12930 8714 13032 8726
rect 2255 8651 2274 8690
rect 2255 8577 2274 8617
rect 2255 8503 2274 8543
rect 2255 8429 2274 8469
rect 2255 8355 2274 8395
rect 2255 8281 2274 8321
rect 2255 8207 2274 8247
rect 2255 8133 2274 8173
rect 2255 8059 2274 8099
rect 2255 7985 2274 8025
rect 2255 7911 2274 7951
rect 2255 7837 2274 7877
rect 2255 7763 2274 7803
rect 2255 7689 2274 7729
rect 2255 7615 2274 7655
rect 2255 7541 2274 7581
rect 2255 7467 2274 7507
rect 2255 7393 2274 7433
rect 2713 8680 2751 8714
rect 2679 8641 2785 8680
rect 2713 8607 2751 8641
rect 2679 8568 2785 8607
rect 2713 8534 2751 8568
rect 2679 8495 2785 8534
rect 2713 8461 2751 8495
rect 2679 8422 2785 8461
rect 2990 8680 3028 8714
rect 2956 8641 3062 8680
rect 2990 8607 3028 8641
rect 2956 8568 3062 8607
rect 2990 8534 3028 8568
rect 2956 8495 3062 8534
rect 2990 8461 3028 8495
rect 2956 8422 3062 8461
rect 3267 8680 3305 8714
rect 3233 8641 3339 8680
rect 3267 8607 3305 8641
rect 3233 8568 3339 8607
rect 3267 8534 3305 8568
rect 3233 8495 3339 8534
rect 3267 8461 3305 8495
rect 3233 8422 3339 8461
rect 3544 8680 3582 8714
rect 3510 8641 3616 8680
rect 3544 8607 3582 8641
rect 3510 8568 3616 8607
rect 3544 8534 3582 8568
rect 3510 8495 3616 8534
rect 3544 8461 3582 8495
rect 3510 8422 3616 8461
rect 3821 8680 3859 8714
rect 3787 8641 3893 8680
rect 3821 8607 3859 8641
rect 3787 8568 3893 8607
rect 3821 8534 3859 8568
rect 3787 8495 3893 8534
rect 3821 8461 3859 8495
rect 3787 8422 3893 8461
rect 4098 8680 4136 8714
rect 4064 8641 4170 8680
rect 4098 8607 4136 8641
rect 4064 8568 4170 8607
rect 4098 8534 4136 8568
rect 4064 8495 4170 8534
rect 4098 8461 4136 8495
rect 4064 8422 4170 8461
rect 4375 8680 4413 8714
rect 4341 8641 4447 8680
rect 4375 8607 4413 8641
rect 4341 8568 4447 8607
rect 4375 8534 4413 8568
rect 4341 8495 4447 8534
rect 4375 8461 4413 8495
rect 4341 8422 4447 8461
rect 4652 8680 4690 8714
rect 4618 8641 4724 8680
rect 4652 8607 4690 8641
rect 4618 8568 4724 8607
rect 4652 8534 4690 8568
rect 4618 8495 4724 8534
rect 4652 8461 4690 8495
rect 4618 8422 4724 8461
rect 4929 8680 4967 8714
rect 4895 8641 5001 8680
rect 4929 8607 4967 8641
rect 4895 8568 5001 8607
rect 4929 8534 4967 8568
rect 4895 8495 5001 8534
rect 4929 8461 4967 8495
rect 4895 8422 5001 8461
rect 5206 8680 5244 8714
rect 5172 8641 5278 8680
rect 5206 8607 5244 8641
rect 5172 8568 5278 8607
rect 5206 8534 5244 8568
rect 5172 8495 5278 8534
rect 5206 8461 5244 8495
rect 5172 8422 5278 8461
rect 5483 8680 5521 8714
rect 5449 8641 5555 8680
rect 5483 8607 5521 8641
rect 5449 8568 5555 8607
rect 5483 8534 5521 8568
rect 5449 8495 5555 8534
rect 5483 8461 5521 8495
rect 5449 8422 5555 8461
rect 5760 8680 5798 8714
rect 5726 8641 5832 8680
rect 5760 8607 5798 8641
rect 5726 8568 5832 8607
rect 5760 8534 5798 8568
rect 5726 8495 5832 8534
rect 5760 8461 5798 8495
rect 5726 8422 5832 8461
rect 6037 8680 6075 8714
rect 6003 8641 6109 8680
rect 6037 8607 6075 8641
rect 6003 8568 6109 8607
rect 6037 8534 6075 8568
rect 6003 8495 6109 8534
rect 6037 8461 6075 8495
rect 6003 8422 6109 8461
rect 6314 8680 6352 8714
rect 6280 8641 6386 8680
rect 6314 8607 6352 8641
rect 6280 8568 6386 8607
rect 6314 8534 6352 8568
rect 6280 8495 6386 8534
rect 6314 8461 6352 8495
rect 6280 8422 6386 8461
rect 6591 8680 6629 8714
rect 6557 8641 6663 8680
rect 6591 8607 6629 8641
rect 6557 8568 6663 8607
rect 6591 8534 6629 8568
rect 6557 8495 6663 8534
rect 6591 8461 6629 8495
rect 6557 8422 6663 8461
rect 6868 8680 6906 8714
rect 6834 8641 6940 8680
rect 6868 8607 6906 8641
rect 6834 8568 6940 8607
rect 6868 8534 6906 8568
rect 6834 8495 6940 8534
rect 6868 8461 6906 8495
rect 6834 8422 6940 8461
rect 7145 8680 7183 8714
rect 7111 8641 7217 8680
rect 7145 8607 7183 8641
rect 7111 8568 7217 8607
rect 7145 8534 7183 8568
rect 7111 8495 7217 8534
rect 7145 8461 7183 8495
rect 7111 8422 7217 8461
rect 7422 8680 7460 8714
rect 7388 8641 7494 8680
rect 7422 8607 7460 8641
rect 7388 8568 7494 8607
rect 7422 8534 7460 8568
rect 7388 8495 7494 8534
rect 7422 8461 7460 8495
rect 7388 8422 7494 8461
rect 7699 8680 7737 8714
rect 7665 8641 7771 8680
rect 7699 8607 7737 8641
rect 7665 8568 7771 8607
rect 7699 8534 7737 8568
rect 7665 8495 7771 8534
rect 7699 8461 7737 8495
rect 7665 8422 7771 8461
rect 7976 8680 8014 8714
rect 7942 8641 8048 8680
rect 7976 8607 8014 8641
rect 7942 8568 8048 8607
rect 7976 8534 8014 8568
rect 7942 8495 8048 8534
rect 7976 8461 8014 8495
rect 7942 8422 8048 8461
rect 8253 8680 8291 8714
rect 8219 8641 8325 8680
rect 8253 8607 8291 8641
rect 8219 8568 8325 8607
rect 8253 8534 8291 8568
rect 8219 8495 8325 8534
rect 8253 8461 8291 8495
rect 8219 8422 8325 8461
rect 8530 8680 8568 8714
rect 8496 8641 8602 8680
rect 8530 8607 8568 8641
rect 8496 8568 8602 8607
rect 8530 8534 8568 8568
rect 8496 8495 8602 8534
rect 8530 8461 8568 8495
rect 8496 8422 8602 8461
rect 8807 8680 8845 8714
rect 8773 8641 8879 8680
rect 8807 8607 8845 8641
rect 8773 8568 8879 8607
rect 8807 8534 8845 8568
rect 8773 8495 8879 8534
rect 8807 8461 8845 8495
rect 8773 8422 8879 8461
rect 9084 8680 9122 8714
rect 9050 8641 9156 8680
rect 9084 8607 9122 8641
rect 9050 8568 9156 8607
rect 9084 8534 9122 8568
rect 9050 8495 9156 8534
rect 9084 8461 9122 8495
rect 9050 8422 9156 8461
rect 9361 8680 9399 8714
rect 9327 8641 9433 8680
rect 9361 8607 9399 8641
rect 9327 8568 9433 8607
rect 9361 8534 9399 8568
rect 9327 8495 9433 8534
rect 9361 8461 9399 8495
rect 9327 8422 9433 8461
rect 9638 8680 9676 8714
rect 9604 8641 9710 8680
rect 9638 8607 9676 8641
rect 9604 8568 9710 8607
rect 9638 8534 9676 8568
rect 9604 8495 9710 8534
rect 9638 8461 9676 8495
rect 9604 8422 9710 8461
rect 9915 8680 9953 8714
rect 9881 8641 9987 8680
rect 9915 8607 9953 8641
rect 9881 8568 9987 8607
rect 9915 8534 9953 8568
rect 9881 8495 9987 8534
rect 9915 8461 9953 8495
rect 9881 8422 9987 8461
rect 10192 8680 10230 8714
rect 10158 8641 10264 8680
rect 10192 8607 10230 8641
rect 10158 8568 10264 8607
rect 10192 8534 10230 8568
rect 10158 8495 10264 8534
rect 10192 8461 10230 8495
rect 10158 8422 10264 8461
rect 10469 8680 10507 8714
rect 10435 8641 10541 8680
rect 10469 8607 10507 8641
rect 10435 8568 10541 8607
rect 10469 8534 10507 8568
rect 10435 8495 10541 8534
rect 10469 8461 10507 8495
rect 10435 8422 10541 8461
rect 10746 8680 10784 8714
rect 10712 8641 10818 8680
rect 10746 8607 10784 8641
rect 10712 8568 10818 8607
rect 10746 8534 10784 8568
rect 10712 8495 10818 8534
rect 10746 8461 10784 8495
rect 10712 8422 10818 8461
rect 11023 8680 11061 8714
rect 10989 8641 11095 8680
rect 11023 8607 11061 8641
rect 10989 8568 11095 8607
rect 11023 8534 11061 8568
rect 10989 8495 11095 8534
rect 11023 8461 11061 8495
rect 10989 8422 11095 8461
rect 11300 8680 11338 8714
rect 11266 8641 11372 8680
rect 11300 8607 11338 8641
rect 11266 8568 11372 8607
rect 11300 8534 11338 8568
rect 11266 8495 11372 8534
rect 11300 8461 11338 8495
rect 11266 8422 11372 8461
rect 11577 8680 11615 8714
rect 11543 8641 11649 8680
rect 11577 8607 11615 8641
rect 11543 8568 11649 8607
rect 11577 8534 11615 8568
rect 11543 8495 11649 8534
rect 11577 8461 11615 8495
rect 11543 8422 11649 8461
rect 11854 8680 11892 8714
rect 11820 8641 11926 8680
rect 11854 8607 11892 8641
rect 11820 8568 11926 8607
rect 11854 8534 11892 8568
rect 11820 8495 11926 8534
rect 11854 8461 11892 8495
rect 11820 8422 11926 8461
rect 12131 8680 12169 8714
rect 12097 8641 12203 8680
rect 12131 8607 12169 8641
rect 12097 8568 12203 8607
rect 12131 8534 12169 8568
rect 12097 8495 12203 8534
rect 12131 8461 12169 8495
rect 12097 8422 12203 8461
rect 12408 8680 12446 8714
rect 12374 8641 12480 8680
rect 12408 8607 12446 8641
rect 12374 8568 12480 8607
rect 12408 8534 12446 8568
rect 12374 8495 12480 8534
rect 12408 8461 12446 8495
rect 12374 8422 12480 8461
rect 12685 8680 12723 8714
rect 12651 8641 12757 8680
rect 12685 8607 12723 8641
rect 12651 8568 12757 8607
rect 12685 8534 12723 8568
rect 12651 8495 12757 8534
rect 12685 8461 12723 8495
rect 12651 8422 12757 8461
rect 12962 8680 13000 8714
rect 12928 8641 13034 8680
rect 12962 8607 13000 8641
rect 12928 8568 13034 8607
rect 12962 8534 13000 8568
rect 12928 8495 13034 8534
rect 12962 8461 13000 8495
rect 12928 8422 13034 8461
rect 13239 8680 13277 8714
rect 13205 8641 13311 8680
rect 13239 8607 13277 8641
rect 13205 8568 13311 8607
rect 13239 8534 13277 8568
rect 13205 8495 13311 8534
rect 13239 8461 13277 8495
rect 13205 8422 13311 8461
rect 2958 7368 3060 7380
rect 3512 7368 3614 7380
rect 4066 7368 4168 7380
rect 4620 7368 4722 7380
rect 5174 7368 5276 7380
rect 5728 7368 5830 7380
rect 6282 7368 6384 7380
rect 6836 7368 6938 7380
rect 7390 7368 7492 7380
rect 7944 7368 8046 7380
rect 8498 7368 8600 7380
rect 9052 7368 9154 7380
rect 9606 7368 9708 7380
rect 10160 7368 10262 7380
rect 10714 7368 10816 7380
rect 11268 7368 11370 7380
rect 11822 7368 11924 7380
rect 12376 7368 12478 7380
rect 12930 7368 13032 7380
rect 2255 7349 2274 7359
rect 2638 7290 2888 7324
rect 2922 7290 2957 7324
rect 2991 7290 3026 7324
rect 3060 7290 3095 7324
rect 3129 7290 3164 7324
rect 3198 7290 3233 7324
rect 3267 7290 3302 7324
rect 3336 7290 3371 7324
rect 3405 7290 3440 7324
rect 3474 7290 3509 7324
rect 3543 7290 3578 7324
rect 3612 7290 3647 7324
rect 3681 7290 3716 7324
rect 3750 7290 3785 7324
rect 3819 7290 3854 7324
rect 3888 7290 3923 7324
rect 3957 7290 3992 7324
rect 4026 7290 4061 7324
rect 4095 7290 4130 7324
rect 4164 7290 4199 7324
rect 4233 7290 4268 7324
rect 4302 7290 4337 7324
rect 4371 7290 4406 7324
rect 4440 7290 4475 7324
rect 4509 7290 4544 7324
rect 4578 7290 4613 7324
rect 4647 7290 4682 7324
rect 4716 7290 4751 7324
rect 4785 7290 4820 7324
rect 4854 7290 4889 7324
rect 4923 7290 4958 7324
rect 4992 7290 5027 7324
rect 5061 7290 5096 7324
rect 5130 7290 5165 7324
rect 5199 7290 5234 7324
rect 5268 7290 5303 7324
rect 5337 7290 5372 7324
rect 5406 7290 5441 7324
rect 5475 7290 5510 7324
rect 5544 7290 5579 7324
rect 5613 7290 5648 7324
rect 5682 7290 5717 7324
rect 5751 7290 5786 7324
rect 5820 7290 5855 7324
rect 5889 7290 5924 7324
rect 5958 7290 5993 7324
rect 6027 7290 6062 7324
rect 6096 7290 6131 7324
rect 6165 7290 6200 7324
rect 6234 7290 6268 7324
rect 6302 7290 6336 7324
rect 6370 7290 6404 7324
rect 6438 7290 6472 7324
rect 6506 7290 6540 7324
rect 6574 7290 6608 7324
rect 6642 7290 6676 7324
rect 6710 7290 6744 7324
rect 6778 7290 6812 7324
rect 6846 7290 6880 7324
rect 6914 7290 6948 7324
rect 6982 7290 7016 7324
rect 7050 7290 7084 7324
rect 7118 7290 7152 7324
rect 7186 7290 7220 7324
rect 7254 7290 7288 7324
rect 7322 7290 7356 7324
rect 7390 7290 7424 7324
rect 7458 7290 7492 7324
rect 7526 7290 7560 7324
rect 7594 7290 7628 7324
rect 7662 7290 7696 7324
rect 7730 7290 7764 7324
rect 7798 7290 7832 7324
rect 7866 7290 7900 7324
rect 7934 7290 7968 7324
rect 8002 7290 8036 7324
rect 8070 7290 8104 7324
rect 8138 7290 8172 7324
rect 8206 7290 8240 7324
rect 8274 7290 8308 7324
rect 8342 7290 8376 7324
rect 8410 7290 8444 7324
rect 8478 7290 8512 7324
rect 8546 7290 8580 7324
rect 8614 7290 8648 7324
rect 8682 7290 8716 7324
rect 8750 7290 8784 7324
rect 8818 7290 8852 7324
rect 8886 7290 8920 7324
rect 8954 7290 8988 7324
rect 9022 7290 9056 7324
rect 9090 7290 9124 7324
rect 9158 7290 9192 7324
rect 9226 7290 9260 7324
rect 9294 7290 9328 7324
rect 9362 7290 9396 7324
rect 9430 7290 9464 7324
rect 9498 7290 9532 7324
rect 9566 7290 9600 7324
rect 9634 7290 9668 7324
rect 9702 7290 9736 7324
rect 9770 7290 9804 7324
rect 9838 7290 9872 7324
rect 9906 7290 9940 7324
rect 9974 7290 10008 7324
rect 10042 7290 10076 7324
rect 10110 7290 10144 7324
rect 10178 7290 10212 7324
rect 10246 7290 10280 7324
rect 10314 7290 10348 7324
rect 10382 7290 10416 7324
rect 10450 7290 10484 7324
rect 10518 7290 10552 7324
rect 10586 7290 10620 7324
rect 10654 7290 10688 7324
rect 10722 7290 10756 7324
rect 10790 7290 10824 7324
rect 10858 7290 10892 7324
rect 10926 7290 10960 7324
rect 10994 7290 11028 7324
rect 11062 7290 11096 7324
rect 11130 7290 11164 7324
rect 11198 7290 11232 7324
rect 11266 7290 11300 7324
rect 11334 7290 11368 7324
rect 11402 7290 11436 7324
rect 11470 7290 11504 7324
rect 11538 7290 11572 7324
rect 11606 7290 11640 7324
rect 11674 7290 11708 7324
rect 11742 7290 11776 7324
rect 11810 7290 11844 7324
rect 11878 7290 11912 7324
rect 11946 7290 11980 7324
rect 12014 7290 12048 7324
rect 12082 7290 12116 7324
rect 12150 7290 12184 7324
rect 12218 7290 12252 7324
rect 12286 7290 12320 7324
rect 12354 7290 12388 7324
rect 12422 7290 12456 7324
rect 12490 7290 12524 7324
rect 12558 7290 12592 7324
rect 12626 7290 12660 7324
rect 12694 7290 12728 7324
rect 12762 7290 12796 7324
rect 12830 7290 12864 7324
rect 12898 7290 12932 7324
rect 12966 7290 13000 7324
rect 13034 7290 13068 7324
rect 13102 7290 13118 7324
rect 2638 7243 13118 7290
rect 2672 7209 2710 7243
rect 2744 7209 13118 7243
rect 2638 7153 13118 7209
rect 2672 7119 2710 7153
rect 2744 7119 13118 7153
rect 2638 7063 13118 7119
rect 2672 7029 2710 7063
rect 2744 7029 13118 7063
rect 2638 6972 13118 7029
rect 2672 6938 2710 6972
rect 2744 6938 13118 6972
rect 2638 6854 13118 6938
rect 2638 6820 2888 6854
rect 2922 6820 2957 6854
rect 2991 6820 3026 6854
rect 3060 6820 3095 6854
rect 3129 6820 3164 6854
rect 3198 6820 3233 6854
rect 3267 6820 3302 6854
rect 3336 6820 3371 6854
rect 3405 6820 3440 6854
rect 3474 6820 3509 6854
rect 3543 6820 3578 6854
rect 3612 6820 3647 6854
rect 3681 6820 3716 6854
rect 3750 6820 3785 6854
rect 3819 6820 3854 6854
rect 3888 6820 3923 6854
rect 3957 6820 3992 6854
rect 4026 6820 4061 6854
rect 4095 6820 4130 6854
rect 4164 6820 4199 6854
rect 4233 6820 4268 6854
rect 4302 6820 4337 6854
rect 4371 6820 4406 6854
rect 4440 6820 4475 6854
rect 4509 6820 4544 6854
rect 4578 6820 4613 6854
rect 4647 6820 4682 6854
rect 4716 6820 4751 6854
rect 4785 6820 4820 6854
rect 4854 6820 4889 6854
rect 4923 6820 4958 6854
rect 4992 6820 5027 6854
rect 5061 6820 5096 6854
rect 5130 6820 5165 6854
rect 5199 6820 5234 6854
rect 5268 6820 5303 6854
rect 5337 6820 5372 6854
rect 5406 6820 5441 6854
rect 5475 6820 5510 6854
rect 5544 6820 5579 6854
rect 5613 6820 5648 6854
rect 5682 6820 5717 6854
rect 5751 6820 5786 6854
rect 5820 6820 5855 6854
rect 5889 6820 5924 6854
rect 5958 6820 5993 6854
rect 6027 6820 6062 6854
rect 6096 6820 6131 6854
rect 6165 6820 6200 6854
rect 6234 6820 6268 6854
rect 6302 6820 6336 6854
rect 6370 6820 6404 6854
rect 6438 6820 6472 6854
rect 6506 6820 6540 6854
rect 6574 6820 6608 6854
rect 6642 6820 6676 6854
rect 6710 6820 6744 6854
rect 6778 6820 6812 6854
rect 6846 6820 6880 6854
rect 6914 6820 6948 6854
rect 6982 6820 7016 6854
rect 7050 6820 7084 6854
rect 7118 6820 7152 6854
rect 7186 6820 7220 6854
rect 7254 6820 7288 6854
rect 7322 6820 7356 6854
rect 7390 6820 7424 6854
rect 7458 6820 7492 6854
rect 7526 6820 7560 6854
rect 7594 6820 7628 6854
rect 7662 6820 7696 6854
rect 7730 6820 7764 6854
rect 7798 6820 7832 6854
rect 7866 6820 7900 6854
rect 7934 6820 7968 6854
rect 8002 6820 8036 6854
rect 8070 6820 8104 6854
rect 8138 6820 8172 6854
rect 8206 6820 8240 6854
rect 8274 6820 8308 6854
rect 8342 6820 8376 6854
rect 8410 6820 8444 6854
rect 8478 6820 8512 6854
rect 8546 6820 8580 6854
rect 8614 6820 8648 6854
rect 8682 6820 8716 6854
rect 8750 6820 8784 6854
rect 8818 6820 8852 6854
rect 8886 6820 8920 6854
rect 8954 6820 8988 6854
rect 9022 6820 9056 6854
rect 9090 6820 9124 6854
rect 9158 6820 9192 6854
rect 9226 6820 9260 6854
rect 9294 6820 9328 6854
rect 9362 6820 9396 6854
rect 9430 6820 9464 6854
rect 9498 6820 9532 6854
rect 9566 6820 9600 6854
rect 9634 6820 9668 6854
rect 9702 6820 9736 6854
rect 9770 6820 9804 6854
rect 9838 6820 9872 6854
rect 9906 6820 9940 6854
rect 9974 6820 10008 6854
rect 10042 6820 10076 6854
rect 10110 6820 10144 6854
rect 10178 6820 10212 6854
rect 10246 6820 10280 6854
rect 10314 6820 10348 6854
rect 10382 6820 10416 6854
rect 10450 6820 10484 6854
rect 10518 6820 10552 6854
rect 10586 6820 10620 6854
rect 10654 6820 10688 6854
rect 10722 6820 10756 6854
rect 10790 6820 10824 6854
rect 10858 6820 10892 6854
rect 10926 6820 10960 6854
rect 10994 6820 11028 6854
rect 11062 6820 11096 6854
rect 11130 6820 11164 6854
rect 11198 6820 11232 6854
rect 11266 6820 11300 6854
rect 11334 6820 11368 6854
rect 11402 6820 11436 6854
rect 11470 6820 11504 6854
rect 11538 6820 11572 6854
rect 11606 6820 11640 6854
rect 11674 6820 11708 6854
rect 11742 6820 11776 6854
rect 11810 6820 11844 6854
rect 11878 6820 11912 6854
rect 11946 6820 11980 6854
rect 12014 6820 12048 6854
rect 12082 6820 12116 6854
rect 12150 6820 12184 6854
rect 12218 6820 12252 6854
rect 12286 6820 12320 6854
rect 12354 6820 12388 6854
rect 12422 6820 12456 6854
rect 12490 6820 12524 6854
rect 12558 6820 12592 6854
rect 12626 6820 12660 6854
rect 12694 6820 12728 6854
rect 12762 6820 12796 6854
rect 12830 6820 12864 6854
rect 12898 6820 12932 6854
rect 12966 6820 13000 6854
rect 13034 6820 13068 6854
rect 13102 6820 13118 6854
rect 1837 6526 1944 6560
rect 2050 6526 2056 6560
rect 1837 6487 1946 6526
rect 2048 6487 2056 6526
rect 1837 6453 1944 6487
rect 2050 6453 2056 6487
rect 1837 6414 1946 6453
rect 2048 6414 2056 6453
rect 1837 6380 1944 6414
rect 2050 6380 2056 6414
rect 1837 6341 1946 6380
rect 2048 6341 2056 6380
rect 1837 6307 1944 6341
rect 2050 6307 2056 6341
rect 1837 6268 1946 6307
rect 2048 6268 2056 6307
rect 1837 6234 1944 6268
rect 2050 6234 2056 6268
rect 1837 6195 1946 6234
rect 2048 6195 2056 6234
rect 1837 6161 1944 6195
rect 2050 6161 2056 6195
rect 1837 6122 1946 6161
rect 2048 6122 2056 6161
rect 1837 6088 1944 6122
rect 2050 6088 2056 6122
rect 1837 6049 1946 6088
rect 2048 6049 2056 6088
rect 1837 6015 1944 6049
rect 2050 6015 2056 6049
rect 1837 5976 1946 6015
rect 2048 5976 2056 6015
rect 1837 5942 1944 5976
rect 2050 5942 2056 5976
rect 1837 5903 1946 5942
rect 2048 5903 2056 5942
rect 1837 5869 1944 5903
rect 2050 5869 2056 5903
rect 1837 5830 1946 5869
rect 2048 5830 2056 5869
rect 1837 5796 1944 5830
rect 2050 5796 2056 5830
rect 1837 5757 1946 5796
rect 2048 5757 2056 5796
rect 1837 5723 1944 5757
rect 2050 5723 2056 5757
rect 1837 5683 1946 5723
rect 2048 5683 2056 5723
rect 1837 5649 1944 5683
rect 2050 5649 2056 5683
rect 1837 5609 1946 5649
rect 2048 5609 2056 5649
rect 1837 5575 1944 5609
rect 2050 5575 2056 5609
rect 1837 5535 1946 5575
rect 2048 5535 2056 5575
rect 1837 5501 1944 5535
rect 1978 5501 2016 5508
rect 2050 5501 2056 5535
rect 1837 5461 2056 5501
rect 1837 5427 1944 5461
rect 1978 5427 2016 5461
rect 2050 5427 2056 5461
rect 1837 5387 2056 5427
rect 1837 5353 1944 5387
rect 1978 5353 2016 5387
rect 2050 5353 2056 5387
rect 1837 5345 2056 5353
rect 1837 5313 1946 5345
rect 2048 5313 2056 5345
rect 1837 5279 1944 5313
rect 2050 5279 2056 5313
rect 1837 5239 1946 5279
rect 2048 5239 2056 5279
rect 1837 5205 1944 5239
rect 2050 5205 2056 5239
rect 1837 5165 1946 5205
rect 2048 5165 2056 5205
rect 1837 5131 1944 5165
rect 2050 5131 2056 5165
rect 1837 5091 1946 5131
rect 2048 5091 2056 5131
rect 1837 5057 1944 5091
rect 2050 5057 2056 5091
rect 1837 5017 1946 5057
rect 2048 5017 2056 5057
rect 1837 4983 1944 5017
rect 2050 4983 2056 5017
rect 2255 6735 2274 6774
rect 2958 6714 3060 6726
rect 3512 6714 3614 6726
rect 4066 6714 4168 6726
rect 4620 6714 4722 6726
rect 5174 6714 5276 6726
rect 5728 6714 5830 6726
rect 6282 6714 6384 6726
rect 6836 6714 6938 6726
rect 7390 6714 7492 6726
rect 7944 6714 8046 6726
rect 8498 6714 8600 6726
rect 9052 6714 9154 6726
rect 9606 6714 9708 6726
rect 10160 6714 10262 6726
rect 10714 6714 10816 6726
rect 11268 6714 11370 6726
rect 11822 6714 11924 6726
rect 12376 6714 12478 6726
rect 12930 6714 13032 6726
rect 2255 6662 2274 6701
rect 2255 6589 2274 6628
rect 2255 6516 2274 6555
rect 2255 6443 2274 6482
rect 2255 6370 2274 6409
rect 2255 6297 2274 6336
rect 2255 6224 2274 6263
rect 2255 6151 2274 6190
rect 2255 6078 2274 6117
rect 2255 6005 2274 6044
rect 2255 5932 2274 5971
rect 2255 5859 2274 5898
rect 2255 5786 2274 5825
rect 2255 5713 2274 5752
rect 2255 5640 2274 5679
rect 2255 5567 2274 5606
rect 2255 5494 2274 5533
rect 2255 5421 2274 5460
rect 2255 5348 2274 5387
rect 2713 6680 2751 6714
rect 2679 6641 2785 6680
rect 2713 6607 2751 6641
rect 2679 6568 2785 6607
rect 2713 6534 2751 6568
rect 2679 6495 2785 6534
rect 2713 6461 2751 6495
rect 2679 6422 2785 6461
rect 2990 6680 3028 6714
rect 2956 6641 3062 6680
rect 2990 6607 3028 6641
rect 2956 6568 3062 6607
rect 2990 6534 3028 6568
rect 2956 6495 3062 6534
rect 2990 6461 3028 6495
rect 2956 6422 3062 6461
rect 3267 6680 3305 6714
rect 3233 6641 3339 6680
rect 3267 6607 3305 6641
rect 3233 6568 3339 6607
rect 3267 6534 3305 6568
rect 3233 6495 3339 6534
rect 3267 6461 3305 6495
rect 3233 6422 3339 6461
rect 3544 6680 3582 6714
rect 3510 6641 3616 6680
rect 3544 6607 3582 6641
rect 3510 6568 3616 6607
rect 3544 6534 3582 6568
rect 3510 6495 3616 6534
rect 3544 6461 3582 6495
rect 3510 6422 3616 6461
rect 3821 6680 3859 6714
rect 3787 6641 3893 6680
rect 3821 6607 3859 6641
rect 3787 6568 3893 6607
rect 3821 6534 3859 6568
rect 3787 6495 3893 6534
rect 3821 6461 3859 6495
rect 3787 6422 3893 6461
rect 4098 6680 4136 6714
rect 4064 6641 4170 6680
rect 4098 6607 4136 6641
rect 4064 6568 4170 6607
rect 4098 6534 4136 6568
rect 4064 6495 4170 6534
rect 4098 6461 4136 6495
rect 4064 6422 4170 6461
rect 4375 6680 4413 6714
rect 4341 6641 4447 6680
rect 4375 6607 4413 6641
rect 4341 6568 4447 6607
rect 4375 6534 4413 6568
rect 4341 6495 4447 6534
rect 4375 6461 4413 6495
rect 4341 6422 4447 6461
rect 4652 6680 4690 6714
rect 4618 6641 4724 6680
rect 4652 6607 4690 6641
rect 4618 6568 4724 6607
rect 4652 6534 4690 6568
rect 4618 6495 4724 6534
rect 4652 6461 4690 6495
rect 4618 6422 4724 6461
rect 4929 6680 4967 6714
rect 4895 6641 5001 6680
rect 4929 6607 4967 6641
rect 4895 6568 5001 6607
rect 4929 6534 4967 6568
rect 4895 6495 5001 6534
rect 4929 6461 4967 6495
rect 4895 6422 5001 6461
rect 5206 6680 5244 6714
rect 5172 6641 5278 6680
rect 5206 6607 5244 6641
rect 5172 6568 5278 6607
rect 5206 6534 5244 6568
rect 5172 6495 5278 6534
rect 5206 6461 5244 6495
rect 5172 6422 5278 6461
rect 5483 6680 5521 6714
rect 5449 6641 5555 6680
rect 5483 6607 5521 6641
rect 5449 6568 5555 6607
rect 5483 6534 5521 6568
rect 5449 6495 5555 6534
rect 5483 6461 5521 6495
rect 5449 6422 5555 6461
rect 5760 6680 5798 6714
rect 5726 6641 5832 6680
rect 5760 6607 5798 6641
rect 5726 6568 5832 6607
rect 5760 6534 5798 6568
rect 5726 6495 5832 6534
rect 5760 6461 5798 6495
rect 5726 6422 5832 6461
rect 6037 6680 6075 6714
rect 6003 6641 6109 6680
rect 6037 6607 6075 6641
rect 6003 6568 6109 6607
rect 6037 6534 6075 6568
rect 6003 6495 6109 6534
rect 6037 6461 6075 6495
rect 6003 6422 6109 6461
rect 6314 6680 6352 6714
rect 6280 6641 6386 6680
rect 6314 6607 6352 6641
rect 6280 6568 6386 6607
rect 6314 6534 6352 6568
rect 6280 6495 6386 6534
rect 6314 6461 6352 6495
rect 6280 6422 6386 6461
rect 6591 6680 6629 6714
rect 6557 6641 6663 6680
rect 6591 6607 6629 6641
rect 6557 6568 6663 6607
rect 6591 6534 6629 6568
rect 6557 6495 6663 6534
rect 6591 6461 6629 6495
rect 6557 6422 6663 6461
rect 6868 6680 6906 6714
rect 6834 6641 6940 6680
rect 6868 6607 6906 6641
rect 6834 6568 6940 6607
rect 6868 6534 6906 6568
rect 6834 6495 6940 6534
rect 6868 6461 6906 6495
rect 6834 6422 6940 6461
rect 7145 6680 7183 6714
rect 7111 6641 7217 6680
rect 7145 6607 7183 6641
rect 7111 6568 7217 6607
rect 7145 6534 7183 6568
rect 7111 6495 7217 6534
rect 7145 6461 7183 6495
rect 7111 6422 7217 6461
rect 7422 6680 7460 6714
rect 7388 6641 7494 6680
rect 7422 6607 7460 6641
rect 7388 6568 7494 6607
rect 7422 6534 7460 6568
rect 7388 6495 7494 6534
rect 7422 6461 7460 6495
rect 7388 6422 7494 6461
rect 7699 6680 7737 6714
rect 7665 6641 7771 6680
rect 7699 6607 7737 6641
rect 7665 6568 7771 6607
rect 7699 6534 7737 6568
rect 7665 6495 7771 6534
rect 7699 6461 7737 6495
rect 7665 6422 7771 6461
rect 7976 6680 8014 6714
rect 7942 6641 8048 6680
rect 7976 6607 8014 6641
rect 7942 6568 8048 6607
rect 7976 6534 8014 6568
rect 7942 6495 8048 6534
rect 7976 6461 8014 6495
rect 7942 6422 8048 6461
rect 8253 6680 8291 6714
rect 8219 6641 8325 6680
rect 8253 6607 8291 6641
rect 8219 6568 8325 6607
rect 8253 6534 8291 6568
rect 8219 6495 8325 6534
rect 8253 6461 8291 6495
rect 8219 6422 8325 6461
rect 8530 6680 8568 6714
rect 8496 6641 8602 6680
rect 8530 6607 8568 6641
rect 8496 6568 8602 6607
rect 8530 6534 8568 6568
rect 8496 6495 8602 6534
rect 8530 6461 8568 6495
rect 8496 6422 8602 6461
rect 8807 6680 8845 6714
rect 8773 6641 8879 6680
rect 8807 6607 8845 6641
rect 8773 6568 8879 6607
rect 8807 6534 8845 6568
rect 8773 6495 8879 6534
rect 8807 6461 8845 6495
rect 8773 6422 8879 6461
rect 9084 6680 9122 6714
rect 9050 6641 9156 6680
rect 9084 6607 9122 6641
rect 9050 6568 9156 6607
rect 9084 6534 9122 6568
rect 9050 6495 9156 6534
rect 9084 6461 9122 6495
rect 9050 6422 9156 6461
rect 9361 6680 9399 6714
rect 9327 6641 9433 6680
rect 9361 6607 9399 6641
rect 9327 6568 9433 6607
rect 9361 6534 9399 6568
rect 9327 6495 9433 6534
rect 9361 6461 9399 6495
rect 9327 6422 9433 6461
rect 9638 6680 9676 6714
rect 9604 6641 9710 6680
rect 9638 6607 9676 6641
rect 9604 6568 9710 6607
rect 9638 6534 9676 6568
rect 9604 6495 9710 6534
rect 9638 6461 9676 6495
rect 9604 6422 9710 6461
rect 9915 6680 9953 6714
rect 9881 6641 9987 6680
rect 9915 6607 9953 6641
rect 9881 6568 9987 6607
rect 9915 6534 9953 6568
rect 9881 6495 9987 6534
rect 9915 6461 9953 6495
rect 9881 6422 9987 6461
rect 10192 6680 10230 6714
rect 10158 6641 10264 6680
rect 10192 6607 10230 6641
rect 10158 6568 10264 6607
rect 10192 6534 10230 6568
rect 10158 6495 10264 6534
rect 10192 6461 10230 6495
rect 10158 6422 10264 6461
rect 10469 6680 10507 6714
rect 10435 6641 10541 6680
rect 10469 6607 10507 6641
rect 10435 6568 10541 6607
rect 10469 6534 10507 6568
rect 10435 6495 10541 6534
rect 10469 6461 10507 6495
rect 10435 6422 10541 6461
rect 10746 6680 10784 6714
rect 10712 6641 10818 6680
rect 10746 6607 10784 6641
rect 10712 6568 10818 6607
rect 10746 6534 10784 6568
rect 10712 6495 10818 6534
rect 10746 6461 10784 6495
rect 10712 6422 10818 6461
rect 11023 6680 11061 6714
rect 10989 6641 11095 6680
rect 11023 6607 11061 6641
rect 10989 6568 11095 6607
rect 11023 6534 11061 6568
rect 10989 6495 11095 6534
rect 11023 6461 11061 6495
rect 10989 6422 11095 6461
rect 11300 6680 11338 6714
rect 11266 6641 11372 6680
rect 11300 6607 11338 6641
rect 11266 6568 11372 6607
rect 11300 6534 11338 6568
rect 11266 6495 11372 6534
rect 11300 6461 11338 6495
rect 11266 6422 11372 6461
rect 11577 6680 11615 6714
rect 11543 6641 11649 6680
rect 11577 6607 11615 6641
rect 11543 6568 11649 6607
rect 11577 6534 11615 6568
rect 11543 6495 11649 6534
rect 11577 6461 11615 6495
rect 11543 6422 11649 6461
rect 11854 6680 11892 6714
rect 11820 6641 11926 6680
rect 11854 6607 11892 6641
rect 11820 6568 11926 6607
rect 11854 6534 11892 6568
rect 11820 6495 11926 6534
rect 11854 6461 11892 6495
rect 11820 6422 11926 6461
rect 12131 6680 12169 6714
rect 12097 6641 12203 6680
rect 12131 6607 12169 6641
rect 12097 6568 12203 6607
rect 12131 6534 12169 6568
rect 12097 6495 12203 6534
rect 12131 6461 12169 6495
rect 12097 6422 12203 6461
rect 12408 6680 12446 6714
rect 12374 6641 12480 6680
rect 12408 6607 12446 6641
rect 12374 6568 12480 6607
rect 12408 6534 12446 6568
rect 12374 6495 12480 6534
rect 12408 6461 12446 6495
rect 12374 6422 12480 6461
rect 12685 6680 12723 6714
rect 12651 6641 12757 6680
rect 12685 6607 12723 6641
rect 12651 6568 12757 6607
rect 12685 6534 12723 6568
rect 12651 6495 12757 6534
rect 12685 6461 12723 6495
rect 12651 6422 12757 6461
rect 12962 6680 13000 6714
rect 12928 6641 13034 6680
rect 12962 6607 13000 6641
rect 12928 6568 13034 6607
rect 12962 6534 13000 6568
rect 12928 6495 13034 6534
rect 12962 6461 13000 6495
rect 12928 6422 13034 6461
rect 13239 6680 13277 6714
rect 13205 6641 13311 6680
rect 13239 6607 13277 6641
rect 13205 6568 13311 6607
rect 13239 6534 13277 6568
rect 13205 6495 13311 6534
rect 13239 6461 13277 6495
rect 13205 6422 13311 6461
rect 2958 5368 3060 5380
rect 3512 5368 3614 5380
rect 4066 5368 4168 5380
rect 4620 5368 4722 5380
rect 5174 5368 5276 5380
rect 5728 5368 5830 5380
rect 6282 5368 6384 5380
rect 6836 5368 6938 5380
rect 7390 5368 7492 5380
rect 7944 5368 8046 5380
rect 8498 5368 8600 5380
rect 9052 5368 9154 5380
rect 9606 5368 9708 5380
rect 10160 5368 10262 5380
rect 10714 5368 10816 5380
rect 11268 5368 11370 5380
rect 11822 5368 11924 5380
rect 12376 5368 12478 5380
rect 12930 5368 13032 5380
rect 2255 5274 2274 5314
rect 2255 5129 2274 5240
rect 2444 5197 13458 5203
rect 2467 5183 2506 5197
rect 2540 5183 2579 5197
rect 2613 5183 2652 5197
rect 2686 5183 2725 5197
rect 2759 5183 2798 5197
rect 2832 5183 2871 5197
rect 2905 5183 2944 5197
rect 2978 5183 3017 5197
rect 3051 5183 3090 5197
rect 3124 5183 3163 5197
rect 3197 5183 3236 5197
rect 3270 5183 3309 5197
rect 3343 5183 3382 5197
rect 3416 5183 3455 5197
rect 3489 5183 3528 5197
rect 3562 5183 3601 5197
rect 3635 5183 3674 5197
rect 3708 5183 3747 5197
rect 3781 5183 3820 5197
rect 3854 5183 3893 5197
rect 3927 5183 3966 5197
rect 4000 5183 4039 5197
rect 4073 5183 4112 5197
rect 4146 5183 4185 5197
rect 4219 5183 4258 5197
rect 4292 5183 4331 5197
rect 4365 5183 4404 5197
rect 4438 5183 4477 5197
rect 4511 5183 4550 5197
rect 4584 5183 4623 5197
rect 4657 5183 4696 5197
rect 4730 5183 4769 5197
rect 4803 5183 4842 5197
rect 4876 5183 4915 5197
rect 4949 5183 4988 5197
rect 5022 5183 5061 5197
rect 5095 5183 5134 5197
rect 5168 5183 5207 5197
rect 5241 5183 5280 5197
rect 5314 5183 5353 5197
rect 5387 5183 5426 5197
rect 2255 5125 2478 5129
rect 2255 5091 2287 5125
rect 2321 5091 2360 5125
rect 2394 5091 2433 5125
rect 2467 5091 2478 5125
rect 2255 5081 2478 5091
rect 13452 5115 13458 5197
rect 13452 5085 13490 5115
rect 13524 5085 13562 5115
rect 13596 5085 13628 5115
rect 2255 5053 5426 5081
rect 2255 5019 2287 5053
rect 2321 5019 2360 5053
rect 2394 5019 2433 5053
rect 2467 5019 2506 5053
rect 2540 5019 2579 5053
rect 2613 5019 2652 5053
rect 2686 5019 2725 5053
rect 2759 5019 2798 5053
rect 2832 5019 2871 5053
rect 2905 5019 2944 5053
rect 2978 5019 3017 5053
rect 3051 5019 3090 5053
rect 3124 5019 3163 5053
rect 3197 5019 3236 5053
rect 3270 5019 3309 5053
rect 3343 5019 3382 5053
rect 3416 5019 3455 5053
rect 3489 5019 3528 5053
rect 3562 5019 3601 5053
rect 3635 5019 3674 5053
rect 3708 5019 3747 5053
rect 3781 5019 3820 5053
rect 3854 5019 3893 5053
rect 3927 5019 3966 5053
rect 4000 5019 4039 5053
rect 4073 5019 4112 5053
rect 4146 5019 4185 5053
rect 4219 5019 4258 5053
rect 4292 5019 4331 5053
rect 4365 5019 4404 5053
rect 4438 5019 4477 5053
rect 4511 5019 4550 5053
rect 4584 5019 4623 5053
rect 4657 5019 4696 5053
rect 4730 5019 4769 5053
rect 4803 5019 4842 5053
rect 4876 5019 4915 5053
rect 4949 5019 4988 5053
rect 5022 5019 5061 5053
rect 5095 5019 5134 5053
rect 5168 5019 5207 5053
rect 5241 5019 5280 5053
rect 5314 5019 5353 5053
rect 5387 5019 5426 5053
rect 13452 5019 13628 5085
rect 2255 5013 13628 5019
rect 13838 6856 13840 6895
rect 13942 6856 13944 6895
rect 13838 6783 13840 6822
rect 13942 6783 13944 6822
rect 13838 6710 13840 6749
rect 13942 6710 13944 6749
rect 13838 6637 13840 6676
rect 13942 6637 13944 6676
rect 13838 6564 13840 6603
rect 13942 6564 13944 6603
rect 13838 6491 13840 6530
rect 13942 6491 13944 6530
rect 13838 6418 13840 6457
rect 13942 6418 13944 6457
rect 13838 6345 13840 6384
rect 13942 6345 13944 6384
rect 13838 6272 13840 6311
rect 13942 6272 13944 6311
rect 13838 6199 13840 6238
rect 13942 6199 13944 6238
rect 13838 6126 13840 6165
rect 13942 6126 13944 6165
rect 13838 6053 13840 6092
rect 13942 6053 13944 6092
rect 13838 5980 13840 6019
rect 13942 5980 13944 6019
rect 13838 5907 13840 5946
rect 13942 5907 13944 5946
rect 13838 5834 13840 5873
rect 13942 5834 13944 5873
rect 13838 5761 13840 5800
rect 13942 5761 13944 5800
rect 13838 5688 13840 5727
rect 13942 5688 13944 5727
rect 13838 5615 13840 5654
rect 13942 5615 13944 5654
rect 13872 5581 13910 5593
rect 13838 5542 13944 5581
rect 13872 5508 13910 5542
rect 13838 5481 13944 5508
rect 13838 5469 13840 5481
rect 13942 5469 13944 5481
rect 13838 5396 13840 5435
rect 13942 5396 13944 5435
rect 13838 5323 13840 5362
rect 13942 5323 13944 5362
rect 13838 5250 13840 5289
rect 13942 5250 13944 5289
rect 13838 5177 13840 5216
rect 13942 5177 13944 5216
rect 13838 5104 13840 5143
rect 13942 5104 13944 5143
rect 13838 5031 13840 5070
rect 13942 5031 13944 5070
rect 1837 4943 1946 4983
rect 2048 4943 2056 4983
rect 1837 4909 1944 4943
rect 2050 4909 2056 4943
rect 1837 4835 1946 4909
rect 2048 4871 2056 4909
rect 13838 4958 13840 4997
rect 13942 4958 13944 4997
rect 13838 4885 13840 4924
rect 13942 4885 13944 4924
rect 2057 4869 2096 4871
rect 2130 4869 2169 4871
rect 2203 4869 2242 4871
rect 2276 4869 2315 4871
rect 2349 4869 2388 4871
rect 2422 4869 2461 4871
rect 2495 4869 2534 4871
rect 2568 4869 2607 4871
rect 2057 4837 2088 4869
rect 2598 4837 2607 4869
rect 2641 4869 2680 4871
rect 2714 4869 2753 4871
rect 2787 4869 2826 4871
rect 2860 4869 2899 4871
rect 2933 4869 2972 4871
rect 3006 4869 3045 4871
rect 3079 4869 3118 4871
rect 3152 4869 3191 4871
rect 3225 4869 3264 4871
rect 3298 4869 3337 4871
rect 3371 4869 3410 4871
rect 3444 4869 3483 4871
rect 3517 4869 3556 4871
rect 3590 4869 3629 4871
rect 3663 4869 3702 4871
rect 3736 4869 3775 4871
rect 3809 4869 3848 4871
rect 3882 4869 3921 4871
rect 3955 4869 3994 4871
rect 4028 4869 4067 4871
rect 4101 4869 4140 4871
rect 4174 4869 4213 4871
rect 4247 4869 4286 4871
rect 4320 4869 4359 4871
rect 4393 4869 4432 4871
rect 4466 4869 4505 4871
rect 4539 4869 4578 4871
rect 4612 4869 4651 4871
rect 4685 4869 4724 4871
rect 4758 4869 4797 4871
rect 4831 4869 4870 4871
rect 4904 4869 4943 4871
rect 4977 4869 5016 4871
rect 5050 4869 5089 4871
rect 5123 4869 5162 4871
rect 5196 4869 5235 4871
rect 13765 4869 13838 4871
rect 2641 4837 2666 4869
rect 2048 4835 2088 4837
rect 1837 4801 2088 4835
rect 1837 4799 2020 4801
rect 2054 4799 2088 4801
rect 2598 4799 2666 4837
rect 1837 4765 1950 4799
rect 1984 4767 2020 4799
rect 2057 4767 2088 4799
rect 2598 4767 2607 4799
rect 1984 4765 2023 4767
rect 2057 4765 2096 4767
rect 2130 4765 2169 4767
rect 2203 4765 2242 4767
rect 2276 4765 2315 4767
rect 2349 4765 2388 4767
rect 2422 4765 2461 4767
rect 2495 4765 2534 4767
rect 2568 4765 2607 4767
rect 2641 4767 2666 4799
rect 13782 4851 13838 4869
rect 13782 4835 13840 4851
rect 13942 4835 13944 4851
rect 13782 4812 13944 4835
rect 13782 4801 13838 4812
rect 13782 4767 13816 4801
rect 13872 4778 13910 4812
rect 13850 4767 13944 4778
rect 2641 4765 2680 4767
rect 2714 4765 2753 4767
rect 2787 4765 2826 4767
rect 2860 4765 2899 4767
rect 2933 4765 2972 4767
rect 3006 4765 3045 4767
rect 3079 4765 3118 4767
rect 3152 4765 3191 4767
rect 3225 4765 3264 4767
rect 3298 4765 3337 4767
rect 3371 4765 3410 4767
rect 3444 4765 3483 4767
rect 3517 4765 3556 4767
rect 3590 4765 3629 4767
rect 3663 4765 3702 4767
rect 3736 4765 3775 4767
rect 3809 4765 3848 4767
rect 3882 4765 3921 4767
rect 3955 4765 3994 4767
rect 4028 4765 4067 4767
rect 4101 4765 4140 4767
rect 4174 4765 4213 4767
rect 4247 4765 4286 4767
rect 4320 4765 4359 4767
rect 4393 4765 4432 4767
rect 4466 4765 4505 4767
rect 4539 4765 4578 4767
rect 4612 4765 4651 4767
rect 4685 4765 4724 4767
rect 4758 4765 4797 4767
rect 4831 4765 4870 4767
rect 4904 4765 4943 4767
rect 4977 4765 5016 4767
rect 5050 4765 5089 4767
rect 5123 4765 5162 4767
rect 5196 4765 5235 4767
rect 13765 4765 13944 4767
rect 352 4606 537 4612
rect 352 4572 423 4606
rect 457 4572 537 4606
rect 1178 4602 2130 4603
rect 352 4529 537 4572
rect 352 4495 423 4529
rect 457 4495 537 4529
rect 352 4452 537 4495
rect 1029 4568 1099 4602
rect 1133 4568 1202 4602
rect 1236 4568 2130 4602
rect 995 4534 2130 4568
rect 995 4500 1887 4534
rect 1921 4500 1955 4534
rect 1989 4500 2130 4534
rect 995 4492 2130 4500
rect 1029 4458 1099 4492
rect 1133 4458 1202 4492
rect 1236 4458 2130 4492
rect 352 4418 423 4452
rect 457 4418 537 4452
rect 352 4375 537 4418
rect 352 4341 423 4375
rect 457 4341 537 4375
rect 352 4298 537 4341
rect 352 4264 423 4298
rect 457 4264 537 4298
rect 352 4220 537 4264
rect 352 4186 423 4220
rect 457 4186 537 4220
rect 352 4142 537 4186
rect 352 4108 423 4142
rect 457 4108 537 4142
rect 352 4028 537 4108
rect 352 3984 1877 4028
rect 352 3950 1668 3984
rect 1702 3950 1753 3984
rect 1787 3950 1838 3984
rect 1872 3950 1877 3984
rect 352 3926 1877 3950
rect 13940 3888 14019 3922
rect 48 3806 64 3840
rect 98 3806 599 3840
rect 48 3772 599 3806
rect 13906 3836 14053 3888
rect 13940 3802 14019 3836
rect 48 3738 64 3772
rect 98 3738 599 3772
rect 48 3589 599 3738
rect 14133 3705 14185 3739
rect 48 3555 368 3589
rect 402 3555 467 3589
rect 501 3555 565 3589
rect 48 3517 599 3555
rect 48 3483 368 3517
rect 402 3483 467 3517
rect 501 3483 565 3517
rect 48 3442 599 3483
rect 1669 3664 3331 3670
rect 1669 3646 1749 3664
rect 1783 3646 1822 3664
rect 1856 3646 1895 3664
rect 1929 3646 1968 3664
rect 2002 3646 2041 3664
rect 2075 3646 2113 3664
rect 2147 3646 2185 3664
rect 2219 3646 2257 3664
rect 2291 3646 2329 3664
rect 2363 3646 2401 3664
rect 2435 3646 2473 3664
rect 2507 3646 2545 3664
rect 2579 3646 2617 3664
rect 2651 3646 2689 3664
rect 2723 3646 2761 3664
rect 1669 3612 1677 3646
rect 1711 3612 1747 3646
rect 1783 3630 1817 3646
rect 1856 3630 1887 3646
rect 1929 3630 1957 3646
rect 2002 3630 2027 3646
rect 2075 3630 2097 3646
rect 2147 3630 2167 3646
rect 2219 3630 2237 3646
rect 2291 3630 2307 3646
rect 2363 3630 2377 3646
rect 2435 3630 2447 3646
rect 2507 3630 2517 3646
rect 2579 3630 2587 3646
rect 2651 3630 2657 3646
rect 2723 3630 2727 3646
rect 1781 3612 1817 3630
rect 1851 3612 1887 3630
rect 1921 3612 1957 3630
rect 1991 3612 2027 3630
rect 2061 3612 2097 3630
rect 2131 3612 2167 3630
rect 2201 3612 2237 3630
rect 2271 3612 2307 3630
rect 2341 3612 2377 3630
rect 2411 3612 2447 3630
rect 2481 3612 2517 3630
rect 2551 3612 2587 3630
rect 2621 3612 2657 3630
rect 2691 3612 2727 3630
rect 2795 3646 2833 3664
rect 2795 3630 2797 3646
rect 2761 3612 2797 3630
rect 2831 3630 2833 3646
rect 2867 3646 2905 3664
rect 2939 3646 2977 3664
rect 3011 3646 3049 3664
rect 3083 3646 3121 3664
rect 3155 3646 3193 3664
rect 3227 3646 3265 3664
rect 3299 3646 3331 3664
rect 2831 3612 2867 3630
rect 2901 3630 2905 3646
rect 2971 3630 2977 3646
rect 3041 3630 3049 3646
rect 3111 3630 3121 3646
rect 3181 3630 3193 3646
rect 3251 3630 3265 3646
rect 2901 3612 2937 3630
rect 2971 3612 3007 3630
rect 3041 3612 3077 3630
rect 3111 3612 3147 3630
rect 3181 3612 3217 3630
rect 3251 3612 3287 3630
rect 3321 3612 3331 3646
rect 1669 3592 3331 3612
rect 1669 3544 1677 3592
rect 1711 3578 3331 3592
rect 1711 3544 1747 3578
rect 1781 3556 1817 3578
rect 1851 3556 1887 3578
rect 1921 3556 1957 3578
rect 1991 3556 2027 3578
rect 2061 3556 2097 3578
rect 2131 3556 2167 3578
rect 2201 3556 2237 3578
rect 2271 3556 2307 3578
rect 1781 3544 1785 3556
rect 1851 3544 1859 3556
rect 1921 3544 1933 3556
rect 1991 3544 2007 3556
rect 2061 3544 2081 3556
rect 2131 3544 2155 3556
rect 2201 3544 2229 3556
rect 2271 3544 2303 3556
rect 2341 3544 2377 3578
rect 2411 3544 2447 3578
rect 2481 3556 2517 3578
rect 2551 3556 2587 3578
rect 2621 3556 2657 3578
rect 2691 3556 2727 3578
rect 2761 3556 2797 3578
rect 2831 3556 2867 3578
rect 2901 3556 2937 3578
rect 2971 3556 3007 3578
rect 2485 3544 2517 3556
rect 2559 3544 2587 3556
rect 2633 3544 2657 3556
rect 2707 3544 2727 3556
rect 2781 3544 2797 3556
rect 2855 3544 2867 3556
rect 2929 3544 2937 3556
rect 3003 3544 3007 3556
rect 3041 3556 3077 3578
rect 3041 3544 3043 3556
rect 1669 3522 1785 3544
rect 1819 3522 1859 3544
rect 1893 3522 1933 3544
rect 1967 3522 2007 3544
rect 2041 3522 2081 3544
rect 2115 3522 2155 3544
rect 2189 3522 2229 3544
rect 2263 3522 2303 3544
rect 2337 3522 2377 3544
rect 2411 3522 2451 3544
rect 2485 3522 2525 3544
rect 2559 3522 2599 3544
rect 2633 3522 2673 3544
rect 2707 3522 2747 3544
rect 2781 3522 2821 3544
rect 2855 3522 2895 3544
rect 2929 3522 2969 3544
rect 3003 3522 3043 3544
rect 3111 3556 3147 3578
rect 3181 3556 3217 3578
rect 3251 3556 3287 3578
rect 3111 3544 3117 3556
rect 3181 3544 3191 3556
rect 3251 3544 3265 3556
rect 3321 3544 3331 3578
rect 3077 3522 3117 3544
rect 3151 3522 3191 3544
rect 3225 3522 3265 3544
rect 3299 3522 3331 3544
rect 1669 3520 3331 3522
rect 1669 3476 1677 3520
rect 1711 3510 3331 3520
rect 3400 3664 11240 3670
rect 3400 3630 3432 3664
rect 3466 3630 3505 3664
rect 3539 3630 3578 3664
rect 3612 3630 3651 3664
rect 3685 3630 3724 3664
rect 3758 3630 3797 3664
rect 3831 3630 3870 3664
rect 3904 3630 3942 3664
rect 3976 3630 4014 3664
rect 4048 3630 4086 3664
rect 4120 3630 4158 3664
rect 4192 3630 4230 3664
rect 4264 3630 4302 3664
rect 4336 3630 4374 3664
rect 4408 3630 4446 3664
rect 4480 3630 4518 3664
rect 4552 3630 4590 3664
rect 4624 3630 4662 3664
rect 4696 3630 4734 3664
rect 4768 3630 4806 3664
rect 4840 3630 4878 3664
rect 4912 3630 4950 3664
rect 4984 3630 5022 3664
rect 5056 3630 5094 3664
rect 5128 3630 5166 3664
rect 5200 3630 5238 3664
rect 5272 3630 5310 3664
rect 5344 3630 5382 3664
rect 5416 3630 5454 3664
rect 5488 3630 5526 3664
rect 5560 3630 5598 3664
rect 5632 3630 5670 3664
rect 5704 3630 5742 3664
rect 5776 3630 5814 3664
rect 5848 3630 5886 3664
rect 5920 3630 5958 3664
rect 5992 3630 6030 3664
rect 6064 3630 6102 3664
rect 6136 3630 6174 3664
rect 6208 3630 6246 3664
rect 6280 3630 6318 3664
rect 6352 3630 6390 3664
rect 6424 3630 6462 3664
rect 6496 3630 6534 3664
rect 6568 3630 6606 3664
rect 6640 3630 6678 3664
rect 6712 3630 6750 3664
rect 6784 3630 6822 3664
rect 6856 3630 6894 3664
rect 6928 3630 6966 3664
rect 7000 3630 7038 3664
rect 7072 3630 7110 3664
rect 7144 3630 7182 3664
rect 7216 3630 7428 3664
rect 7462 3630 7501 3664
rect 7535 3630 7574 3664
rect 7608 3630 7646 3664
rect 7680 3630 7718 3664
rect 7752 3630 7790 3664
rect 7824 3630 7862 3664
rect 7896 3630 7934 3664
rect 7968 3630 8006 3664
rect 8040 3630 8078 3664
rect 8112 3630 8150 3664
rect 8184 3630 8222 3664
rect 8256 3630 8294 3664
rect 8328 3630 8366 3664
rect 8400 3630 8438 3664
rect 8472 3630 8510 3664
rect 8544 3630 8582 3664
rect 8616 3630 8654 3664
rect 8688 3630 8726 3664
rect 8760 3630 8798 3664
rect 8832 3630 8870 3664
rect 8904 3630 8942 3664
rect 8976 3630 9014 3664
rect 9048 3630 9086 3664
rect 9120 3630 9158 3664
rect 9192 3630 9230 3664
rect 9264 3630 9302 3664
rect 9336 3630 9374 3664
rect 9408 3630 9446 3664
rect 9480 3630 9518 3664
rect 9552 3630 9590 3664
rect 9624 3630 9662 3664
rect 9696 3630 9734 3664
rect 9768 3630 9806 3664
rect 9840 3630 9878 3664
rect 9912 3630 9950 3664
rect 9984 3630 10022 3664
rect 10056 3630 10094 3664
rect 10128 3630 10166 3664
rect 10200 3630 10238 3664
rect 10272 3630 10310 3664
rect 10344 3630 10382 3664
rect 10416 3630 10454 3664
rect 10488 3630 10526 3664
rect 10560 3630 10598 3664
rect 10632 3630 10670 3664
rect 10704 3630 10742 3664
rect 10776 3630 10814 3664
rect 10848 3630 10886 3664
rect 10920 3630 10958 3664
rect 10992 3630 11030 3664
rect 11064 3630 11102 3664
rect 11136 3630 11174 3664
rect 11208 3630 11240 3664
rect 3400 3556 11240 3630
rect 14099 3626 14219 3705
rect 14133 3592 14185 3626
rect 3400 3522 3432 3556
rect 3466 3522 3505 3556
rect 3539 3522 3578 3556
rect 3612 3522 3651 3556
rect 3685 3522 3724 3556
rect 3758 3522 3797 3556
rect 3831 3522 3870 3556
rect 3904 3522 3942 3556
rect 3976 3522 4014 3556
rect 4048 3522 4086 3556
rect 4120 3522 4158 3556
rect 4192 3522 4230 3556
rect 4264 3522 4302 3556
rect 4336 3522 4374 3556
rect 4408 3522 4446 3556
rect 4480 3522 4518 3556
rect 4552 3522 4590 3556
rect 4624 3522 4662 3556
rect 4696 3522 4734 3556
rect 4768 3522 4806 3556
rect 4840 3522 4878 3556
rect 4912 3522 4950 3556
rect 4984 3522 5022 3556
rect 5056 3522 5094 3556
rect 5128 3522 5166 3556
rect 5200 3522 5238 3556
rect 5272 3522 5310 3556
rect 5344 3522 5382 3556
rect 5416 3522 5454 3556
rect 5488 3522 5526 3556
rect 5560 3522 5598 3556
rect 5632 3522 5670 3556
rect 5704 3522 5742 3556
rect 5776 3522 5814 3556
rect 5848 3522 5886 3556
rect 5920 3522 5958 3556
rect 5992 3522 6030 3556
rect 6064 3522 6102 3556
rect 6136 3522 6174 3556
rect 6208 3522 6246 3556
rect 6280 3522 6318 3556
rect 6352 3522 6390 3556
rect 6424 3522 6462 3556
rect 6496 3522 6534 3556
rect 6568 3522 6606 3556
rect 6640 3522 6678 3556
rect 6712 3522 6750 3556
rect 6784 3522 6822 3556
rect 6856 3522 6894 3556
rect 6928 3522 6966 3556
rect 7000 3522 7038 3556
rect 7072 3522 7110 3556
rect 7144 3522 7182 3556
rect 7216 3522 7428 3556
rect 7462 3522 7501 3556
rect 7535 3522 7574 3556
rect 7608 3522 7646 3556
rect 7680 3522 7718 3556
rect 7752 3522 7790 3556
rect 7824 3522 7862 3556
rect 7896 3522 7934 3556
rect 7968 3522 8006 3556
rect 8040 3522 8078 3556
rect 8112 3522 8150 3556
rect 8184 3522 8222 3556
rect 8256 3522 8294 3556
rect 8328 3522 8366 3556
rect 8400 3522 8438 3556
rect 8472 3522 8510 3556
rect 8544 3522 8582 3556
rect 8616 3522 8654 3556
rect 8688 3522 8726 3556
rect 8760 3522 8798 3556
rect 8832 3522 8870 3556
rect 8904 3522 8942 3556
rect 8976 3522 9014 3556
rect 9048 3522 9086 3556
rect 9120 3522 9158 3556
rect 9192 3522 9230 3556
rect 9264 3522 9302 3556
rect 9336 3522 9374 3556
rect 9408 3522 9446 3556
rect 9480 3522 9518 3556
rect 9552 3522 9590 3556
rect 9624 3522 9662 3556
rect 9696 3522 9734 3556
rect 9768 3522 9806 3556
rect 9840 3522 9878 3556
rect 9912 3522 9950 3556
rect 9984 3522 10022 3556
rect 10056 3522 10094 3556
rect 10128 3522 10166 3556
rect 10200 3522 10238 3556
rect 10272 3522 10310 3556
rect 10344 3522 10382 3556
rect 10416 3522 10454 3556
rect 10488 3522 10526 3556
rect 10560 3522 10598 3556
rect 10632 3522 10670 3556
rect 10704 3522 10742 3556
rect 10776 3522 10814 3556
rect 10848 3522 10886 3556
rect 10920 3522 10958 3556
rect 10992 3522 11030 3556
rect 11064 3522 11102 3556
rect 11136 3522 11174 3556
rect 11208 3522 11240 3556
rect 3400 3516 11240 3522
rect 1711 3476 1747 3510
rect 1781 3484 1817 3510
rect 1781 3476 1785 3484
rect 1851 3476 1887 3510
rect 1921 3476 1957 3510
rect 1991 3476 2027 3510
rect 2061 3476 2097 3510
rect 2131 3476 2167 3510
rect 2201 3476 2237 3510
rect 2271 3476 2307 3510
rect 2341 3476 2377 3510
rect 2411 3476 2447 3510
rect 2481 3476 2517 3510
rect 2551 3476 2587 3510
rect 2621 3476 2657 3510
rect 2691 3476 2727 3510
rect 2761 3476 2797 3510
rect 2831 3476 2867 3510
rect 2901 3476 2937 3510
rect 2971 3476 3007 3510
rect 3041 3476 3077 3510
rect 3111 3476 3147 3510
rect 3181 3476 3217 3510
rect 3251 3476 3287 3510
rect 3321 3476 3331 3510
rect 1669 3450 1785 3476
rect 1819 3461 3331 3476
rect 1819 3450 1892 3461
rect 1669 3448 1892 3450
rect 270 3408 345 3442
rect 402 3408 420 3442
rect 470 3408 494 3442
rect 538 3408 568 3442
rect 606 3408 640 3442
rect 676 3408 708 3442
rect 750 3408 776 3442
rect 825 3408 844 3442
rect 900 3408 912 3442
rect 975 3408 980 3442
rect 1014 3408 1016 3442
rect 1082 3408 1091 3442
rect 1150 3408 1166 3442
rect 1218 3408 1241 3442
rect 1286 3408 1316 3442
rect 1354 3408 1422 3442
rect 270 3374 304 3408
rect 270 3306 304 3336
rect 1388 3370 1422 3408
rect 270 3238 304 3263
rect 270 3170 304 3190
rect 270 3102 304 3117
rect 270 3034 304 3044
rect 270 2966 304 2971
rect 270 2859 304 2864
rect 270 2786 304 2796
rect 270 2713 304 2728
rect 270 2640 304 2660
rect 270 2567 304 2592
rect 270 2494 304 2524
rect 270 2422 304 2456
rect 270 2354 304 2387
rect 270 2286 304 2314
rect 270 2218 304 2242
rect 270 2150 304 2170
rect 270 2082 304 2098
rect 270 2014 304 2026
rect 270 1946 304 1954
rect 369 3248 403 3288
rect 369 3174 403 3214
rect 369 3100 403 3140
rect 553 3248 587 3288
rect 553 3174 587 3214
rect 553 3100 587 3140
rect 369 3026 403 3066
rect 369 2951 403 2992
rect 369 2876 403 2917
rect 369 2801 403 2842
rect 369 2726 403 2767
rect 369 2651 403 2692
rect 369 2576 403 2617
rect 369 2501 403 2542
rect 369 2426 403 2467
rect 369 2351 403 2392
rect 369 2276 403 2317
rect 369 2201 403 2242
rect 369 2126 403 2167
rect 369 2051 403 2092
rect 461 3015 495 3054
rect 461 2942 495 2981
rect 461 2869 495 2908
rect 461 2796 495 2835
rect 461 2723 495 2762
rect 461 2650 495 2689
rect 461 2577 495 2616
rect 461 2504 495 2543
rect 461 2431 495 2470
rect 461 2358 495 2397
rect 461 2284 495 2324
rect 461 2210 495 2250
rect 461 2136 495 2176
rect 461 2062 495 2102
rect 737 3248 771 3288
rect 737 3174 771 3214
rect 737 3100 771 3140
rect 553 3026 587 3066
rect 553 2951 587 2992
rect 553 2876 587 2917
rect 553 2801 587 2842
rect 553 2726 587 2767
rect 553 2651 587 2692
rect 553 2576 587 2617
rect 553 2501 587 2542
rect 553 2426 587 2467
rect 553 2351 587 2392
rect 553 2276 587 2317
rect 553 2201 587 2242
rect 553 2126 587 2167
rect 553 2051 587 2092
rect 369 1976 403 2017
rect 645 3015 679 3054
rect 645 2942 679 2981
rect 645 2869 679 2908
rect 645 2796 679 2835
rect 645 2723 679 2762
rect 645 2650 679 2689
rect 645 2577 679 2616
rect 645 2504 679 2543
rect 645 2431 679 2470
rect 645 2358 679 2397
rect 645 2284 679 2324
rect 645 2210 679 2250
rect 645 2136 679 2176
rect 645 2062 679 2102
rect 921 3248 955 3288
rect 921 3174 955 3214
rect 921 3100 955 3140
rect 737 3026 771 3066
rect 737 2951 771 2992
rect 737 2876 771 2917
rect 737 2801 771 2842
rect 737 2726 771 2767
rect 737 2651 771 2692
rect 737 2576 771 2617
rect 737 2501 771 2542
rect 737 2426 771 2467
rect 737 2351 771 2392
rect 737 2276 771 2317
rect 737 2201 771 2242
rect 737 2126 771 2167
rect 737 2051 771 2092
rect 553 1976 587 2017
rect 829 3015 863 3054
rect 829 2942 863 2981
rect 829 2869 863 2908
rect 829 2796 863 2835
rect 829 2723 863 2762
rect 829 2650 863 2689
rect 829 2577 863 2616
rect 829 2504 863 2543
rect 829 2431 863 2470
rect 829 2358 863 2397
rect 829 2284 863 2324
rect 829 2210 863 2250
rect 829 2136 863 2176
rect 829 2062 863 2102
rect 1105 3248 1139 3288
rect 1105 3174 1139 3214
rect 1105 3100 1139 3140
rect 921 3026 955 3066
rect 921 2951 955 2992
rect 921 2876 955 2917
rect 921 2801 955 2842
rect 921 2726 955 2767
rect 921 2651 955 2692
rect 921 2576 955 2617
rect 921 2501 955 2542
rect 921 2426 955 2467
rect 921 2351 955 2392
rect 921 2276 955 2317
rect 921 2201 955 2242
rect 921 2126 955 2167
rect 921 2051 955 2092
rect 737 1976 771 2017
rect 1013 3015 1047 3054
rect 1013 2942 1047 2981
rect 1013 2869 1047 2908
rect 1013 2796 1047 2835
rect 1013 2723 1047 2762
rect 1013 2650 1047 2689
rect 1013 2577 1047 2616
rect 1013 2504 1047 2543
rect 1013 2431 1047 2470
rect 1013 2358 1047 2397
rect 1013 2284 1047 2324
rect 1013 2210 1047 2250
rect 1013 2136 1047 2176
rect 1013 2062 1047 2102
rect 1289 3248 1323 3288
rect 1289 3174 1323 3214
rect 1289 3100 1323 3140
rect 1105 3026 1139 3066
rect 1105 2951 1139 2992
rect 1105 2876 1139 2917
rect 1105 2801 1139 2842
rect 1105 2726 1139 2767
rect 1105 2651 1139 2692
rect 1105 2576 1139 2617
rect 1105 2501 1139 2542
rect 1105 2426 1139 2467
rect 1105 2351 1139 2392
rect 1105 2276 1139 2317
rect 1105 2201 1139 2242
rect 1105 2126 1139 2167
rect 1105 2051 1139 2092
rect 921 1976 955 2017
rect 1197 3015 1231 3054
rect 1197 2942 1231 2981
rect 1197 2869 1231 2908
rect 1197 2796 1231 2835
rect 1197 2723 1231 2762
rect 1197 2650 1231 2689
rect 1197 2577 1231 2616
rect 1197 2504 1231 2543
rect 1197 2431 1231 2470
rect 1197 2358 1231 2397
rect 1197 2284 1231 2324
rect 1197 2210 1231 2250
rect 1197 2136 1231 2176
rect 1197 2062 1231 2102
rect 1289 3026 1323 3066
rect 1289 2951 1323 2992
rect 1289 2876 1323 2917
rect 1289 2801 1323 2842
rect 1289 2726 1323 2767
rect 1289 2651 1323 2692
rect 1289 2576 1323 2617
rect 1289 2501 1323 2542
rect 1289 2426 1323 2467
rect 1289 2351 1323 2392
rect 1289 2276 1323 2317
rect 1289 2201 1323 2242
rect 1289 2126 1323 2167
rect 1289 2051 1323 2092
rect 1105 1976 1139 2017
rect 1289 1976 1323 2017
rect 1388 3298 1422 3332
rect 1388 3230 1422 3264
rect 1388 3162 1422 3192
rect 1388 3094 1422 3120
rect 1388 3026 1422 3048
rect 1388 2958 1422 2976
rect 1388 2890 1422 2904
rect 1388 2822 1422 2832
rect 1388 2754 1422 2760
rect 1388 2686 1422 2688
rect 1388 2650 1422 2652
rect 1388 2578 1422 2584
rect 1388 2506 1422 2516
rect 1388 2434 1422 2448
rect 1388 2362 1422 2380
rect 1388 2290 1422 2312
rect 1388 2218 1422 2244
rect 1388 2146 1422 2176
rect 1388 2074 1422 2108
rect 1388 2006 1422 2040
rect 1388 1938 1422 1968
rect 270 1878 304 1882
rect 414 1852 430 1886
rect 464 1852 503 1886
rect 537 1852 576 1886
rect 610 1852 649 1886
rect 683 1852 722 1886
rect 756 1852 795 1886
rect 829 1852 868 1886
rect 902 1852 940 1886
rect 974 1852 1012 1886
rect 1046 1852 1084 1886
rect 1118 1852 1156 1886
rect 1190 1852 1228 1886
rect 1262 1852 1278 1886
rect 1388 1870 1422 1896
rect 1388 1802 1422 1824
rect 270 1772 304 1776
rect 270 1700 304 1708
rect 270 1628 304 1640
rect 270 1556 304 1572
rect 270 1484 304 1504
rect 270 1412 304 1436
rect 270 1340 304 1368
rect 270 1268 304 1300
rect 270 1198 304 1232
rect 270 1130 304 1162
rect 270 1062 304 1090
rect 270 994 304 1018
rect 270 926 304 946
rect 270 858 304 874
rect 270 790 304 824
rect 270 722 304 756
rect 270 654 304 688
rect 369 1718 403 1758
rect 369 1644 403 1684
rect 369 1570 403 1610
rect 369 1496 403 1536
rect 369 1422 403 1462
rect 369 1348 403 1388
rect 369 1274 403 1314
rect 369 1200 403 1240
rect 369 1126 403 1166
rect 369 1052 403 1092
rect 369 978 403 1018
rect 369 903 403 944
rect 369 828 403 869
rect 369 753 403 794
rect 369 678 403 719
rect 461 1718 495 1758
rect 461 1644 495 1684
rect 461 1570 495 1610
rect 461 1496 495 1536
rect 461 1422 495 1462
rect 461 1348 495 1388
rect 461 1274 495 1314
rect 461 1200 495 1240
rect 461 1126 495 1166
rect 461 1052 495 1092
rect 461 978 495 1018
rect 461 904 495 944
rect 461 830 495 870
rect 461 756 495 796
rect 461 682 495 722
rect 270 586 304 620
rect 270 518 304 552
rect 461 607 495 648
rect 553 1718 587 1758
rect 553 1644 587 1684
rect 553 1570 587 1610
rect 553 1496 587 1536
rect 553 1422 587 1462
rect 553 1348 587 1388
rect 553 1274 587 1314
rect 553 1200 587 1240
rect 553 1126 587 1166
rect 553 1052 587 1092
rect 553 978 587 1018
rect 553 903 587 944
rect 553 828 587 869
rect 553 753 587 794
rect 553 678 587 719
rect 645 1718 679 1758
rect 645 1644 679 1684
rect 645 1570 679 1610
rect 645 1496 679 1536
rect 645 1422 679 1462
rect 645 1348 679 1388
rect 645 1274 679 1314
rect 645 1200 679 1240
rect 645 1126 679 1166
rect 645 1052 679 1092
rect 645 978 679 1018
rect 645 904 679 944
rect 645 830 679 870
rect 645 756 679 796
rect 645 682 679 722
rect 461 532 495 573
rect 645 607 679 648
rect 737 1718 771 1758
rect 737 1644 771 1684
rect 737 1570 771 1610
rect 737 1496 771 1536
rect 737 1422 771 1462
rect 737 1348 771 1388
rect 737 1274 771 1314
rect 737 1200 771 1240
rect 737 1126 771 1166
rect 737 1052 771 1092
rect 737 978 771 1018
rect 737 903 771 944
rect 737 828 771 869
rect 737 753 771 794
rect 737 678 771 719
rect 829 1718 863 1758
rect 829 1644 863 1684
rect 829 1570 863 1610
rect 829 1496 863 1536
rect 829 1422 863 1462
rect 829 1348 863 1388
rect 829 1274 863 1314
rect 829 1200 863 1240
rect 829 1126 863 1166
rect 829 1052 863 1092
rect 829 978 863 1018
rect 829 904 863 944
rect 829 830 863 870
rect 829 756 863 796
rect 829 682 863 722
rect 645 532 679 573
rect 829 607 863 648
rect 921 1718 955 1758
rect 921 1644 955 1684
rect 921 1570 955 1610
rect 921 1496 955 1536
rect 921 1422 955 1462
rect 921 1348 955 1388
rect 921 1274 955 1314
rect 921 1200 955 1240
rect 921 1126 955 1166
rect 921 1052 955 1092
rect 921 978 955 1018
rect 921 903 955 944
rect 921 828 955 869
rect 921 753 955 794
rect 921 678 955 719
rect 1013 1718 1047 1758
rect 1013 1644 1047 1684
rect 1013 1570 1047 1610
rect 1013 1496 1047 1536
rect 1013 1422 1047 1462
rect 1013 1348 1047 1388
rect 1013 1274 1047 1314
rect 1013 1200 1047 1240
rect 1013 1126 1047 1166
rect 1013 1052 1047 1092
rect 1013 978 1047 1018
rect 1013 904 1047 944
rect 1013 830 1047 870
rect 1013 756 1047 796
rect 1013 682 1047 722
rect 829 532 863 573
rect 1013 607 1047 648
rect 1105 1718 1139 1758
rect 1105 1644 1139 1684
rect 1105 1570 1139 1610
rect 1105 1496 1139 1536
rect 1105 1422 1139 1462
rect 1105 1348 1139 1388
rect 1105 1274 1139 1314
rect 1105 1200 1139 1240
rect 1105 1126 1139 1166
rect 1105 1052 1139 1092
rect 1105 978 1139 1018
rect 1105 903 1139 944
rect 1105 828 1139 869
rect 1105 753 1139 794
rect 1105 678 1139 719
rect 1197 1718 1231 1758
rect 1197 1644 1231 1684
rect 1197 1570 1231 1610
rect 1197 1496 1231 1536
rect 1197 1422 1231 1462
rect 1197 1348 1231 1388
rect 1197 1274 1231 1314
rect 1197 1200 1231 1240
rect 1197 1126 1231 1166
rect 1197 1052 1231 1092
rect 1197 978 1231 1018
rect 1197 904 1231 944
rect 1197 830 1231 870
rect 1197 756 1231 796
rect 1197 682 1231 722
rect 1013 532 1047 573
rect 1197 607 1231 648
rect 1197 532 1231 573
rect 1289 1718 1323 1758
rect 1289 1644 1323 1684
rect 1289 1570 1323 1610
rect 1289 1496 1323 1536
rect 1289 1421 1323 1462
rect 1289 1346 1323 1387
rect 1289 1271 1323 1312
rect 1289 1196 1323 1237
rect 1289 1121 1323 1162
rect 1289 1046 1323 1087
rect 1289 971 1323 1012
rect 1289 896 1323 937
rect 1289 821 1323 862
rect 1289 746 1323 787
rect 1289 671 1323 712
rect 1289 596 1323 637
rect 1289 521 1323 562
rect 270 450 304 484
rect 270 382 304 416
rect 1289 446 1323 487
rect 1388 1734 1422 1751
rect 1388 1666 1422 1678
rect 1388 1598 1422 1605
rect 1388 1530 1422 1532
rect 1388 1493 1422 1496
rect 1388 1420 1422 1428
rect 1388 1347 1422 1360
rect 1388 1274 1422 1292
rect 1388 1201 1422 1224
rect 1388 1128 1422 1156
rect 1388 1055 1422 1088
rect 1388 986 1422 1020
rect 1388 918 1422 948
rect 1388 850 1422 875
rect 1388 782 1422 802
rect 1388 714 1422 729
rect 1388 646 1422 656
rect 1388 578 1422 612
rect 1388 510 1422 544
rect 1388 442 1422 476
rect 1388 374 1422 408
rect 270 238 304 348
rect 414 322 426 356
rect 464 322 500 356
rect 537 322 574 356
rect 610 322 648 356
rect 683 322 721 356
rect 756 322 794 356
rect 829 322 867 356
rect 902 322 940 356
rect 974 322 1012 356
rect 1047 322 1084 356
rect 1120 322 1156 356
rect 1193 322 1228 356
rect 1266 322 1278 356
rect 1388 306 1422 340
rect 1669 3408 1677 3448
rect 1711 3442 1892 3448
rect 1926 3442 1967 3461
rect 2001 3442 2042 3461
rect 2076 3442 2117 3461
rect 2151 3442 2192 3461
rect 2226 3442 2266 3461
rect 2300 3442 2340 3461
rect 2374 3442 2414 3461
rect 2448 3442 2488 3461
rect 2522 3442 2562 3461
rect 2596 3442 2636 3461
rect 2670 3442 2710 3461
rect 2744 3442 2784 3461
rect 2818 3442 2858 3461
rect 2892 3442 2932 3461
rect 2966 3442 3006 3461
rect 3040 3442 3080 3461
rect 3114 3442 3154 3461
rect 3188 3442 3228 3461
rect 3262 3442 3331 3461
rect 1711 3408 1747 3442
rect 1781 3412 1817 3442
rect 1781 3408 1785 3412
rect 1851 3408 1887 3442
rect 1926 3427 1957 3442
rect 2001 3427 2027 3442
rect 2076 3427 2097 3442
rect 2151 3427 2167 3442
rect 2226 3427 2237 3442
rect 2300 3427 2307 3442
rect 2374 3427 2377 3442
rect 1921 3408 1957 3427
rect 1991 3408 2027 3427
rect 2061 3408 2097 3427
rect 2131 3408 2167 3427
rect 2201 3408 2237 3427
rect 2271 3408 2307 3427
rect 2341 3408 2377 3427
rect 2411 3427 2414 3442
rect 2481 3427 2488 3442
rect 2551 3427 2562 3442
rect 2621 3427 2636 3442
rect 2691 3427 2710 3442
rect 2761 3427 2784 3442
rect 2831 3427 2858 3442
rect 2901 3427 2932 3442
rect 2971 3427 3006 3442
rect 2411 3408 2447 3427
rect 2481 3408 2517 3427
rect 2551 3408 2587 3427
rect 2621 3408 2657 3427
rect 2691 3408 2727 3427
rect 2761 3408 2797 3427
rect 2831 3408 2867 3427
rect 2901 3408 2937 3427
rect 2971 3408 3007 3427
rect 3041 3408 3077 3442
rect 3114 3427 3147 3442
rect 3188 3427 3217 3442
rect 3262 3427 3287 3442
rect 3111 3408 3147 3427
rect 3181 3408 3217 3427
rect 3251 3408 3287 3427
rect 3321 3408 3331 3442
rect 1669 3378 1785 3408
rect 1819 3389 3331 3408
rect 1819 3378 1892 3389
rect 1669 3376 1892 3378
rect 1669 3340 1677 3376
rect 1711 3374 1892 3376
rect 1926 3374 1967 3389
rect 2001 3374 2042 3389
rect 2076 3374 2117 3389
rect 2151 3374 2192 3389
rect 2226 3374 2266 3389
rect 2300 3374 2340 3389
rect 2374 3374 2414 3389
rect 2448 3374 2488 3389
rect 2522 3374 2562 3389
rect 2596 3374 2636 3389
rect 2670 3374 2710 3389
rect 2744 3374 2784 3389
rect 2818 3374 2858 3389
rect 2892 3374 2932 3389
rect 2966 3374 3006 3389
rect 3040 3374 3080 3389
rect 3114 3374 3154 3389
rect 3188 3374 3228 3389
rect 3262 3374 3331 3389
rect 13523 3420 13621 3454
rect 13657 3420 13689 3454
rect 13723 3420 13747 3454
rect 13791 3420 13821 3454
rect 13859 3420 13893 3454
rect 13929 3420 13961 3454
rect 14003 3420 14029 3454
rect 14078 3420 14097 3454
rect 14153 3420 14165 3454
rect 14228 3420 14233 3454
rect 14267 3420 14269 3454
rect 14335 3420 14344 3454
rect 14403 3420 14419 3454
rect 14471 3420 14494 3454
rect 14539 3420 14569 3454
rect 14607 3420 14675 3454
rect 13523 3386 13557 3420
rect 1711 3340 1747 3374
rect 1781 3340 1817 3374
rect 1851 3340 1887 3374
rect 1926 3355 1957 3374
rect 2001 3355 2027 3374
rect 2076 3355 2097 3374
rect 2151 3355 2167 3374
rect 2226 3355 2237 3374
rect 2300 3355 2307 3374
rect 2374 3355 2377 3374
rect 1921 3340 1957 3355
rect 1991 3340 2027 3355
rect 2061 3340 2097 3355
rect 2131 3340 2167 3355
rect 2201 3340 2237 3355
rect 2271 3340 2307 3355
rect 2341 3340 2377 3355
rect 2411 3355 2414 3374
rect 2481 3355 2488 3374
rect 2551 3355 2562 3374
rect 2621 3355 2636 3374
rect 2691 3355 2710 3374
rect 2761 3355 2784 3374
rect 2831 3355 2858 3374
rect 2901 3355 2932 3374
rect 2971 3355 3006 3374
rect 2411 3340 2447 3355
rect 2481 3340 2517 3355
rect 2551 3340 2587 3355
rect 2621 3340 2657 3355
rect 2691 3340 2727 3355
rect 2761 3340 2797 3355
rect 2831 3340 2867 3355
rect 2901 3340 2937 3355
rect 2971 3340 3007 3355
rect 3041 3340 3077 3374
rect 3114 3355 3147 3374
rect 3188 3355 3217 3374
rect 3262 3355 3287 3374
rect 3111 3340 3147 3355
rect 3181 3340 3217 3355
rect 3251 3340 3287 3355
rect 3321 3340 3331 3374
rect 1669 3306 1785 3340
rect 1819 3317 3331 3340
rect 1819 3306 1892 3317
rect 1926 3306 1967 3317
rect 2001 3306 2042 3317
rect 2076 3306 2117 3317
rect 2151 3306 2192 3317
rect 2226 3306 2266 3317
rect 2300 3306 2340 3317
rect 2374 3306 2414 3317
rect 2448 3306 2488 3317
rect 2522 3306 2562 3317
rect 2596 3306 2636 3317
rect 2670 3306 2710 3317
rect 2744 3306 2784 3317
rect 2818 3306 2858 3317
rect 2892 3306 2932 3317
rect 2966 3306 3006 3317
rect 3040 3306 3080 3317
rect 3114 3306 3154 3317
rect 3188 3306 3228 3317
rect 3262 3306 3331 3317
rect 1669 3270 1677 3306
rect 1711 3272 1747 3306
rect 1781 3272 1817 3306
rect 1851 3272 1887 3306
rect 1926 3283 1957 3306
rect 2001 3283 2027 3306
rect 2076 3283 2097 3306
rect 2151 3283 2167 3306
rect 2226 3283 2237 3306
rect 2300 3283 2307 3306
rect 2374 3283 2377 3306
rect 1921 3272 1957 3283
rect 1991 3272 2027 3283
rect 2061 3272 2097 3283
rect 2131 3272 2167 3283
rect 2201 3272 2237 3283
rect 2271 3272 2307 3283
rect 2341 3272 2377 3283
rect 2411 3283 2414 3306
rect 2481 3283 2488 3306
rect 2551 3283 2562 3306
rect 2621 3283 2636 3306
rect 2691 3283 2710 3306
rect 2761 3283 2784 3306
rect 2831 3283 2858 3306
rect 2901 3283 2932 3306
rect 2971 3283 3006 3306
rect 2411 3272 2447 3283
rect 2481 3272 2517 3283
rect 2551 3272 2587 3283
rect 2621 3272 2657 3283
rect 2691 3272 2727 3283
rect 2761 3272 2797 3283
rect 2831 3272 2867 3283
rect 2901 3272 2937 3283
rect 2971 3272 3007 3283
rect 3041 3272 3077 3306
rect 3114 3283 3147 3306
rect 3188 3283 3217 3306
rect 3262 3283 3287 3306
rect 3111 3272 3147 3283
rect 3181 3272 3217 3283
rect 3251 3272 3287 3283
rect 3321 3272 3331 3306
rect 13523 3318 13557 3348
rect 14641 3382 14675 3420
rect 1711 3270 3331 3272
rect 1669 3268 3331 3270
rect 1669 3238 1785 3268
rect 1819 3245 3331 3268
rect 1819 3238 1892 3245
rect 1926 3238 1967 3245
rect 2001 3238 2042 3245
rect 2076 3238 2117 3245
rect 2151 3238 2192 3245
rect 2226 3238 2266 3245
rect 2300 3238 2340 3245
rect 2374 3238 2414 3245
rect 2448 3238 2488 3245
rect 2522 3238 2562 3245
rect 2596 3238 2636 3245
rect 2670 3238 2710 3245
rect 2744 3238 2784 3245
rect 2818 3238 2858 3245
rect 2892 3238 2932 3245
rect 2966 3238 3006 3245
rect 3040 3238 3080 3245
rect 3114 3238 3154 3245
rect 3188 3238 3228 3245
rect 3262 3238 3331 3245
rect 1669 3198 1677 3238
rect 1711 3204 1747 3238
rect 1781 3234 1785 3238
rect 1781 3204 1817 3234
rect 1851 3204 1887 3238
rect 1926 3211 1957 3238
rect 2001 3211 2027 3238
rect 2076 3211 2097 3238
rect 2151 3211 2167 3238
rect 2226 3211 2237 3238
rect 2300 3211 2307 3238
rect 2374 3211 2377 3238
rect 1921 3204 1957 3211
rect 1991 3204 2027 3211
rect 2061 3204 2097 3211
rect 2131 3204 2167 3211
rect 2201 3204 2237 3211
rect 2271 3204 2307 3211
rect 2341 3204 2377 3211
rect 2411 3211 2414 3238
rect 2481 3211 2488 3238
rect 2551 3211 2562 3238
rect 2621 3211 2636 3238
rect 2691 3211 2710 3238
rect 2761 3211 2784 3238
rect 2831 3211 2858 3238
rect 2901 3211 2932 3238
rect 2971 3211 3006 3238
rect 2411 3204 2447 3211
rect 2481 3204 2517 3211
rect 2551 3204 2587 3211
rect 2621 3204 2657 3211
rect 2691 3204 2727 3211
rect 2761 3204 2797 3211
rect 2831 3204 2867 3211
rect 2901 3204 2937 3211
rect 2971 3204 3007 3211
rect 3041 3204 3077 3238
rect 3114 3211 3147 3238
rect 3188 3211 3217 3238
rect 3262 3211 3287 3238
rect 3111 3204 3147 3211
rect 3181 3204 3217 3211
rect 3251 3204 3287 3211
rect 3321 3204 3331 3238
rect 1711 3198 3331 3204
rect 1669 3196 3331 3198
rect 1669 3169 1785 3196
rect 1819 3173 3331 3196
rect 1819 3169 1892 3173
rect 1926 3169 1967 3173
rect 2001 3169 2042 3173
rect 2076 3169 2117 3173
rect 2151 3169 2192 3173
rect 2226 3169 2266 3173
rect 2300 3169 2340 3173
rect 2374 3169 2414 3173
rect 2448 3169 2488 3173
rect 2522 3169 2562 3173
rect 2596 3169 2636 3173
rect 2670 3169 2710 3173
rect 2744 3169 2784 3173
rect 2818 3169 2858 3173
rect 2892 3169 2932 3173
rect 2966 3169 3006 3173
rect 3040 3169 3080 3173
rect 3114 3169 3154 3173
rect 3188 3169 3228 3173
rect 3262 3169 3331 3173
rect 1669 3126 1677 3169
rect 1711 3135 1747 3169
rect 1781 3162 1785 3169
rect 1781 3135 1817 3162
rect 1851 3135 1887 3169
rect 1926 3139 1957 3169
rect 2001 3139 2027 3169
rect 2076 3139 2097 3169
rect 2151 3139 2167 3169
rect 2226 3139 2237 3169
rect 2300 3139 2307 3169
rect 2374 3139 2377 3169
rect 1921 3135 1957 3139
rect 1991 3135 2027 3139
rect 2061 3135 2097 3139
rect 2131 3135 2167 3139
rect 2201 3135 2237 3139
rect 2271 3135 2307 3139
rect 2341 3135 2377 3139
rect 2411 3139 2414 3169
rect 2481 3139 2488 3169
rect 2551 3139 2562 3169
rect 2621 3139 2636 3169
rect 2691 3139 2710 3169
rect 2761 3139 2784 3169
rect 2831 3139 2858 3169
rect 2901 3139 2932 3169
rect 2971 3139 3006 3169
rect 2411 3135 2447 3139
rect 2481 3135 2517 3139
rect 2551 3135 2587 3139
rect 2621 3135 2657 3139
rect 2691 3135 2727 3139
rect 2761 3135 2797 3139
rect 2831 3135 2867 3139
rect 2901 3135 2937 3139
rect 2971 3135 3007 3139
rect 3041 3135 3077 3169
rect 3114 3139 3147 3169
rect 3188 3139 3217 3169
rect 3262 3139 3287 3169
rect 3111 3135 3147 3139
rect 3181 3135 3217 3139
rect 3251 3135 3287 3139
rect 3321 3135 3331 3169
rect 1711 3126 3331 3135
rect 1669 3124 3331 3126
rect 1669 3100 1785 3124
rect 1819 3100 3331 3124
rect 1669 3054 1677 3100
rect 1711 3066 1747 3100
rect 1781 3090 1785 3100
rect 1781 3066 1817 3090
rect 1851 3066 1887 3100
rect 1921 3066 1957 3100
rect 1991 3066 2027 3100
rect 2061 3066 2097 3100
rect 2131 3066 2167 3100
rect 2201 3066 2237 3100
rect 2271 3066 2307 3100
rect 2341 3066 2377 3100
rect 2411 3066 2447 3100
rect 2481 3066 2517 3100
rect 2551 3066 2587 3100
rect 2621 3066 2657 3100
rect 2691 3066 2727 3100
rect 2761 3066 2797 3100
rect 2831 3066 2867 3100
rect 2901 3066 2937 3100
rect 2971 3066 3007 3100
rect 3041 3066 3077 3100
rect 3111 3066 3147 3100
rect 3181 3066 3217 3100
rect 3251 3066 3287 3100
rect 3321 3066 3331 3100
rect 1711 3054 3331 3066
rect 1669 3052 3331 3054
rect 1669 3031 1785 3052
rect 1819 3031 3331 3052
rect 1669 2982 1677 3031
rect 1711 2997 1747 3031
rect 1781 3018 1785 3031
rect 1781 2997 1817 3018
rect 1851 2997 1887 3031
rect 1921 2997 1957 3031
rect 1991 2997 2027 3031
rect 2061 2997 2097 3031
rect 2131 2997 2167 3031
rect 2201 2997 2237 3031
rect 2271 2997 2307 3031
rect 2341 2997 2377 3031
rect 2411 2997 2447 3031
rect 2481 2997 2517 3031
rect 2551 2997 2587 3031
rect 2621 2997 2657 3031
rect 2691 2997 2727 3031
rect 2761 2997 2797 3031
rect 2831 2997 2867 3031
rect 2901 2997 2937 3031
rect 2971 2997 3007 3031
rect 3041 2997 3077 3031
rect 3111 2997 3147 3031
rect 3181 2997 3217 3031
rect 3251 2997 3287 3031
rect 3321 2997 3331 3031
rect 1711 2982 3331 2997
rect 1669 2980 3331 2982
rect 1669 2962 1785 2980
rect 1819 2962 3331 2980
rect 1669 2910 1677 2962
rect 1711 2928 1747 2962
rect 1781 2946 1785 2962
rect 1781 2928 1817 2946
rect 1851 2928 1887 2962
rect 1921 2928 1957 2962
rect 1991 2928 2027 2962
rect 2061 2928 2097 2962
rect 2131 2928 2167 2962
rect 2201 2928 2237 2962
rect 2271 2928 2307 2962
rect 2341 2928 2377 2962
rect 2411 2928 2447 2962
rect 2481 2928 2517 2962
rect 2551 2928 2587 2962
rect 2621 2928 2657 2962
rect 2691 2928 2727 2962
rect 2761 2928 2797 2962
rect 2831 2928 2867 2962
rect 2901 2928 2937 2962
rect 2971 2928 3007 2962
rect 3041 2928 3077 2962
rect 3111 2928 3147 2962
rect 3181 2928 3217 2962
rect 3251 2928 3287 2962
rect 3321 2928 3331 2962
rect 1711 2910 3331 2928
rect 1669 2908 3331 2910
rect 1669 2893 1785 2908
rect 1819 2893 3331 2908
rect 1669 2838 1677 2893
rect 1711 2859 1747 2893
rect 1781 2874 1785 2893
rect 1781 2859 1817 2874
rect 1851 2859 1887 2893
rect 1921 2859 1957 2893
rect 1991 2859 2027 2893
rect 2061 2859 2097 2893
rect 2131 2859 2167 2893
rect 2201 2859 2237 2893
rect 2271 2859 2307 2893
rect 2341 2859 2377 2893
rect 2411 2859 2447 2893
rect 2481 2859 2517 2893
rect 2551 2859 2587 2893
rect 2621 2859 2657 2893
rect 2691 2859 2727 2893
rect 2761 2859 2797 2893
rect 2831 2859 2867 2893
rect 2901 2859 2937 2893
rect 2971 2859 3007 2893
rect 3041 2859 3077 2893
rect 3111 2859 3147 2893
rect 3181 2859 3217 2893
rect 3251 2859 3287 2893
rect 3321 2859 3331 2893
rect 1711 2838 3331 2859
rect 1669 2836 3331 2838
rect 1669 2824 1785 2836
rect 1819 2824 3331 2836
rect 1669 2766 1677 2824
rect 1711 2790 1747 2824
rect 1781 2802 1785 2824
rect 1781 2790 1817 2802
rect 1851 2790 1887 2824
rect 1921 2790 1957 2824
rect 1991 2790 2027 2824
rect 2061 2790 2097 2824
rect 2131 2790 2167 2824
rect 2201 2790 2237 2824
rect 2271 2790 2307 2824
rect 2341 2790 2377 2824
rect 2411 2790 2447 2824
rect 2481 2790 2517 2824
rect 2551 2790 2587 2824
rect 2621 2790 2657 2824
rect 2691 2790 2727 2824
rect 2761 2790 2797 2824
rect 2831 2790 2867 2824
rect 2901 2790 2937 2824
rect 2971 2790 3007 2824
rect 3041 2790 3077 2824
rect 3111 2790 3147 2824
rect 3181 2790 3217 2824
rect 3251 2790 3287 2824
rect 3321 2790 3331 2824
rect 1711 2766 3331 2790
rect 1669 2764 3331 2766
rect 1669 2755 1785 2764
rect 1819 2755 3331 2764
rect 1669 2694 1677 2755
rect 1711 2721 1747 2755
rect 1781 2730 1785 2755
rect 1781 2721 1817 2730
rect 1851 2721 1887 2755
rect 1921 2721 1957 2755
rect 1991 2721 2027 2755
rect 2061 2721 2097 2755
rect 2131 2721 2167 2755
rect 2201 2721 2237 2755
rect 2271 2721 2307 2755
rect 2341 2721 2377 2755
rect 2411 2721 2447 2755
rect 2481 2721 2517 2755
rect 2551 2721 2587 2755
rect 2621 2721 2657 2755
rect 2691 2721 2727 2755
rect 2761 2721 2797 2755
rect 2831 2721 2867 2755
rect 2901 2721 2937 2755
rect 2971 2721 3007 2755
rect 3041 2721 3077 2755
rect 3111 2721 3147 2755
rect 3181 2721 3217 2755
rect 3251 2721 3287 2755
rect 3321 2721 3331 2755
rect 1711 2694 3331 2721
rect 1669 2692 3331 2694
rect 1669 2686 1785 2692
rect 1819 2686 3331 2692
rect 1669 2622 1677 2686
rect 1711 2652 1747 2686
rect 1781 2658 1785 2686
rect 1781 2652 1817 2658
rect 1851 2652 1887 2686
rect 1921 2652 1957 2686
rect 1991 2652 2027 2686
rect 2061 2652 2097 2686
rect 2131 2652 2167 2686
rect 2201 2652 2237 2686
rect 2271 2652 2307 2686
rect 2341 2652 2377 2686
rect 2411 2652 2447 2686
rect 2481 2652 2517 2686
rect 2551 2652 2587 2686
rect 2621 2652 2657 2686
rect 2691 2652 2727 2686
rect 2761 2652 2797 2686
rect 2831 2652 2867 2686
rect 2901 2652 2937 2686
rect 2971 2652 3007 2686
rect 3041 2652 3077 2686
rect 3111 2652 3147 2686
rect 3181 2652 3217 2686
rect 3251 2652 3287 2686
rect 3321 2652 3331 2686
rect 1711 2622 3331 2652
rect 1669 2620 3331 2622
rect 1669 2617 1785 2620
rect 1819 2617 3331 2620
rect 1669 2550 1677 2617
rect 1711 2583 1747 2617
rect 1781 2586 1785 2617
rect 1781 2583 1817 2586
rect 1851 2583 1887 2617
rect 1921 2583 1957 2617
rect 1991 2583 2027 2617
rect 2061 2583 2097 2617
rect 2131 2583 2167 2617
rect 2201 2583 2237 2617
rect 2271 2583 2307 2617
rect 2341 2583 2377 2617
rect 2411 2583 2447 2617
rect 2481 2583 2517 2617
rect 2551 2583 2587 2617
rect 2621 2583 2657 2617
rect 2691 2583 2727 2617
rect 2761 2583 2797 2617
rect 2831 2583 2867 2617
rect 2901 2583 2937 2617
rect 2971 2583 3007 2617
rect 3041 2583 3077 2617
rect 3111 2583 3147 2617
rect 3181 2583 3217 2617
rect 3251 2583 3287 2617
rect 3321 2583 3331 2617
rect 1711 2550 3331 2583
rect 1669 2548 3331 2550
rect 1669 2514 1677 2548
rect 1711 2514 1747 2548
rect 1781 2547 1817 2548
rect 1781 2514 1785 2547
rect 1851 2514 1887 2548
rect 1921 2514 1957 2548
rect 1991 2514 2027 2548
rect 2061 2514 2097 2548
rect 2131 2514 2167 2548
rect 2201 2514 2237 2548
rect 2271 2514 2307 2548
rect 2341 2514 2377 2548
rect 2411 2514 2447 2548
rect 2481 2514 2517 2548
rect 2551 2514 2587 2548
rect 2621 2514 2657 2548
rect 2691 2514 2727 2548
rect 2761 2514 2797 2548
rect 2831 2514 2867 2548
rect 2901 2514 2937 2548
rect 2971 2514 3007 2548
rect 3041 2514 3077 2548
rect 3111 2514 3147 2548
rect 3181 2514 3217 2548
rect 3251 2514 3287 2548
rect 3321 2514 3331 2548
rect 1669 2513 1785 2514
rect 1819 2513 3331 2514
rect 1669 2511 3331 2513
rect 1669 2445 1677 2511
rect 1711 2479 3331 2511
rect 1711 2445 1747 2479
rect 1781 2474 1817 2479
rect 1781 2445 1785 2474
rect 1851 2445 1887 2479
rect 1921 2445 1957 2479
rect 1991 2445 2027 2479
rect 2061 2445 2097 2479
rect 2131 2445 2167 2479
rect 2201 2445 2237 2479
rect 2271 2445 2307 2479
rect 2341 2445 2377 2479
rect 2411 2445 2447 2479
rect 2481 2445 2517 2479
rect 2551 2445 2587 2479
rect 2621 2445 2657 2479
rect 2691 2445 2727 2479
rect 2761 2445 2797 2479
rect 2831 2445 2867 2479
rect 2901 2445 2937 2479
rect 2971 2445 3007 2479
rect 3041 2445 3077 2479
rect 3111 2445 3147 2479
rect 3181 2445 3217 2479
rect 3251 2445 3287 2479
rect 3321 2445 3331 2479
rect 1669 2440 1785 2445
rect 1819 2440 3331 2445
rect 1669 2438 3331 2440
rect 1669 2376 1677 2438
rect 1711 2410 3331 2438
rect 1711 2376 1747 2410
rect 1781 2401 1817 2410
rect 1781 2376 1785 2401
rect 1851 2376 1887 2410
rect 1921 2376 1957 2410
rect 1991 2376 2027 2410
rect 2061 2376 2097 2410
rect 2131 2376 2167 2410
rect 2201 2376 2237 2410
rect 2271 2376 2307 2410
rect 2341 2376 2377 2410
rect 2411 2376 2447 2410
rect 2481 2376 2517 2410
rect 2551 2376 2587 2410
rect 2621 2376 2657 2410
rect 2691 2376 2727 2410
rect 2761 2376 2797 2410
rect 2831 2376 2867 2410
rect 2901 2376 2937 2410
rect 2971 2376 3007 2410
rect 3041 2376 3077 2410
rect 3111 2376 3147 2410
rect 3181 2376 3217 2410
rect 3251 2376 3287 2410
rect 3321 2376 3331 2410
rect 1669 2367 1785 2376
rect 1819 2367 3331 2376
rect 1669 2365 3331 2367
rect 1669 2307 1677 2365
rect 1711 2341 3331 2365
rect 1711 2307 1747 2341
rect 1781 2328 1817 2341
rect 1781 2307 1785 2328
rect 1851 2307 1887 2341
rect 1921 2307 1957 2341
rect 1991 2307 2027 2341
rect 2061 2307 2097 2341
rect 2131 2307 2167 2341
rect 2201 2307 2237 2341
rect 2271 2307 2307 2341
rect 2341 2307 2377 2341
rect 2411 2307 2447 2341
rect 2481 2307 2517 2341
rect 2551 2307 2587 2341
rect 2621 2307 2657 2341
rect 2691 2307 2727 2341
rect 2761 2307 2797 2341
rect 2831 2307 2867 2341
rect 2901 2307 2937 2341
rect 2971 2307 3007 2341
rect 3041 2307 3077 2341
rect 3111 2307 3147 2341
rect 3181 2307 3217 2341
rect 3251 2307 3287 2341
rect 3321 2307 3331 2341
rect 1669 2294 1785 2307
rect 1819 2294 3331 2307
rect 1669 2292 3331 2294
rect 1669 2238 1677 2292
rect 1711 2272 3331 2292
rect 1711 2238 1747 2272
rect 1781 2255 1817 2272
rect 1781 2238 1785 2255
rect 1851 2238 1887 2272
rect 1921 2238 1957 2272
rect 1991 2238 2027 2272
rect 2061 2238 2097 2272
rect 2131 2238 2167 2272
rect 2201 2238 2237 2272
rect 2271 2238 2307 2272
rect 2341 2238 2377 2272
rect 2411 2238 2447 2272
rect 2481 2238 2517 2272
rect 2551 2238 2587 2272
rect 2621 2238 2657 2272
rect 2691 2238 2727 2272
rect 2761 2238 2797 2272
rect 2831 2238 2867 2272
rect 2901 2238 2937 2272
rect 2971 2238 3007 2272
rect 3041 2238 3077 2272
rect 3111 2238 3147 2272
rect 3181 2238 3217 2272
rect 3251 2238 3287 2272
rect 3321 2238 3331 2272
rect 1669 2221 1785 2238
rect 1819 2221 3331 2238
rect 1669 2219 3331 2221
rect 1669 2169 1677 2219
rect 1711 2203 3331 2219
rect 1711 2169 1747 2203
rect 1781 2182 1817 2203
rect 1781 2169 1785 2182
rect 1851 2169 1887 2203
rect 1921 2169 1957 2203
rect 1991 2169 2027 2203
rect 2061 2169 2097 2203
rect 2131 2169 2167 2203
rect 2201 2169 2237 2203
rect 2271 2169 2307 2203
rect 2341 2169 2377 2203
rect 2411 2169 2447 2203
rect 2481 2169 2517 2203
rect 2551 2169 2587 2203
rect 2621 2169 2657 2203
rect 2691 2169 2727 2203
rect 2761 2169 2797 2203
rect 2831 2169 2867 2203
rect 2901 2169 2937 2203
rect 2971 2169 3007 2203
rect 3041 2169 3077 2203
rect 3111 2169 3147 2203
rect 3181 2169 3217 2203
rect 3251 2169 3287 2203
rect 3321 2169 3331 2203
rect 1669 2148 1785 2169
rect 1819 2148 3331 2169
rect 1669 2146 3331 2148
rect 1669 2100 1677 2146
rect 1711 2134 3331 2146
rect 1711 2100 1747 2134
rect 1781 2109 1817 2134
rect 1781 2100 1785 2109
rect 1851 2100 1887 2134
rect 1921 2100 1957 2134
rect 1991 2100 2027 2134
rect 2061 2100 2097 2134
rect 2131 2100 2167 2134
rect 2201 2100 2237 2134
rect 2271 2100 2307 2134
rect 2341 2100 2377 2134
rect 2411 2100 2447 2134
rect 2481 2100 2517 2134
rect 2551 2100 2587 2134
rect 2621 2100 2657 2134
rect 2691 2100 2727 2134
rect 2761 2100 2797 2134
rect 2831 2100 2867 2134
rect 2901 2100 2937 2134
rect 2971 2100 3007 2134
rect 3041 2100 3077 2134
rect 3111 2100 3147 2134
rect 3181 2100 3217 2134
rect 3251 2100 3287 2134
rect 3321 2100 3331 2134
rect 1669 2075 1785 2100
rect 1819 2075 3331 2100
rect 1669 2073 3331 2075
rect 1669 2031 1677 2073
rect 1711 2065 3331 2073
rect 1711 2031 1747 2065
rect 1781 2036 1817 2065
rect 1781 2031 1785 2036
rect 1851 2031 1887 2065
rect 1921 2031 1957 2065
rect 1991 2031 2027 2065
rect 2061 2031 2097 2065
rect 2131 2031 2167 2065
rect 2201 2031 2237 2065
rect 2271 2031 2307 2065
rect 2341 2031 2377 2065
rect 2411 2031 2447 2065
rect 2481 2031 2517 2065
rect 2551 2031 2587 2065
rect 2621 2031 2657 2065
rect 2691 2031 2727 2065
rect 2761 2031 2797 2065
rect 2831 2031 2867 2065
rect 2901 2031 2937 2065
rect 2971 2031 3007 2065
rect 3041 2031 3077 2065
rect 3111 2031 3147 2065
rect 3181 2031 3217 2065
rect 3251 2031 3287 2065
rect 3321 2031 3331 2065
rect 1669 2002 1785 2031
rect 1819 2002 3331 2031
rect 1669 2000 3331 2002
rect 1669 1962 1677 2000
rect 1711 1996 3331 2000
rect 1711 1962 1747 1996
rect 1781 1963 1817 1996
rect 1781 1962 1785 1963
rect 1851 1962 1887 1996
rect 1921 1962 1957 1996
rect 1991 1962 2027 1996
rect 2061 1962 2097 1996
rect 2131 1962 2167 1996
rect 2201 1962 2237 1996
rect 2271 1962 2307 1996
rect 2341 1962 2377 1996
rect 2411 1962 2447 1996
rect 2481 1962 2517 1996
rect 2551 1962 2587 1996
rect 2621 1962 2657 1996
rect 2691 1962 2727 1996
rect 2761 1962 2797 1996
rect 2831 1962 2867 1996
rect 2901 1962 2937 1996
rect 2971 1962 3007 1996
rect 3041 1962 3077 1996
rect 3111 1962 3147 1996
rect 3181 1962 3217 1996
rect 3251 1962 3287 1996
rect 3321 1962 3331 1996
rect 1669 1929 1785 1962
rect 1819 1929 3331 1962
rect 1669 1927 3331 1929
rect 1669 1893 1677 1927
rect 1711 1893 1747 1927
rect 1781 1893 1817 1927
rect 1851 1893 1887 1927
rect 1921 1893 1957 1927
rect 1991 1893 2027 1927
rect 2061 1893 2097 1927
rect 2131 1893 2167 1927
rect 2201 1893 2237 1927
rect 2271 1893 2307 1927
rect 2341 1893 2377 1927
rect 2411 1893 2447 1927
rect 2481 1893 2517 1927
rect 2551 1893 2587 1927
rect 2621 1893 2657 1927
rect 2691 1893 2727 1927
rect 2761 1893 2797 1927
rect 2831 1893 2867 1927
rect 2901 1893 2937 1927
rect 2971 1893 3007 1927
rect 3041 1893 3077 1927
rect 3111 1893 3147 1927
rect 3181 1893 3217 1927
rect 3251 1893 3287 1927
rect 3321 1893 3331 1927
rect 1669 1890 3331 1893
rect 1669 1858 1785 1890
rect 1819 1858 3331 1890
rect 1669 1820 1677 1858
rect 1711 1824 1747 1858
rect 1781 1856 1785 1858
rect 1781 1824 1817 1856
rect 1851 1824 1887 1858
rect 1921 1824 1957 1858
rect 1991 1824 2027 1858
rect 2061 1824 2097 1858
rect 2131 1824 2167 1858
rect 2201 1824 2237 1858
rect 2271 1824 2307 1858
rect 2341 1824 2377 1858
rect 2411 1824 2447 1858
rect 2481 1824 2517 1858
rect 2551 1824 2587 1858
rect 2621 1824 2657 1858
rect 2691 1824 2727 1858
rect 2761 1824 2797 1858
rect 2831 1824 2867 1858
rect 2901 1824 2937 1858
rect 2971 1824 3007 1858
rect 3041 1824 3077 1858
rect 3111 1824 3147 1858
rect 3181 1824 3217 1858
rect 3251 1824 3287 1858
rect 3321 1824 3331 1858
rect 1711 1820 3331 1824
rect 1669 1817 3331 1820
rect 1669 1789 1785 1817
rect 1819 1789 3331 1817
rect 1669 1747 1677 1789
rect 1711 1755 1747 1789
rect 1781 1783 1785 1789
rect 1781 1755 1817 1783
rect 1851 1755 1887 1789
rect 1921 1755 1957 1789
rect 1991 1755 2027 1789
rect 2061 1755 2097 1789
rect 2131 1755 2167 1789
rect 2201 1755 2237 1789
rect 2271 1755 2307 1789
rect 2341 1755 2377 1789
rect 2411 1755 2447 1789
rect 2481 1755 2517 1789
rect 2551 1755 2587 1789
rect 2621 1755 2657 1789
rect 2691 1755 2727 1789
rect 2761 1755 2797 1789
rect 2831 1755 2867 1789
rect 2901 1755 2937 1789
rect 2971 1755 3007 1789
rect 3041 1755 3077 1789
rect 3111 1755 3147 1789
rect 3181 1755 3217 1789
rect 3251 1755 3287 1789
rect 3321 1755 3331 1789
rect 1711 1747 3331 1755
rect 1669 1744 3331 1747
rect 1669 1720 1785 1744
rect 1819 1720 3331 1744
rect 1669 1674 1677 1720
rect 1711 1686 1747 1720
rect 1781 1710 1785 1720
rect 1781 1686 1817 1710
rect 1851 1686 1887 1720
rect 1921 1686 1957 1720
rect 1991 1686 2027 1720
rect 2061 1686 2097 1720
rect 2131 1686 2167 1720
rect 2201 1686 2237 1720
rect 2271 1686 2307 1720
rect 2341 1686 2377 1720
rect 2411 1686 2447 1720
rect 2481 1686 2517 1720
rect 2551 1686 2587 1720
rect 2621 1686 2657 1720
rect 2691 1686 2727 1720
rect 2761 1686 2797 1720
rect 2831 1686 2867 1720
rect 2901 1686 2937 1720
rect 2971 1686 3007 1720
rect 3041 1686 3077 1720
rect 3111 1686 3147 1720
rect 3181 1686 3217 1720
rect 3251 1686 3287 1720
rect 3321 1686 3331 1720
rect 1711 1674 3331 1686
rect 1669 1671 3331 1674
rect 1669 1651 1785 1671
rect 1819 1651 3331 1671
rect 1669 1601 1677 1651
rect 1711 1617 1747 1651
rect 1781 1637 1785 1651
rect 1781 1617 1817 1637
rect 1851 1617 1887 1651
rect 1921 1617 1957 1651
rect 1991 1617 2027 1651
rect 2061 1617 2097 1651
rect 2131 1617 2167 1651
rect 2201 1617 2237 1651
rect 2271 1617 2307 1651
rect 2341 1617 2377 1651
rect 2411 1617 2447 1651
rect 2481 1617 2517 1651
rect 2551 1617 2587 1651
rect 2621 1617 2657 1651
rect 2691 1617 2727 1651
rect 2761 1617 2797 1651
rect 2831 1617 2867 1651
rect 2901 1617 2937 1651
rect 2971 1617 3007 1651
rect 3041 1617 3077 1651
rect 3111 1617 3147 1651
rect 3181 1617 3217 1651
rect 3251 1617 3287 1651
rect 3321 1617 3331 1651
rect 1711 1601 3331 1617
rect 1669 1598 3331 1601
rect 1669 1582 1785 1598
rect 1819 1582 3331 1598
rect 1669 1528 1677 1582
rect 1711 1548 1747 1582
rect 1781 1564 1785 1582
rect 1781 1548 1817 1564
rect 1851 1548 1887 1582
rect 1921 1548 1957 1582
rect 1991 1548 2027 1582
rect 2061 1548 2097 1582
rect 2131 1548 2167 1582
rect 2201 1548 2237 1582
rect 2271 1548 2307 1582
rect 2341 1548 2377 1582
rect 2411 1548 2447 1582
rect 2481 1548 2517 1582
rect 2551 1548 2587 1582
rect 2621 1548 2657 1582
rect 2691 1548 2727 1582
rect 2761 1548 2797 1582
rect 2831 1548 2867 1582
rect 2901 1548 2937 1582
rect 2971 1548 3007 1582
rect 3041 1548 3077 1582
rect 3111 1548 3147 1582
rect 3181 1548 3217 1582
rect 3251 1548 3287 1582
rect 3321 1548 3331 1582
rect 1711 1528 3331 1548
rect 1669 1525 3331 1528
rect 1669 1513 1785 1525
rect 1819 1513 3331 1525
rect 1669 1455 1677 1513
rect 1711 1479 1747 1513
rect 1781 1491 1785 1513
rect 1781 1479 1817 1491
rect 1851 1479 1887 1513
rect 1921 1479 1957 1513
rect 1991 1479 2027 1513
rect 2061 1479 2097 1513
rect 2131 1479 2167 1513
rect 2201 1479 2237 1513
rect 2271 1479 2307 1513
rect 2341 1479 2377 1513
rect 2411 1479 2447 1513
rect 2481 1479 2517 1513
rect 2551 1479 2587 1513
rect 2621 1479 2657 1513
rect 2691 1479 2727 1513
rect 2761 1479 2797 1513
rect 2831 1479 2867 1513
rect 2901 1479 2937 1513
rect 2971 1479 3007 1513
rect 3041 1479 3077 1513
rect 3111 1479 3147 1513
rect 3181 1479 3217 1513
rect 3251 1479 3287 1513
rect 3321 1479 3331 1513
rect 1711 1455 3331 1479
rect 1669 1452 3331 1455
rect 1669 1444 1785 1452
rect 1819 1444 3331 1452
rect 1669 1382 1677 1444
rect 1711 1410 1747 1444
rect 1781 1418 1785 1444
rect 1781 1410 1817 1418
rect 1851 1410 1887 1444
rect 1921 1410 1957 1444
rect 1991 1410 2027 1444
rect 2061 1410 2097 1444
rect 2131 1410 2167 1444
rect 2201 1410 2237 1444
rect 2271 1410 2307 1444
rect 2341 1410 2377 1444
rect 2411 1410 2447 1444
rect 2481 1410 2517 1444
rect 2551 1410 2587 1444
rect 2621 1410 2657 1444
rect 2691 1410 2727 1444
rect 2761 1410 2797 1444
rect 2831 1410 2867 1444
rect 2901 1410 2937 1444
rect 2971 1410 3007 1444
rect 3041 1410 3077 1444
rect 3111 1410 3147 1444
rect 3181 1410 3217 1444
rect 3251 1410 3287 1444
rect 3321 1410 3331 1444
rect 1711 1382 3331 1410
rect 1669 1379 3331 1382
rect 1669 1375 1785 1379
rect 1819 1375 3331 1379
rect 1669 1309 1677 1375
rect 1711 1341 1747 1375
rect 1781 1345 1785 1375
rect 1781 1341 1817 1345
rect 1851 1341 1887 1375
rect 1921 1341 1957 1375
rect 1991 1341 2027 1375
rect 2061 1341 2097 1375
rect 2131 1341 2167 1375
rect 2201 1341 2237 1375
rect 2271 1341 2307 1375
rect 2341 1341 2377 1375
rect 2411 1341 2447 1375
rect 2481 1341 2517 1375
rect 2551 1341 2587 1375
rect 2621 1341 2657 1375
rect 2691 1341 2727 1375
rect 2761 1341 2797 1375
rect 2831 1341 2867 1375
rect 2901 1341 2937 1375
rect 2971 1341 3007 1375
rect 3041 1341 3077 1375
rect 3111 1341 3147 1375
rect 3181 1341 3217 1375
rect 3251 1341 3287 1375
rect 3321 1341 3331 1375
rect 1711 1309 3331 1341
rect 1669 1306 3331 1309
rect 1669 1272 1677 1306
rect 1711 1272 1747 1306
rect 1781 1272 1785 1306
rect 1851 1272 1887 1306
rect 1921 1272 1957 1306
rect 1991 1272 2027 1306
rect 2061 1272 2097 1306
rect 2131 1272 2167 1306
rect 2201 1272 2237 1306
rect 2271 1272 2307 1306
rect 2341 1272 2377 1306
rect 2411 1272 2447 1306
rect 2481 1272 2517 1306
rect 2551 1272 2587 1306
rect 2621 1272 2657 1306
rect 2691 1272 2727 1306
rect 2761 1272 2797 1306
rect 2831 1272 2867 1306
rect 2901 1272 2937 1306
rect 2971 1272 3007 1306
rect 3041 1272 3077 1306
rect 3111 1272 3147 1306
rect 3181 1272 3217 1306
rect 3251 1272 3287 1306
rect 3321 1272 3331 1306
rect 1669 1270 3331 1272
rect 1669 1203 1677 1270
rect 1711 1237 3331 1270
rect 1711 1203 1747 1237
rect 1781 1233 1817 1237
rect 1781 1203 1785 1233
rect 1851 1203 1887 1237
rect 1921 1203 1957 1237
rect 1991 1203 2027 1237
rect 2061 1203 2097 1237
rect 2131 1203 2167 1237
rect 2201 1203 2237 1237
rect 2271 1203 2307 1237
rect 2341 1203 2377 1237
rect 2411 1203 2447 1237
rect 2481 1203 2517 1237
rect 2551 1203 2587 1237
rect 2621 1203 2657 1237
rect 2691 1203 2727 1237
rect 2761 1203 2797 1237
rect 2831 1203 2867 1237
rect 2901 1203 2937 1237
rect 2971 1203 3007 1237
rect 3041 1203 3077 1237
rect 3111 1203 3147 1237
rect 3181 1203 3217 1237
rect 3251 1203 3287 1237
rect 3321 1203 3331 1237
rect 1669 1199 1785 1203
rect 1819 1199 3331 1203
rect 1669 1197 3331 1199
rect 1669 1134 1677 1197
rect 1711 1168 3331 1197
rect 1711 1134 1747 1168
rect 1781 1160 1817 1168
rect 1781 1134 1785 1160
rect 1851 1134 1887 1168
rect 1921 1134 1957 1168
rect 1991 1134 2027 1168
rect 2061 1134 2097 1168
rect 2131 1134 2167 1168
rect 2201 1134 2237 1168
rect 2271 1134 2307 1168
rect 2341 1134 2377 1168
rect 2411 1134 2447 1168
rect 2481 1134 2517 1168
rect 2551 1134 2587 1168
rect 2621 1134 2657 1168
rect 2691 1134 2727 1168
rect 2761 1134 2797 1168
rect 2831 1134 2867 1168
rect 2901 1134 2937 1168
rect 2971 1134 3007 1168
rect 3041 1134 3077 1168
rect 3111 1134 3147 1168
rect 3181 1134 3217 1168
rect 3251 1134 3287 1168
rect 3321 1134 3331 1168
rect 1669 1126 1785 1134
rect 1819 1126 3331 1134
rect 1669 1124 3331 1126
rect 1669 1065 1677 1124
rect 1711 1099 3331 1124
rect 1711 1065 1747 1099
rect 1781 1087 1817 1099
rect 1781 1065 1785 1087
rect 1851 1065 1887 1099
rect 1921 1065 1957 1099
rect 1991 1065 2027 1099
rect 2061 1065 2097 1099
rect 2131 1065 2167 1099
rect 2201 1065 2237 1099
rect 2271 1065 2307 1099
rect 2341 1065 2377 1099
rect 2411 1065 2447 1099
rect 2481 1065 2517 1099
rect 2551 1065 2587 1099
rect 2621 1065 2657 1099
rect 2691 1065 2727 1099
rect 2761 1065 2797 1099
rect 2831 1065 2867 1099
rect 2901 1065 2937 1099
rect 2971 1065 3007 1099
rect 3041 1065 3077 1099
rect 3111 1065 3147 1099
rect 3181 1065 3217 1099
rect 3251 1065 3287 1099
rect 3321 1065 3331 1099
rect 1669 1053 1785 1065
rect 1819 1053 3331 1065
rect 1669 1051 3331 1053
rect 1669 996 1677 1051
rect 1711 1030 3331 1051
rect 1711 996 1747 1030
rect 1781 1014 1817 1030
rect 1781 996 1785 1014
rect 1851 996 1887 1030
rect 1921 996 1957 1030
rect 1991 996 2027 1030
rect 2061 996 2097 1030
rect 2131 996 2167 1030
rect 2201 996 2237 1030
rect 2271 996 2307 1030
rect 2341 996 2377 1030
rect 2411 996 2447 1030
rect 2481 996 2517 1030
rect 2551 996 2587 1030
rect 2621 996 2657 1030
rect 2691 996 2727 1030
rect 2761 996 2797 1030
rect 2831 996 2867 1030
rect 2901 996 2937 1030
rect 2971 996 3007 1030
rect 3041 996 3077 1030
rect 3111 996 3147 1030
rect 3181 996 3217 1030
rect 3251 996 3287 1030
rect 3321 996 3331 1030
rect 1669 980 1785 996
rect 1819 980 3331 996
rect 1669 978 3331 980
rect 1669 927 1677 978
rect 1711 961 3331 978
rect 1711 927 1747 961
rect 1781 941 1817 961
rect 1781 927 1785 941
rect 1851 927 1887 961
rect 1921 927 1957 961
rect 1991 927 2027 961
rect 2061 927 2097 961
rect 2131 927 2167 961
rect 2201 927 2237 961
rect 2271 927 2307 961
rect 2341 927 2377 961
rect 2411 927 2447 961
rect 2481 927 2517 961
rect 2551 927 2587 961
rect 2621 927 2657 961
rect 2691 927 2727 961
rect 2761 927 2797 961
rect 2831 927 2867 961
rect 2901 927 2937 961
rect 2971 927 3007 961
rect 3041 927 3077 961
rect 3111 927 3147 961
rect 3181 927 3217 961
rect 3251 927 3287 961
rect 3321 927 3331 961
rect 1669 907 1785 927
rect 1819 907 3331 927
rect 1669 905 3331 907
rect 1669 858 1677 905
rect 1711 892 3331 905
rect 1711 858 1747 892
rect 1781 868 1817 892
rect 1781 858 1785 868
rect 1851 858 1887 892
rect 1921 858 1957 892
rect 1991 858 2027 892
rect 2061 858 2097 892
rect 2131 858 2167 892
rect 2201 858 2237 892
rect 2271 858 2307 892
rect 2341 858 2377 892
rect 2411 858 2447 892
rect 2481 858 2517 892
rect 2551 858 2587 892
rect 2621 858 2657 892
rect 2691 858 2727 892
rect 2761 858 2797 892
rect 2831 858 2867 892
rect 2901 858 2937 892
rect 2971 858 3007 892
rect 3041 858 3077 892
rect 3111 858 3147 892
rect 3181 858 3217 892
rect 3251 858 3287 892
rect 3321 858 3331 892
rect 1669 834 1785 858
rect 1819 834 3331 858
rect 1669 832 3331 834
rect 1669 789 1677 832
rect 1711 823 3331 832
rect 1711 789 1747 823
rect 1781 795 1817 823
rect 1781 789 1785 795
rect 1851 789 1887 823
rect 1921 789 1957 823
rect 1991 789 2027 823
rect 2061 789 2097 823
rect 2131 789 2167 823
rect 2201 789 2237 823
rect 2271 789 2307 823
rect 2341 789 2377 823
rect 2411 789 2447 823
rect 2481 789 2517 823
rect 2551 789 2587 823
rect 2621 789 2657 823
rect 2691 789 2727 823
rect 2761 789 2797 823
rect 2831 789 2867 823
rect 2901 789 2937 823
rect 2971 789 3007 823
rect 3041 789 3077 823
rect 3111 789 3147 823
rect 3181 789 3217 823
rect 3251 789 3287 823
rect 3321 789 3331 823
rect 1669 761 1785 789
rect 1819 761 3331 789
rect 1669 759 3331 761
rect 1669 720 1677 759
rect 1711 754 3331 759
rect 1711 720 1747 754
rect 1781 722 1817 754
rect 1781 720 1785 722
rect 1851 720 1887 754
rect 1921 720 1957 754
rect 1991 720 2027 754
rect 2061 720 2097 754
rect 2131 720 2167 754
rect 2201 720 2237 754
rect 2271 720 2307 754
rect 2341 720 2377 754
rect 2411 720 2447 754
rect 2481 720 2517 754
rect 2551 720 2587 754
rect 2621 720 2657 754
rect 2691 720 2727 754
rect 2761 720 2797 754
rect 2831 720 2867 754
rect 2901 720 2937 754
rect 2971 720 3007 754
rect 3041 720 3077 754
rect 3111 720 3147 754
rect 3181 720 3217 754
rect 3251 720 3287 754
rect 3321 720 3331 754
rect 1669 688 1785 720
rect 1819 688 3331 720
rect 1669 686 3331 688
rect 1669 651 1677 686
rect 1711 685 3331 686
rect 1711 651 1747 685
rect 1781 651 1817 685
rect 1851 651 1887 685
rect 1921 651 1957 685
rect 1991 651 2027 685
rect 2061 651 2097 685
rect 2131 651 2167 685
rect 2201 651 2237 685
rect 2271 651 2307 685
rect 2341 651 2377 685
rect 2411 651 2447 685
rect 2481 651 2517 685
rect 2551 651 2587 685
rect 2621 651 2657 685
rect 2691 651 2727 685
rect 2761 651 2797 685
rect 2831 651 2867 685
rect 2901 651 2937 685
rect 2971 651 3007 685
rect 3041 651 3077 685
rect 3111 651 3147 685
rect 3181 651 3217 685
rect 3251 651 3287 685
rect 3321 651 3331 685
rect 1669 649 3331 651
rect 1669 616 1785 649
rect 1819 616 3331 649
rect 1669 579 1677 616
rect 1711 582 1747 616
rect 1781 615 1785 616
rect 1781 582 1817 615
rect 1851 582 1887 616
rect 1921 582 1957 616
rect 1991 582 2027 616
rect 2061 582 2097 616
rect 2131 582 2167 616
rect 2201 582 2237 616
rect 2271 582 2307 616
rect 2341 582 2377 616
rect 2411 582 2447 616
rect 2481 582 2517 616
rect 2551 582 2587 616
rect 2621 582 2657 616
rect 2691 582 2727 616
rect 2761 582 2797 616
rect 2831 582 2867 616
rect 2901 582 2937 616
rect 2971 582 3007 616
rect 3041 582 3077 616
rect 3111 582 3147 616
rect 3181 582 3217 616
rect 3251 582 3287 616
rect 3321 582 3331 616
rect 1711 579 1892 582
rect 1669 576 1892 579
rect 1669 547 1785 576
rect 1819 548 1892 576
rect 1926 548 1967 582
rect 2001 548 2042 582
rect 2076 548 2117 582
rect 2151 548 2192 582
rect 2226 548 2266 582
rect 2300 548 2340 582
rect 2374 548 2414 582
rect 2448 548 2488 582
rect 2522 548 2562 582
rect 2596 548 2636 582
rect 2670 548 2710 582
rect 2744 548 2784 582
rect 2818 548 2858 582
rect 2892 548 2932 582
rect 2966 548 3006 582
rect 3040 548 3080 582
rect 3114 548 3154 582
rect 3188 548 3228 582
rect 3262 548 3331 582
rect 1819 547 3331 548
rect 1669 506 1677 547
rect 1711 513 1747 547
rect 1781 542 1785 547
rect 1781 513 1817 542
rect 1851 513 1887 547
rect 1921 513 1957 547
rect 1991 513 2027 547
rect 2061 513 2097 547
rect 2131 513 2167 547
rect 2201 513 2237 547
rect 2271 513 2307 547
rect 2341 513 2377 547
rect 2411 513 2447 547
rect 2481 513 2517 547
rect 2551 513 2587 547
rect 2621 513 2657 547
rect 2691 513 2727 547
rect 2761 513 2797 547
rect 2831 513 2867 547
rect 2901 513 2937 547
rect 2971 513 3007 547
rect 3041 513 3077 547
rect 3111 513 3147 547
rect 3181 513 3217 547
rect 3251 513 3287 547
rect 3321 513 3331 547
rect 1711 510 3331 513
rect 1711 506 1892 510
rect 1669 503 1892 506
rect 1669 478 1785 503
rect 1819 478 1892 503
rect 1926 478 1967 510
rect 2001 478 2042 510
rect 2076 478 2117 510
rect 2151 478 2192 510
rect 2226 478 2266 510
rect 2300 478 2340 510
rect 2374 478 2414 510
rect 2448 478 2488 510
rect 2522 478 2562 510
rect 2596 478 2636 510
rect 2670 478 2710 510
rect 2744 478 2784 510
rect 2818 478 2858 510
rect 2892 478 2932 510
rect 2966 478 3006 510
rect 3040 478 3080 510
rect 3114 478 3154 510
rect 3188 478 3228 510
rect 3262 478 3331 510
rect 1669 433 1677 478
rect 1711 444 1747 478
rect 1781 469 1785 478
rect 1781 444 1817 469
rect 1851 444 1887 478
rect 1926 476 1957 478
rect 2001 476 2027 478
rect 2076 476 2097 478
rect 2151 476 2167 478
rect 2226 476 2237 478
rect 2300 476 2307 478
rect 2374 476 2377 478
rect 1921 444 1957 476
rect 1991 444 2027 476
rect 2061 444 2097 476
rect 2131 444 2167 476
rect 2201 444 2237 476
rect 2271 444 2307 476
rect 2341 444 2377 476
rect 2411 476 2414 478
rect 2481 476 2488 478
rect 2551 476 2562 478
rect 2621 476 2636 478
rect 2691 476 2710 478
rect 2761 476 2784 478
rect 2831 476 2858 478
rect 2901 476 2932 478
rect 2971 476 3006 478
rect 2411 444 2447 476
rect 2481 444 2517 476
rect 2551 444 2587 476
rect 2621 444 2657 476
rect 2691 444 2727 476
rect 2761 444 2797 476
rect 2831 444 2867 476
rect 2901 444 2937 476
rect 2971 444 3007 476
rect 3041 444 3077 478
rect 3114 476 3147 478
rect 3188 476 3217 478
rect 3262 476 3287 478
rect 3111 444 3147 476
rect 3181 444 3217 476
rect 3251 444 3287 476
rect 3321 444 3331 478
rect 1711 433 3331 444
rect 1669 430 3331 433
rect 1669 409 1785 430
rect 1819 409 1860 430
rect 1894 409 1935 430
rect 1969 409 2010 430
rect 2044 409 2085 430
rect 2119 409 2160 430
rect 2194 409 2235 430
rect 2269 409 2310 430
rect 2344 409 2385 430
rect 2419 409 2460 430
rect 2494 409 2535 430
rect 2569 409 2610 430
rect 2644 409 2685 430
rect 2719 409 2760 430
rect 2794 409 2835 430
rect 2869 409 2910 430
rect 2944 409 2985 430
rect 3019 409 3060 430
rect 3094 409 3135 430
rect 3169 409 3210 430
rect 3244 409 3331 430
rect 1669 360 1677 409
rect 1711 375 1747 409
rect 1781 396 1785 409
rect 1851 396 1860 409
rect 1921 396 1935 409
rect 1991 396 2010 409
rect 2061 396 2085 409
rect 2131 396 2160 409
rect 2201 396 2235 409
rect 1781 375 1817 396
rect 1851 375 1887 396
rect 1921 375 1957 396
rect 1991 375 2027 396
rect 2061 375 2097 396
rect 2131 375 2167 396
rect 2201 375 2237 396
rect 2271 375 2307 409
rect 2344 396 2377 409
rect 2419 396 2447 409
rect 2494 396 2517 409
rect 2569 396 2587 409
rect 2644 396 2657 409
rect 2719 396 2727 409
rect 2794 396 2797 409
rect 2341 375 2377 396
rect 2411 375 2447 396
rect 2481 375 2517 396
rect 2551 375 2587 396
rect 2621 375 2657 396
rect 2691 375 2727 396
rect 2761 375 2797 396
rect 2831 396 2835 409
rect 2901 396 2910 409
rect 2971 396 2985 409
rect 3041 396 3060 409
rect 3111 396 3135 409
rect 3181 396 3210 409
rect 2831 375 2867 396
rect 2901 375 2937 396
rect 2971 375 3007 396
rect 3041 375 3077 396
rect 3111 375 3147 396
rect 3181 375 3217 396
rect 3251 375 3287 409
rect 3321 375 3331 409
rect 1711 360 3331 375
rect 1669 340 3331 360
rect 13523 3250 13557 3275
rect 13523 3182 13557 3202
rect 13523 3114 13557 3129
rect 13523 3046 13557 3056
rect 13523 2978 13557 2983
rect 13523 2871 13557 2876
rect 13523 2798 13557 2808
rect 13523 2725 13557 2740
rect 13523 2652 13557 2672
rect 13523 2579 13557 2604
rect 13523 2506 13557 2536
rect 13523 2434 13557 2468
rect 13523 2366 13557 2399
rect 13523 2298 13557 2326
rect 13523 2230 13557 2253
rect 13523 2162 13557 2180
rect 13523 2094 13557 2107
rect 13523 2026 13557 2034
rect 13523 1958 13557 1961
rect 13622 3260 13656 3300
rect 13622 3186 13656 3226
rect 13622 3112 13656 3152
rect 13806 3260 13840 3300
rect 13806 3186 13840 3226
rect 13622 3038 13656 3078
rect 13622 2963 13656 3004
rect 13622 2888 13656 2929
rect 13622 2813 13656 2854
rect 13622 2738 13656 2779
rect 13622 2663 13656 2704
rect 13622 2588 13656 2629
rect 13622 2513 13656 2554
rect 13622 2438 13656 2479
rect 13622 2363 13656 2404
rect 13622 2288 13656 2329
rect 13622 2213 13656 2254
rect 13622 2138 13656 2179
rect 13622 2063 13656 2104
rect 13714 3057 13748 3098
rect 13714 2982 13748 3023
rect 13714 2907 13748 2948
rect 13714 2832 13748 2873
rect 13714 2757 13748 2798
rect 13714 2682 13748 2723
rect 13714 2606 13748 2648
rect 13714 2530 13748 2572
rect 13714 2454 13748 2496
rect 13714 2378 13748 2420
rect 13714 2302 13748 2344
rect 13714 2226 13748 2268
rect 13714 2150 13748 2192
rect 13714 2074 13748 2116
rect 13806 3112 13840 3152
rect 13990 3260 14024 3300
rect 13990 3186 14024 3226
rect 13806 3038 13840 3078
rect 13806 2963 13840 3004
rect 13806 2888 13840 2929
rect 13806 2813 13840 2854
rect 13806 2738 13840 2779
rect 13806 2663 13840 2704
rect 13806 2588 13840 2629
rect 13806 2513 13840 2554
rect 13806 2438 13840 2479
rect 13806 2363 13840 2404
rect 13806 2288 13840 2329
rect 13806 2213 13840 2254
rect 13806 2138 13840 2179
rect 13806 2063 13840 2104
rect 13622 1988 13656 2029
rect 13898 3057 13932 3098
rect 13898 2982 13932 3023
rect 13898 2907 13932 2948
rect 13898 2832 13932 2873
rect 13898 2757 13932 2798
rect 13898 2682 13932 2723
rect 13898 2606 13932 2648
rect 13898 2530 13932 2572
rect 13898 2454 13932 2496
rect 13898 2378 13932 2420
rect 13898 2302 13932 2344
rect 13898 2226 13932 2268
rect 13898 2150 13932 2192
rect 13898 2074 13932 2116
rect 13990 3112 14024 3152
rect 14174 3260 14208 3300
rect 14174 3186 14208 3226
rect 13990 3038 14024 3078
rect 13990 2963 14024 3004
rect 13990 2888 14024 2929
rect 13990 2813 14024 2854
rect 13990 2738 14024 2779
rect 13990 2663 14024 2704
rect 13990 2588 14024 2629
rect 13990 2513 14024 2554
rect 13990 2438 14024 2479
rect 13990 2363 14024 2404
rect 13990 2288 14024 2329
rect 13990 2213 14024 2254
rect 13990 2138 14024 2179
rect 13990 2063 14024 2104
rect 13806 1988 13840 2029
rect 14082 3057 14116 3098
rect 14082 2982 14116 3023
rect 14082 2907 14116 2948
rect 14082 2832 14116 2873
rect 14082 2757 14116 2798
rect 14082 2682 14116 2723
rect 14082 2606 14116 2648
rect 14082 2530 14116 2572
rect 14082 2454 14116 2496
rect 14082 2378 14116 2420
rect 14082 2302 14116 2344
rect 14082 2226 14116 2268
rect 14082 2150 14116 2192
rect 14082 2074 14116 2116
rect 14174 3112 14208 3152
rect 14358 3260 14392 3300
rect 14358 3186 14392 3226
rect 14174 3038 14208 3078
rect 14174 2963 14208 3004
rect 14174 2888 14208 2929
rect 14174 2813 14208 2854
rect 14174 2738 14208 2779
rect 14174 2663 14208 2704
rect 14174 2588 14208 2629
rect 14174 2513 14208 2554
rect 14174 2438 14208 2479
rect 14174 2363 14208 2404
rect 14174 2288 14208 2329
rect 14174 2213 14208 2254
rect 14174 2138 14208 2179
rect 14174 2063 14208 2104
rect 13990 1988 14024 2029
rect 14266 3057 14300 3098
rect 14266 2982 14300 3023
rect 14266 2907 14300 2948
rect 14266 2832 14300 2873
rect 14266 2757 14300 2798
rect 14266 2682 14300 2723
rect 14266 2606 14300 2648
rect 14266 2530 14300 2572
rect 14266 2454 14300 2496
rect 14266 2378 14300 2420
rect 14266 2302 14300 2344
rect 14266 2226 14300 2268
rect 14266 2150 14300 2192
rect 14266 2074 14300 2116
rect 14358 3112 14392 3152
rect 14542 3260 14576 3300
rect 14542 3186 14576 3226
rect 14358 3038 14392 3078
rect 14358 2963 14392 3004
rect 14358 2888 14392 2929
rect 14358 2813 14392 2854
rect 14358 2738 14392 2779
rect 14358 2663 14392 2704
rect 14358 2588 14392 2629
rect 14358 2513 14392 2554
rect 14358 2438 14392 2479
rect 14358 2363 14392 2404
rect 14358 2288 14392 2329
rect 14358 2213 14392 2254
rect 14358 2138 14392 2179
rect 14358 2063 14392 2104
rect 14174 1988 14208 2029
rect 14450 3057 14484 3098
rect 14450 2982 14484 3023
rect 14450 2907 14484 2948
rect 14450 2832 14484 2873
rect 14450 2757 14484 2798
rect 14450 2682 14484 2723
rect 14450 2606 14484 2648
rect 14450 2530 14484 2572
rect 14450 2454 14484 2496
rect 14450 2378 14484 2420
rect 14450 2302 14484 2344
rect 14450 2226 14484 2268
rect 14450 2150 14484 2192
rect 14450 2074 14484 2116
rect 14542 3112 14576 3152
rect 14542 3038 14576 3078
rect 14542 2963 14576 3004
rect 14542 2888 14576 2929
rect 14542 2813 14576 2854
rect 14542 2738 14576 2779
rect 14542 2663 14576 2704
rect 14542 2588 14576 2629
rect 14542 2513 14576 2554
rect 14542 2438 14576 2479
rect 14542 2363 14576 2404
rect 14542 2288 14576 2329
rect 14542 2213 14576 2254
rect 14542 2138 14576 2179
rect 14542 2063 14576 2104
rect 14358 1988 14392 2029
rect 14542 1988 14576 2029
rect 14641 3310 14675 3344
rect 14641 3242 14675 3276
rect 14641 3174 14675 3204
rect 14641 3106 14675 3132
rect 14641 3038 14675 3060
rect 14641 2970 14675 2988
rect 14641 2902 14675 2916
rect 14641 2834 14675 2843
rect 14641 2766 14675 2770
rect 14641 2731 14675 2732
rect 14641 2658 14675 2664
rect 14641 2585 14675 2596
rect 14641 2512 14675 2528
rect 14641 2439 14675 2460
rect 14641 2366 14675 2392
rect 14641 2293 14675 2324
rect 14641 2222 14675 2256
rect 14641 2154 14675 2186
rect 14641 2086 14675 2113
rect 14641 2018 14675 2040
rect 13523 1922 13557 1924
rect 14641 1950 14675 1967
rect 13667 1864 13683 1898
rect 13717 1864 13756 1898
rect 13790 1864 13829 1898
rect 13863 1864 13902 1898
rect 13936 1864 13975 1898
rect 14009 1864 14048 1898
rect 14082 1864 14121 1898
rect 14155 1864 14193 1898
rect 14227 1864 14265 1898
rect 14299 1864 14337 1898
rect 14371 1864 14409 1898
rect 14443 1864 14481 1898
rect 14515 1864 14531 1898
rect 14641 1882 14675 1894
rect 13523 1849 13557 1856
rect 14641 1814 14675 1821
rect 13523 1776 13557 1788
rect 13523 1703 13557 1720
rect 13523 1630 13557 1652
rect 13523 1557 13557 1584
rect 13523 1484 13557 1516
rect 13523 1414 13557 1448
rect 13523 1346 13557 1377
rect 13523 1278 13557 1304
rect 13523 1210 13557 1232
rect 13523 1142 13557 1160
rect 13523 1074 13557 1088
rect 13523 1006 13557 1016
rect 13523 938 13557 944
rect 13523 870 13557 872
rect 13523 834 13557 836
rect 13523 762 13557 768
rect 13523 690 13557 700
rect 13622 1730 13656 1770
rect 13622 1656 13656 1696
rect 13622 1582 13656 1622
rect 13622 1508 13656 1548
rect 13622 1434 13656 1474
rect 13622 1360 13656 1400
rect 13622 1286 13656 1326
rect 13622 1212 13656 1252
rect 13622 1138 13656 1178
rect 13622 1064 13656 1104
rect 13622 990 13656 1030
rect 13622 915 13656 956
rect 13622 840 13656 881
rect 13622 765 13656 806
rect 13622 690 13656 731
rect 13714 1730 13748 1770
rect 13714 1656 13748 1696
rect 13714 1582 13748 1622
rect 13714 1508 13748 1548
rect 13714 1434 13748 1474
rect 13714 1360 13748 1400
rect 13714 1286 13748 1326
rect 13714 1212 13748 1252
rect 13714 1138 13748 1178
rect 13714 1064 13748 1104
rect 13714 990 13748 1030
rect 13714 916 13748 956
rect 13714 842 13748 882
rect 13714 768 13748 808
rect 13714 694 13748 734
rect 13523 598 13557 632
rect 13523 530 13557 564
rect 13714 619 13748 660
rect 13806 1730 13840 1770
rect 13806 1656 13840 1696
rect 13806 1582 13840 1622
rect 13806 1508 13840 1548
rect 13806 1434 13840 1474
rect 13806 1360 13840 1400
rect 13806 1286 13840 1326
rect 13806 1212 13840 1252
rect 13806 1138 13840 1178
rect 13806 1064 13840 1104
rect 13806 990 13840 1030
rect 13806 915 13840 956
rect 13806 840 13840 881
rect 13806 765 13840 806
rect 13806 690 13840 731
rect 13898 1730 13932 1770
rect 13898 1656 13932 1696
rect 13898 1582 13932 1622
rect 13898 1508 13932 1548
rect 13898 1434 13932 1474
rect 13898 1360 13932 1400
rect 13898 1286 13932 1326
rect 13898 1212 13932 1252
rect 13898 1138 13932 1178
rect 13898 1064 13932 1104
rect 13898 990 13932 1030
rect 13898 916 13932 956
rect 13898 842 13932 882
rect 13898 768 13932 808
rect 13898 694 13932 734
rect 13714 544 13748 585
rect 13898 619 13932 660
rect 13990 1730 14024 1770
rect 13990 1656 14024 1696
rect 13990 1582 14024 1622
rect 13990 1508 14024 1548
rect 13990 1434 14024 1474
rect 13990 1360 14024 1400
rect 13990 1286 14024 1326
rect 13990 1212 14024 1252
rect 13990 1138 14024 1178
rect 13990 1064 14024 1104
rect 13990 990 14024 1030
rect 13990 915 14024 956
rect 13990 840 14024 881
rect 13990 765 14024 806
rect 13990 690 14024 731
rect 14082 1730 14116 1770
rect 14082 1656 14116 1696
rect 14082 1582 14116 1622
rect 14082 1508 14116 1548
rect 14082 1434 14116 1474
rect 14082 1360 14116 1400
rect 14082 1286 14116 1326
rect 14082 1212 14116 1252
rect 14082 1138 14116 1178
rect 14082 1064 14116 1104
rect 14082 990 14116 1030
rect 14082 916 14116 956
rect 14082 842 14116 882
rect 14082 768 14116 808
rect 14082 694 14116 734
rect 13898 544 13932 585
rect 14082 619 14116 660
rect 14174 1730 14208 1770
rect 14174 1656 14208 1696
rect 14174 1582 14208 1622
rect 14174 1508 14208 1548
rect 14174 1434 14208 1474
rect 14174 1360 14208 1400
rect 14174 1286 14208 1326
rect 14174 1212 14208 1252
rect 14174 1138 14208 1178
rect 14174 1064 14208 1104
rect 14174 990 14208 1030
rect 14174 915 14208 956
rect 14174 840 14208 881
rect 14174 765 14208 806
rect 14174 690 14208 731
rect 14266 1730 14300 1770
rect 14266 1656 14300 1696
rect 14266 1582 14300 1622
rect 14266 1508 14300 1548
rect 14266 1434 14300 1474
rect 14266 1360 14300 1400
rect 14266 1286 14300 1326
rect 14266 1212 14300 1252
rect 14266 1138 14300 1178
rect 14266 1064 14300 1104
rect 14266 990 14300 1030
rect 14266 916 14300 956
rect 14266 842 14300 882
rect 14266 768 14300 808
rect 14266 694 14300 734
rect 14082 544 14116 585
rect 14266 619 14300 660
rect 14358 1730 14392 1770
rect 14358 1656 14392 1696
rect 14358 1582 14392 1622
rect 14358 1508 14392 1548
rect 14358 1434 14392 1474
rect 14358 1360 14392 1400
rect 14358 1286 14392 1326
rect 14358 1212 14392 1252
rect 14358 1138 14392 1178
rect 14358 1064 14392 1104
rect 14358 990 14392 1030
rect 14358 915 14392 956
rect 14358 840 14392 881
rect 14358 765 14392 806
rect 14358 690 14392 731
rect 14450 1730 14484 1770
rect 14450 1656 14484 1696
rect 14450 1582 14484 1622
rect 14450 1508 14484 1548
rect 14450 1434 14484 1474
rect 14450 1360 14484 1400
rect 14450 1286 14484 1326
rect 14450 1212 14484 1252
rect 14450 1138 14484 1178
rect 14450 1064 14484 1104
rect 14450 990 14484 1030
rect 14450 916 14484 956
rect 14450 842 14484 882
rect 14450 768 14484 808
rect 14450 694 14484 734
rect 14266 544 14300 585
rect 14450 619 14484 660
rect 14450 544 14484 585
rect 14542 1730 14576 1770
rect 14542 1656 14576 1696
rect 14542 1582 14576 1622
rect 14542 1508 14576 1548
rect 14542 1433 14576 1474
rect 14542 1358 14576 1399
rect 14542 1283 14576 1324
rect 14542 1208 14576 1249
rect 14542 1133 14576 1174
rect 14542 1058 14576 1099
rect 14542 983 14576 1024
rect 14542 908 14576 949
rect 14542 833 14576 874
rect 14542 758 14576 799
rect 14542 683 14576 724
rect 14542 608 14576 649
rect 14542 533 14576 574
rect 13523 462 13557 496
rect 13523 394 13557 428
rect 14542 458 14576 499
rect 14641 1746 14675 1748
rect 14641 1709 14675 1712
rect 14641 1636 14675 1644
rect 14641 1563 14675 1576
rect 14641 1490 14675 1508
rect 14641 1417 14675 1440
rect 14641 1344 14675 1372
rect 14641 1271 14675 1304
rect 14641 1202 14675 1236
rect 14641 1134 14675 1164
rect 14641 1066 14675 1091
rect 14641 998 14675 1018
rect 14641 930 14675 945
rect 14641 862 14675 872
rect 14641 794 14675 799
rect 14641 687 14675 692
rect 14641 614 14675 624
rect 14641 541 14675 556
rect 14641 468 14675 488
rect 14641 395 14675 420
rect 1669 306 1677 340
rect 1711 306 1747 340
rect 1781 322 1817 340
rect 1851 322 1887 340
rect 1921 322 1957 340
rect 1991 322 2027 340
rect 2061 322 2097 340
rect 2131 322 2167 340
rect 2201 322 2237 340
rect 2271 322 2307 340
rect 2341 322 2377 340
rect 2411 322 2447 340
rect 2481 322 2517 340
rect 1784 306 1817 322
rect 1857 306 1887 322
rect 1930 306 1957 322
rect 2003 306 2027 322
rect 2076 306 2097 322
rect 2149 306 2167 322
rect 2222 306 2237 322
rect 2295 306 2307 322
rect 2368 306 2377 322
rect 2441 306 2447 322
rect 2514 306 2517 322
rect 2551 322 2587 340
rect 2551 306 2553 322
rect 1669 288 1750 306
rect 1784 288 1823 306
rect 1857 288 1896 306
rect 1930 288 1969 306
rect 2003 288 2042 306
rect 2076 288 2115 306
rect 2149 288 2188 306
rect 2222 288 2261 306
rect 2295 288 2334 306
rect 2368 288 2407 306
rect 2441 288 2480 306
rect 2514 288 2553 306
rect 2621 322 2657 340
rect 2691 322 2727 340
rect 2761 322 2797 340
rect 2831 322 2867 340
rect 2901 322 2937 340
rect 2971 322 3007 340
rect 3041 322 3077 340
rect 3111 322 3147 340
rect 3181 322 3217 340
rect 2621 306 2626 322
rect 2691 306 2699 322
rect 2761 306 2772 322
rect 2831 306 2845 322
rect 2901 306 2918 322
rect 2971 306 2991 322
rect 3041 306 3064 322
rect 3111 306 3137 322
rect 3181 306 3210 322
rect 3251 306 3287 340
rect 3321 306 3331 340
rect 2587 288 2626 306
rect 2660 288 2699 306
rect 2733 288 2772 306
rect 2806 288 2845 306
rect 2879 288 2918 306
rect 2952 288 2991 306
rect 3025 288 3064 306
rect 3098 288 3137 306
rect 3171 288 3210 306
rect 3244 288 3331 306
rect 1669 282 3331 288
rect 1388 238 1422 272
rect 13523 250 13557 360
rect 13667 334 13679 368
rect 13717 334 13753 368
rect 13790 334 13827 368
rect 13863 334 13901 368
rect 13936 334 13974 368
rect 14009 334 14047 368
rect 14082 334 14120 368
rect 14155 334 14193 368
rect 14227 334 14265 368
rect 14300 334 14337 368
rect 14373 334 14409 368
rect 14446 334 14481 368
rect 14519 334 14531 368
rect 14641 322 14675 352
rect 14641 250 14675 284
rect 270 204 338 238
rect 372 204 406 238
rect 440 204 474 238
rect 508 204 542 238
rect 576 204 610 238
rect 644 204 678 238
rect 712 204 746 238
rect 780 204 814 238
rect 848 204 882 238
rect 916 204 950 238
rect 984 204 1018 238
rect 1052 204 1086 238
rect 1120 204 1154 238
rect 1188 204 1222 238
rect 1256 204 1290 238
rect 1324 204 1422 238
rect 13556 216 13591 250
rect 13631 216 13659 250
rect 13706 216 13727 250
rect 13781 216 13795 250
rect 13856 216 13863 250
rect 13965 216 13972 250
rect 14033 216 14047 250
rect 14101 216 14122 250
rect 14169 216 14197 250
rect 14237 216 14271 250
rect 14305 216 14339 250
rect 14379 216 14407 250
rect 14453 216 14475 250
rect 14527 216 14543 250
rect 14601 216 14675 250
<< viali >>
rect 14775 39522 14809 39556
rect 14917 39522 14951 39556
rect 2163 39474 10189 39476
rect 10228 39474 10262 39476
rect 10301 39474 10335 39476
rect 10374 39474 10408 39476
rect 10447 39474 10481 39476
rect 10520 39474 10554 39476
rect 10593 39474 10627 39476
rect 10666 39474 10700 39476
rect 10739 39474 10773 39476
rect 10812 39474 10846 39476
rect 10885 39474 10919 39476
rect 10958 39474 10992 39476
rect 11031 39474 11065 39476
rect 11104 39474 11138 39476
rect 11177 39474 11211 39476
rect 11250 39474 11284 39476
rect 11323 39474 11357 39476
rect 11396 39474 11430 39476
rect 11469 39474 11503 39476
rect 11542 39474 11576 39476
rect 11615 39474 11649 39476
rect 11688 39474 11722 39476
rect 11761 39474 11795 39476
rect 11834 39474 11868 39476
rect 11907 39474 11941 39476
rect 11980 39474 12014 39476
rect 12053 39474 12087 39476
rect 12126 39474 12160 39476
rect 12199 39474 12233 39476
rect 12272 39474 12306 39476
rect 12345 39474 12379 39476
rect 12418 39474 12452 39476
rect 12491 39474 12525 39476
rect 12564 39474 12598 39476
rect 12637 39474 12671 39476
rect 12710 39474 12744 39476
rect 12783 39474 12817 39476
rect 12856 39474 12890 39476
rect 12929 39474 12963 39476
rect 13002 39474 13036 39476
rect 13075 39474 13109 39476
rect 13148 39474 13182 39476
rect 13221 39474 13255 39476
rect 13294 39474 13328 39476
rect 13367 39474 13401 39476
rect 13440 39474 13474 39476
rect 13513 39474 13547 39476
rect 13586 39474 13620 39476
rect 13659 39474 13693 39476
rect 13732 39474 13766 39476
rect 1684 39272 1718 39284
rect 1684 39250 1718 39272
rect 1684 39204 1718 39212
rect 1684 39178 1718 39204
rect 1944 39406 2050 39470
rect 1944 34108 1946 39406
rect 1946 34108 2048 39406
rect 2048 34108 2050 39406
rect 2163 39372 10189 39474
rect 10228 39442 10262 39474
rect 10301 39442 10335 39474
rect 10374 39442 10408 39474
rect 10447 39442 10481 39474
rect 10520 39442 10554 39474
rect 10593 39442 10627 39474
rect 10666 39442 10700 39474
rect 10739 39442 10773 39474
rect 10812 39442 10846 39474
rect 10885 39442 10919 39474
rect 10958 39442 10992 39474
rect 11031 39442 11065 39474
rect 11104 39442 11138 39474
rect 11177 39442 11211 39474
rect 11250 39442 11284 39474
rect 11323 39442 11357 39474
rect 11396 39442 11430 39474
rect 11469 39442 11503 39474
rect 11542 39442 11576 39474
rect 11615 39442 11649 39474
rect 11688 39442 11722 39474
rect 11761 39442 11795 39474
rect 11834 39442 11868 39474
rect 11907 39442 11941 39474
rect 11980 39442 12014 39474
rect 12053 39442 12087 39474
rect 12126 39442 12160 39474
rect 12199 39442 12233 39474
rect 12272 39442 12306 39474
rect 12345 39442 12379 39474
rect 12418 39442 12452 39474
rect 12491 39442 12525 39474
rect 12564 39442 12598 39474
rect 12637 39442 12671 39474
rect 12710 39442 12744 39474
rect 12783 39442 12817 39474
rect 12856 39442 12890 39474
rect 12929 39442 12963 39474
rect 13002 39442 13036 39474
rect 13075 39442 13109 39474
rect 13148 39442 13182 39474
rect 13221 39442 13255 39474
rect 13294 39442 13328 39474
rect 13367 39442 13401 39474
rect 13440 39442 13474 39474
rect 13513 39442 13547 39474
rect 13586 39442 13620 39474
rect 13659 39442 13693 39474
rect 13732 39442 13766 39474
rect 10228 39372 10262 39404
rect 10301 39372 10335 39404
rect 10374 39372 10408 39404
rect 10447 39372 10481 39404
rect 10520 39372 10554 39404
rect 10593 39372 10627 39404
rect 10666 39372 10700 39404
rect 10739 39372 10773 39404
rect 10812 39372 10846 39404
rect 10885 39372 10919 39404
rect 10958 39372 10992 39404
rect 11031 39372 11065 39404
rect 11104 39372 11138 39404
rect 11177 39372 11211 39404
rect 11250 39372 11284 39404
rect 11323 39372 11357 39404
rect 11396 39372 11430 39404
rect 11469 39372 11503 39404
rect 11542 39372 11576 39404
rect 11615 39372 11649 39404
rect 11688 39372 11722 39404
rect 11761 39372 11795 39404
rect 11834 39372 11868 39404
rect 11907 39372 11941 39404
rect 11980 39372 12014 39404
rect 12053 39372 12087 39404
rect 12126 39372 12160 39404
rect 12199 39372 12233 39404
rect 12272 39372 12306 39404
rect 12345 39372 12379 39404
rect 12418 39372 12452 39404
rect 12491 39372 12525 39404
rect 12564 39372 12598 39404
rect 12637 39372 12671 39404
rect 12710 39372 12744 39404
rect 12783 39372 12817 39404
rect 12856 39372 12890 39404
rect 12929 39372 12963 39404
rect 13002 39372 13036 39404
rect 13075 39372 13109 39404
rect 13148 39372 13182 39404
rect 13221 39372 13255 39404
rect 13294 39372 13328 39404
rect 13367 39372 13401 39404
rect 13440 39372 13474 39404
rect 13513 39372 13547 39404
rect 13586 39372 13620 39404
rect 13659 39372 13693 39404
rect 13732 39372 13766 39404
rect 13838 39372 13874 39470
rect 13874 39372 13944 39470
rect 14775 39384 14809 39418
rect 14917 39384 14951 39418
rect 2163 39370 10189 39372
rect 10228 39370 10262 39372
rect 10301 39370 10335 39372
rect 10374 39370 10408 39372
rect 10447 39370 10481 39372
rect 10520 39370 10554 39372
rect 10593 39370 10627 39372
rect 10666 39370 10700 39372
rect 10739 39370 10773 39372
rect 10812 39370 10846 39372
rect 10885 39370 10919 39372
rect 10958 39370 10992 39372
rect 11031 39370 11065 39372
rect 11104 39370 11138 39372
rect 11177 39370 11211 39372
rect 11250 39370 11284 39372
rect 11323 39370 11357 39372
rect 11396 39370 11430 39372
rect 11469 39370 11503 39372
rect 11542 39370 11576 39372
rect 11615 39370 11649 39372
rect 11688 39370 11722 39372
rect 11761 39370 11795 39372
rect 11834 39370 11868 39372
rect 11907 39370 11941 39372
rect 11980 39370 12014 39372
rect 12053 39370 12087 39372
rect 12126 39370 12160 39372
rect 12199 39370 12233 39372
rect 12272 39370 12306 39372
rect 12345 39370 12379 39372
rect 12418 39370 12452 39372
rect 12491 39370 12525 39372
rect 12564 39370 12598 39372
rect 12637 39370 12671 39372
rect 12710 39370 12744 39372
rect 12783 39370 12817 39372
rect 12856 39370 12890 39372
rect 12929 39370 12963 39372
rect 13002 39370 13036 39372
rect 13075 39370 13109 39372
rect 13148 39370 13182 39372
rect 13221 39370 13255 39372
rect 13294 39370 13328 39372
rect 13367 39370 13401 39372
rect 13440 39370 13474 39372
rect 13513 39370 13547 39372
rect 13586 39370 13620 39372
rect 13659 39370 13693 39372
rect 13732 39370 13766 39372
rect 13838 39355 13944 39372
rect 13838 39321 13908 39355
rect 13908 39321 13942 39355
rect 13942 39321 13944 39355
rect 13838 39287 13944 39321
rect 1944 34035 1946 34069
rect 1946 34035 1978 34069
rect 2016 34035 2048 34069
rect 2048 34035 2050 34069
rect 1944 33962 1946 33996
rect 1946 33962 1978 33996
rect 2016 33962 2048 33996
rect 2048 33962 2050 33996
rect 1944 33889 1946 33923
rect 1946 33889 1978 33923
rect 2016 33889 2048 33923
rect 2048 33889 2050 33923
rect 1944 33816 1946 33850
rect 1946 33816 1978 33850
rect 2016 33816 2048 33850
rect 2048 33816 2050 33850
rect 1944 33743 1946 33777
rect 1946 33743 1978 33777
rect 2016 33743 2048 33777
rect 2048 33743 2050 33777
rect 1944 33670 1946 33704
rect 1946 33670 1978 33704
rect 2016 33670 2048 33704
rect 2048 33670 2050 33704
rect 1837 19864 1871 19898
rect 1909 19864 1943 19898
rect 1837 19787 1871 19821
rect 1909 19787 1943 19821
rect 1837 19710 1871 19744
rect 1909 19710 1943 19744
rect 1837 19633 1871 19667
rect 1909 19633 1943 19667
rect 2291 39153 9957 39171
rect 9996 39153 10030 39171
rect 10069 39153 10103 39171
rect 10142 39153 10176 39171
rect 10215 39153 10249 39171
rect 2291 39119 2482 39153
rect 2482 39119 2516 39153
rect 2516 39119 2550 39153
rect 2550 39119 2584 39153
rect 2584 39119 2618 39153
rect 2618 39119 2652 39153
rect 2652 39119 2686 39153
rect 2686 39119 2720 39153
rect 2720 39119 2754 39153
rect 2754 39119 2788 39153
rect 2788 39119 2822 39153
rect 2822 39119 2856 39153
rect 2856 39119 2890 39153
rect 2890 39119 2924 39153
rect 2924 39119 2958 39153
rect 2958 39119 2992 39153
rect 2992 39119 3026 39153
rect 3026 39119 3060 39153
rect 3060 39119 3094 39153
rect 3094 39119 3128 39153
rect 3128 39119 3162 39153
rect 3162 39119 3196 39153
rect 3196 39119 3230 39153
rect 3230 39119 3264 39153
rect 3264 39119 3298 39153
rect 3298 39119 3332 39153
rect 3332 39119 3366 39153
rect 3366 39119 3400 39153
rect 3400 39119 3434 39153
rect 3434 39119 3468 39153
rect 3468 39119 3502 39153
rect 3502 39119 3536 39153
rect 3536 39119 3570 39153
rect 3570 39119 3604 39153
rect 3604 39119 3638 39153
rect 3638 39119 3672 39153
rect 3672 39119 3706 39153
rect 3706 39119 3740 39153
rect 3740 39119 3774 39153
rect 3774 39119 3808 39153
rect 3808 39119 3842 39153
rect 3842 39119 3876 39153
rect 3876 39119 3910 39153
rect 3910 39119 3944 39153
rect 3944 39119 3978 39153
rect 3978 39119 4012 39153
rect 4012 39119 4046 39153
rect 4046 39119 4080 39153
rect 4080 39119 4114 39153
rect 4114 39119 4148 39153
rect 4148 39119 4182 39153
rect 4182 39119 4216 39153
rect 4216 39119 4250 39153
rect 4250 39119 4284 39153
rect 4284 39119 4318 39153
rect 4318 39119 4352 39153
rect 4352 39119 4386 39153
rect 4386 39119 4420 39153
rect 4420 39119 4454 39153
rect 4454 39119 4488 39153
rect 4488 39119 4522 39153
rect 4522 39119 4556 39153
rect 4556 39119 4590 39153
rect 4590 39119 4624 39153
rect 4624 39119 4658 39153
rect 4658 39119 4692 39153
rect 4692 39119 4726 39153
rect 4726 39119 4760 39153
rect 4760 39119 4794 39153
rect 4794 39119 4828 39153
rect 4828 39119 4862 39153
rect 4862 39119 4896 39153
rect 4896 39119 4930 39153
rect 4930 39119 4964 39153
rect 4964 39119 4998 39153
rect 4998 39119 5032 39153
rect 5032 39119 5066 39153
rect 5066 39119 5100 39153
rect 5100 39119 5134 39153
rect 5134 39119 5168 39153
rect 5168 39119 5202 39153
rect 5202 39119 5236 39153
rect 5236 39119 5270 39153
rect 5270 39119 5304 39153
rect 5304 39119 5338 39153
rect 5338 39119 5372 39153
rect 5372 39119 5406 39153
rect 5406 39119 5440 39153
rect 5440 39119 5474 39153
rect 5474 39119 5508 39153
rect 5508 39119 5542 39153
rect 5542 39119 5576 39153
rect 5576 39119 5610 39153
rect 5610 39119 5644 39153
rect 5644 39119 5678 39153
rect 5678 39119 5712 39153
rect 5712 39119 5746 39153
rect 5746 39119 5780 39153
rect 5780 39119 5814 39153
rect 5814 39119 5848 39153
rect 5848 39119 5882 39153
rect 5882 39119 5916 39153
rect 5916 39119 5950 39153
rect 5950 39119 5984 39153
rect 5984 39119 6018 39153
rect 6018 39119 6052 39153
rect 6052 39119 6086 39153
rect 6086 39119 6120 39153
rect 6120 39119 6154 39153
rect 6154 39119 6188 39153
rect 6188 39119 6222 39153
rect 6222 39119 6256 39153
rect 6256 39119 6290 39153
rect 6290 39119 6324 39153
rect 6324 39119 6358 39153
rect 6358 39119 6392 39153
rect 6392 39119 6426 39153
rect 6426 39119 6460 39153
rect 6460 39119 6494 39153
rect 6494 39119 6528 39153
rect 6528 39119 6562 39153
rect 6562 39119 6596 39153
rect 6596 39119 6630 39153
rect 6630 39119 6664 39153
rect 6664 39119 6698 39153
rect 6698 39119 6732 39153
rect 6732 39119 6766 39153
rect 6766 39119 6800 39153
rect 6800 39119 6834 39153
rect 6834 39119 6868 39153
rect 6868 39119 6902 39153
rect 6902 39119 6936 39153
rect 6936 39119 6970 39153
rect 6970 39119 7004 39153
rect 7004 39119 7038 39153
rect 7038 39119 7072 39153
rect 7072 39119 7106 39153
rect 7106 39119 7140 39153
rect 7140 39119 7174 39153
rect 7174 39119 7208 39153
rect 7208 39119 7242 39153
rect 7242 39119 7276 39153
rect 7276 39119 7310 39153
rect 7310 39119 7344 39153
rect 7344 39119 7378 39153
rect 7378 39119 7412 39153
rect 7412 39119 7446 39153
rect 7446 39119 7480 39153
rect 7480 39119 7514 39153
rect 7514 39119 7548 39153
rect 7548 39119 7582 39153
rect 7582 39119 7616 39153
rect 7616 39119 7650 39153
rect 7650 39119 7684 39153
rect 7684 39119 7718 39153
rect 7718 39119 7752 39153
rect 7752 39119 7786 39153
rect 7786 39119 7820 39153
rect 7820 39119 7854 39153
rect 7854 39119 7888 39153
rect 7888 39119 7922 39153
rect 7922 39119 7956 39153
rect 7956 39119 7990 39153
rect 7990 39119 8024 39153
rect 8024 39119 8058 39153
rect 8058 39119 8092 39153
rect 8092 39119 8126 39153
rect 8126 39119 8160 39153
rect 8160 39119 8194 39153
rect 8194 39119 8228 39153
rect 8228 39119 8262 39153
rect 8262 39119 8296 39153
rect 8296 39119 8330 39153
rect 8330 39119 8364 39153
rect 8364 39119 8398 39153
rect 8398 39119 8432 39153
rect 8432 39119 8466 39153
rect 8466 39119 8500 39153
rect 8500 39119 8534 39153
rect 8534 39119 8568 39153
rect 8568 39119 8602 39153
rect 8602 39119 8636 39153
rect 8636 39119 8670 39153
rect 8670 39119 8704 39153
rect 8704 39119 8738 39153
rect 8738 39119 8772 39153
rect 8772 39119 8806 39153
rect 8806 39119 8840 39153
rect 8840 39119 8874 39153
rect 8874 39119 8908 39153
rect 8908 39119 8943 39153
rect 8943 39119 8977 39153
rect 8977 39119 9012 39153
rect 9012 39119 9046 39153
rect 9046 39119 9081 39153
rect 9081 39119 9115 39153
rect 9115 39119 9150 39153
rect 9150 39119 9184 39153
rect 9184 39119 9219 39153
rect 9219 39119 9253 39153
rect 9253 39119 9288 39153
rect 9288 39119 9322 39153
rect 9322 39119 9357 39153
rect 9357 39119 9391 39153
rect 9391 39119 9426 39153
rect 9426 39119 9460 39153
rect 9460 39119 9495 39153
rect 9495 39119 9529 39153
rect 9529 39119 9564 39153
rect 9564 39119 9598 39153
rect 9598 39119 9633 39153
rect 9633 39119 9667 39153
rect 9667 39119 9702 39153
rect 9702 39119 9736 39153
rect 9736 39119 9771 39153
rect 9771 39119 9805 39153
rect 9805 39119 9840 39153
rect 9840 39119 9874 39153
rect 9874 39119 9909 39153
rect 9909 39119 9943 39153
rect 9943 39119 9957 39153
rect 9996 39137 10012 39153
rect 10012 39137 10030 39153
rect 10069 39137 10081 39153
rect 10081 39137 10103 39153
rect 10142 39137 10150 39153
rect 10150 39137 10176 39153
rect 10215 39137 10219 39153
rect 10219 39137 10249 39153
rect 10288 39137 10322 39171
rect 10361 39153 10395 39171
rect 10434 39153 10468 39171
rect 10507 39153 10541 39171
rect 10580 39153 10614 39171
rect 10653 39153 10687 39171
rect 10726 39153 10760 39171
rect 10799 39153 10833 39171
rect 10872 39153 10906 39171
rect 10945 39153 10979 39171
rect 11018 39153 11052 39171
rect 11091 39153 11125 39171
rect 11164 39153 11198 39171
rect 11237 39153 11271 39171
rect 11310 39153 11344 39171
rect 11383 39153 11417 39171
rect 11456 39153 11490 39171
rect 11529 39153 11563 39171
rect 11602 39153 11636 39171
rect 11675 39153 11709 39171
rect 11748 39153 11782 39171
rect 11821 39153 11855 39171
rect 11894 39153 11928 39171
rect 11967 39153 12001 39171
rect 12040 39153 12074 39171
rect 12113 39153 12147 39171
rect 12186 39153 12220 39171
rect 12259 39153 12293 39171
rect 12332 39153 12366 39171
rect 12405 39153 12439 39171
rect 12478 39153 12512 39171
rect 12551 39153 12585 39171
rect 12624 39153 12658 39171
rect 12697 39153 12731 39171
rect 12770 39153 12804 39171
rect 12843 39153 12877 39171
rect 12916 39153 12950 39171
rect 12989 39153 13095 39171
rect 13137 39153 13171 39171
rect 13213 39153 13247 39171
rect 13289 39153 13323 39171
rect 13365 39153 13399 39171
rect 13441 39153 13475 39171
rect 10361 39137 10392 39153
rect 10392 39137 10395 39153
rect 10434 39137 10461 39153
rect 10461 39137 10468 39153
rect 10507 39137 10530 39153
rect 10530 39137 10541 39153
rect 10580 39137 10599 39153
rect 10599 39137 10614 39153
rect 10653 39137 10668 39153
rect 10668 39137 10687 39153
rect 10726 39137 10737 39153
rect 10737 39137 10760 39153
rect 10799 39137 10806 39153
rect 10806 39137 10833 39153
rect 10872 39137 10875 39153
rect 10875 39137 10906 39153
rect 10945 39137 10978 39153
rect 10978 39137 10979 39153
rect 11018 39137 11047 39153
rect 11047 39137 11052 39153
rect 11091 39137 11116 39153
rect 11116 39137 11125 39153
rect 11164 39137 11185 39153
rect 11185 39137 11198 39153
rect 11237 39137 11254 39153
rect 11254 39137 11271 39153
rect 11310 39137 11323 39153
rect 11323 39137 11344 39153
rect 11383 39137 11392 39153
rect 11392 39137 11417 39153
rect 11456 39137 11461 39153
rect 11461 39137 11490 39153
rect 11529 39137 11530 39153
rect 11530 39137 11563 39153
rect 11602 39137 11634 39153
rect 11634 39137 11636 39153
rect 11675 39137 11703 39153
rect 11703 39137 11709 39153
rect 11748 39137 11772 39153
rect 11772 39137 11782 39153
rect 11821 39137 11841 39153
rect 11841 39137 11855 39153
rect 11894 39137 11910 39153
rect 11910 39137 11928 39153
rect 11967 39137 11979 39153
rect 11979 39137 12001 39153
rect 12040 39137 12048 39153
rect 12048 39137 12074 39153
rect 12113 39137 12117 39153
rect 12117 39137 12147 39153
rect 12186 39137 12220 39153
rect 12259 39137 12289 39153
rect 12289 39137 12293 39153
rect 12332 39137 12358 39153
rect 12358 39137 12366 39153
rect 12405 39137 12427 39153
rect 12427 39137 12439 39153
rect 12478 39137 12496 39153
rect 12496 39137 12512 39153
rect 12551 39137 12565 39153
rect 12565 39137 12585 39153
rect 12624 39137 12634 39153
rect 12634 39137 12658 39153
rect 12697 39137 12703 39153
rect 12703 39137 12731 39153
rect 12770 39137 12772 39153
rect 12772 39137 12804 39153
rect 12843 39137 12876 39153
rect 12876 39137 12877 39153
rect 12916 39137 12945 39153
rect 12945 39137 12950 39153
rect 12989 39119 13014 39153
rect 13014 39119 13048 39153
rect 13048 39119 13083 39153
rect 13083 39119 13095 39153
rect 13137 39137 13152 39153
rect 13152 39137 13171 39153
rect 13213 39137 13221 39153
rect 13221 39137 13247 39153
rect 13289 39137 13290 39153
rect 13290 39137 13323 39153
rect 13365 39137 13393 39153
rect 13393 39137 13399 39153
rect 13441 39137 13462 39153
rect 13462 39137 13475 39153
rect 13517 39137 13551 39171
rect 13593 39137 13627 39171
rect 2219 39065 2253 39099
rect 2291 39065 2444 39119
rect 2219 38992 2253 39026
rect 2291 38992 2325 39026
rect 2363 38993 2444 39065
rect 2444 39027 9957 39119
rect 9996 39065 10030 39099
rect 10069 39065 10103 39099
rect 10142 39065 10176 39099
rect 10215 39065 10249 39099
rect 10288 39065 10322 39099
rect 10361 39065 10395 39099
rect 10434 39065 10468 39099
rect 10507 39065 10541 39099
rect 10580 39065 10614 39099
rect 10653 39065 10687 39099
rect 10726 39065 10760 39099
rect 10799 39065 10833 39099
rect 10872 39065 10906 39099
rect 10945 39065 10979 39099
rect 11018 39065 11052 39099
rect 11091 39065 11125 39099
rect 11164 39065 11198 39099
rect 11237 39065 11271 39099
rect 11310 39065 11344 39099
rect 11383 39065 11417 39099
rect 11456 39065 11490 39099
rect 11529 39065 11563 39099
rect 11602 39065 11636 39099
rect 11675 39065 11709 39099
rect 11748 39065 11782 39099
rect 11821 39065 11855 39099
rect 11894 39065 11928 39099
rect 11967 39065 12001 39099
rect 12040 39065 12074 39099
rect 12113 39065 12147 39099
rect 12186 39065 12220 39099
rect 12259 39065 12293 39099
rect 12332 39065 12366 39099
rect 12405 39065 12439 39099
rect 12478 39065 12512 39099
rect 12551 39065 12585 39099
rect 12624 39065 12658 39099
rect 12697 39065 12731 39099
rect 12770 39065 12804 39099
rect 12843 39065 12877 39099
rect 12916 39065 12950 39099
rect 12989 39027 13095 39119
rect 13137 39065 13171 39099
rect 13213 39065 13247 39099
rect 13289 39065 13323 39099
rect 13365 39065 13399 39099
rect 13441 39065 13475 39099
rect 13517 39065 13551 39099
rect 13593 39027 13617 39099
rect 2444 38993 2482 39027
rect 2482 38993 2516 39027
rect 2516 38993 2550 39027
rect 2550 38993 2584 39027
rect 2584 38993 2618 39027
rect 2618 38993 2652 39027
rect 2652 38993 2686 39027
rect 2686 38993 2720 39027
rect 2720 38993 2754 39027
rect 2754 38993 2788 39027
rect 2788 38993 2822 39027
rect 2822 38993 2856 39027
rect 2856 38993 2890 39027
rect 2890 38993 2924 39027
rect 2924 38993 2958 39027
rect 2958 38993 2992 39027
rect 2992 38993 3026 39027
rect 3026 38993 3060 39027
rect 3060 38993 3094 39027
rect 3094 38993 3128 39027
rect 3128 38993 3162 39027
rect 3162 38993 3196 39027
rect 3196 38993 3230 39027
rect 3230 38993 3264 39027
rect 3264 38993 3298 39027
rect 3298 38993 3332 39027
rect 3332 38993 3366 39027
rect 3366 38993 3400 39027
rect 3400 38993 3434 39027
rect 3434 38993 3468 39027
rect 3468 38993 3502 39027
rect 3502 38993 3536 39027
rect 3536 38993 3570 39027
rect 3570 38993 3604 39027
rect 3604 38993 3638 39027
rect 3638 38993 3672 39027
rect 3672 38993 3706 39027
rect 3706 38993 3740 39027
rect 3740 38993 3774 39027
rect 3774 38993 3808 39027
rect 3808 38993 3842 39027
rect 3842 38993 3876 39027
rect 3876 38993 3910 39027
rect 3910 38993 3944 39027
rect 3944 38993 3978 39027
rect 3978 38993 4012 39027
rect 4012 38993 4046 39027
rect 4046 38993 4080 39027
rect 4080 38993 4114 39027
rect 4114 38993 4148 39027
rect 4148 38993 4182 39027
rect 4182 38993 4216 39027
rect 4216 38993 4250 39027
rect 4250 38993 4284 39027
rect 4284 38993 4318 39027
rect 4318 38993 4352 39027
rect 4352 38993 4386 39027
rect 4386 38993 4420 39027
rect 4420 38993 4454 39027
rect 4454 38993 4488 39027
rect 4488 38993 4522 39027
rect 4522 38993 4556 39027
rect 4556 38993 4590 39027
rect 4590 38993 4624 39027
rect 4624 38993 4658 39027
rect 4658 38993 4692 39027
rect 4692 38993 4726 39027
rect 4726 38993 4760 39027
rect 4760 38993 4794 39027
rect 4794 38993 4828 39027
rect 4828 38993 4862 39027
rect 4862 38993 4896 39027
rect 4896 38993 4930 39027
rect 4930 38993 4964 39027
rect 4964 38993 4998 39027
rect 4998 38993 5032 39027
rect 5032 38993 5066 39027
rect 5066 38993 5100 39027
rect 5100 38993 5134 39027
rect 5134 38993 5168 39027
rect 5168 38993 5202 39027
rect 5202 38993 5236 39027
rect 5236 38993 5270 39027
rect 5270 38993 5304 39027
rect 5304 38993 5338 39027
rect 5338 38993 5372 39027
rect 5372 38993 5406 39027
rect 5406 38993 5440 39027
rect 5440 38993 5474 39027
rect 5474 38993 5508 39027
rect 5508 38993 5542 39027
rect 5542 38993 5576 39027
rect 5576 38993 5610 39027
rect 5610 38993 5644 39027
rect 5644 38993 5678 39027
rect 5678 38993 5712 39027
rect 5712 38993 5746 39027
rect 5746 38993 5780 39027
rect 5780 38993 5814 39027
rect 5814 38993 5848 39027
rect 5848 38993 5882 39027
rect 5882 38993 5916 39027
rect 5916 38993 5950 39027
rect 5950 38993 5984 39027
rect 5984 38993 6018 39027
rect 6018 38993 6052 39027
rect 6052 38993 6086 39027
rect 6086 38993 6120 39027
rect 6120 38993 6154 39027
rect 6154 38993 6188 39027
rect 6188 38993 6222 39027
rect 6222 38993 6256 39027
rect 6256 38993 6290 39027
rect 6290 38993 6324 39027
rect 6324 38993 6358 39027
rect 6358 38993 6392 39027
rect 6392 38993 6426 39027
rect 6426 38993 6460 39027
rect 6460 38993 6494 39027
rect 6494 38993 6528 39027
rect 6528 38993 6562 39027
rect 6562 38993 6596 39027
rect 6596 38993 6630 39027
rect 6630 38993 6664 39027
rect 6664 38993 6698 39027
rect 6698 38993 6732 39027
rect 6732 38993 6766 39027
rect 6766 38993 6800 39027
rect 6800 38993 6834 39027
rect 6834 38993 6868 39027
rect 6868 38993 6902 39027
rect 6902 38993 6936 39027
rect 6936 38993 6970 39027
rect 6970 38993 7004 39027
rect 7004 38993 7038 39027
rect 7038 38993 7072 39027
rect 7072 38993 7106 39027
rect 7106 38993 7140 39027
rect 7140 38993 7174 39027
rect 7174 38993 7208 39027
rect 7208 38993 7242 39027
rect 7242 38993 7276 39027
rect 7276 38993 7310 39027
rect 7310 38993 7344 39027
rect 7344 38993 7378 39027
rect 7378 38993 7412 39027
rect 7412 38993 7446 39027
rect 7446 38993 7480 39027
rect 7480 38993 7514 39027
rect 7514 38993 7548 39027
rect 7548 38993 7582 39027
rect 7582 38993 7616 39027
rect 7616 38993 7650 39027
rect 7650 38993 7684 39027
rect 7684 38993 7718 39027
rect 7718 38993 7752 39027
rect 7752 38993 7786 39027
rect 7786 38993 7820 39027
rect 7820 38993 7854 39027
rect 7854 38993 7888 39027
rect 7888 38993 7922 39027
rect 7922 38993 7956 39027
rect 7956 38993 7990 39027
rect 7990 38993 8024 39027
rect 8024 38993 8058 39027
rect 8058 38993 8092 39027
rect 8092 38993 8126 39027
rect 8126 38993 8160 39027
rect 8160 38993 8194 39027
rect 8194 38993 8228 39027
rect 8228 38993 8262 39027
rect 8262 38993 8296 39027
rect 8296 38993 8330 39027
rect 8330 38993 8364 39027
rect 8364 38993 8398 39027
rect 8398 38993 8432 39027
rect 8432 38993 8466 39027
rect 8466 38993 8500 39027
rect 8500 38993 8534 39027
rect 8534 38993 8568 39027
rect 8568 38993 8602 39027
rect 8602 38993 8636 39027
rect 8636 38993 8670 39027
rect 8670 38993 8704 39027
rect 8704 38993 8738 39027
rect 8738 38993 8772 39027
rect 8772 38993 8806 39027
rect 8806 38993 8840 39027
rect 8840 38993 8874 39027
rect 8874 38993 8908 39027
rect 8908 38993 8943 39027
rect 8943 38993 8977 39027
rect 8977 38993 9012 39027
rect 9012 38993 9046 39027
rect 9046 38993 9081 39027
rect 9081 38993 9115 39027
rect 9115 38993 9150 39027
rect 9150 38993 9184 39027
rect 9184 38993 9219 39027
rect 9219 38993 9253 39027
rect 9253 38993 9288 39027
rect 9288 38993 9322 39027
rect 9322 38993 9357 39027
rect 9357 38993 9391 39027
rect 9391 38993 9426 39027
rect 9426 38993 9460 39027
rect 9460 38993 9495 39027
rect 9495 38993 9529 39027
rect 9529 38993 9564 39027
rect 9564 38993 9598 39027
rect 9598 38993 9633 39027
rect 9633 38993 9667 39027
rect 9667 38993 9702 39027
rect 9702 38993 9736 39027
rect 9736 38993 9771 39027
rect 9771 38993 9805 39027
rect 9805 38993 9840 39027
rect 9840 38993 9874 39027
rect 9874 38993 9909 39027
rect 9909 38993 9943 39027
rect 9943 38993 9957 39027
rect 9996 38993 10012 39027
rect 10012 38993 10030 39027
rect 10069 38993 10081 39027
rect 10081 38993 10103 39027
rect 10142 38993 10150 39027
rect 10150 38993 10176 39027
rect 10215 38993 10219 39027
rect 10219 38993 10249 39027
rect 10288 38993 10322 39027
rect 10361 38993 10392 39027
rect 10392 38993 10395 39027
rect 10434 38993 10461 39027
rect 10461 38993 10468 39027
rect 10507 38993 10530 39027
rect 10530 38993 10541 39027
rect 10580 38993 10599 39027
rect 10599 38993 10614 39027
rect 10653 38993 10668 39027
rect 10668 38993 10687 39027
rect 10726 38993 10737 39027
rect 10737 38993 10760 39027
rect 10799 38993 10806 39027
rect 10806 38993 10833 39027
rect 10872 38993 10875 39027
rect 10875 38993 10906 39027
rect 10945 38993 10978 39027
rect 10978 38993 10979 39027
rect 11018 38993 11047 39027
rect 11047 38993 11052 39027
rect 11091 38993 11116 39027
rect 11116 38993 11125 39027
rect 11164 38993 11185 39027
rect 11185 38993 11198 39027
rect 11237 38993 11254 39027
rect 11254 38993 11271 39027
rect 11310 38993 11323 39027
rect 11323 38993 11344 39027
rect 11383 38993 11392 39027
rect 11392 38993 11417 39027
rect 11456 38993 11461 39027
rect 11461 38993 11490 39027
rect 11529 38993 11530 39027
rect 11530 38993 11563 39027
rect 11602 38993 11634 39027
rect 11634 38993 11636 39027
rect 11675 38993 11703 39027
rect 11703 38993 11709 39027
rect 11748 38993 11772 39027
rect 11772 38993 11782 39027
rect 11821 38993 11841 39027
rect 11841 38993 11855 39027
rect 11894 38993 11910 39027
rect 11910 38993 11928 39027
rect 11967 38993 11979 39027
rect 11979 38993 12001 39027
rect 12040 38993 12048 39027
rect 12048 38993 12074 39027
rect 12113 38993 12117 39027
rect 12117 38993 12147 39027
rect 12186 38993 12220 39027
rect 12259 38993 12289 39027
rect 12289 38993 12293 39027
rect 12332 38993 12358 39027
rect 12358 38993 12366 39027
rect 12405 38993 12427 39027
rect 12427 38993 12439 39027
rect 12478 38993 12496 39027
rect 12496 38993 12512 39027
rect 12551 38993 12565 39027
rect 12565 38993 12585 39027
rect 12624 38993 12634 39027
rect 12634 38993 12658 39027
rect 12697 38993 12703 39027
rect 12703 38993 12731 39027
rect 12770 38993 12772 39027
rect 12772 38993 12804 39027
rect 12843 38993 12876 39027
rect 12876 38993 12877 39027
rect 12916 38993 12945 39027
rect 12945 38993 12950 39027
rect 12989 38993 13014 39027
rect 13014 38993 13048 39027
rect 13048 38993 13083 39027
rect 13083 38993 13095 39027
rect 13137 38993 13152 39027
rect 13152 38993 13171 39027
rect 13213 38993 13221 39027
rect 13221 38993 13247 39027
rect 13290 38993 13324 39027
rect 13367 38993 13393 39027
rect 13393 38993 13401 39027
rect 13444 38993 13462 39027
rect 13462 38993 13478 39027
rect 2219 38919 2253 38953
rect 2291 38919 2325 38953
rect 2363 38920 2397 38954
rect 2219 38846 2253 38880
rect 2291 38846 2325 38880
rect 2363 38847 2397 38881
rect 2884 38820 2888 38854
rect 2888 38820 2918 38854
rect 2957 38820 2991 38854
rect 3030 38820 3060 38854
rect 3060 38820 3064 38854
rect 3103 38820 3129 38854
rect 3129 38820 3137 38854
rect 3176 38820 3198 38854
rect 3198 38820 3210 38854
rect 3249 38820 3267 38854
rect 3267 38820 3283 38854
rect 3322 38820 3336 38854
rect 3336 38820 3356 38854
rect 3395 38820 3405 38854
rect 3405 38820 3429 38854
rect 3468 38820 3474 38854
rect 3474 38820 3502 38854
rect 3541 38820 3543 38854
rect 3543 38820 3575 38854
rect 3614 38820 3647 38854
rect 3647 38820 3648 38854
rect 3687 38820 3716 38854
rect 3716 38820 3721 38854
rect 3760 38820 3785 38854
rect 3785 38820 3794 38854
rect 3833 38820 3854 38854
rect 3854 38820 3867 38854
rect 3906 38820 3923 38854
rect 3923 38820 3940 38854
rect 3979 38820 3992 38854
rect 3992 38820 4013 38854
rect 4052 38820 4061 38854
rect 4061 38820 4086 38854
rect 4125 38820 4130 38854
rect 4130 38820 4159 38854
rect 4198 38820 4199 38854
rect 4199 38820 4232 38854
rect 4271 38820 4302 38854
rect 4302 38820 4305 38854
rect 4344 38820 4371 38854
rect 4371 38820 4378 38854
rect 4417 38820 4440 38854
rect 4440 38820 4451 38854
rect 4490 38820 4509 38854
rect 4509 38820 4524 38854
rect 4563 38820 4578 38854
rect 4578 38820 4597 38854
rect 4636 38820 4647 38854
rect 4647 38820 4670 38854
rect 4709 38820 4716 38854
rect 4716 38820 4743 38854
rect 4782 38820 4785 38854
rect 4785 38820 4816 38854
rect 4855 38820 4889 38854
rect 4928 38820 4958 38854
rect 4958 38820 4962 38854
rect 5001 38820 5027 38854
rect 5027 38820 5035 38854
rect 5074 38820 5096 38854
rect 5096 38820 5108 38854
rect 5147 38820 5165 38854
rect 5165 38820 5181 38854
rect 5220 38820 5234 38854
rect 5234 38820 5254 38854
rect 5293 38820 5303 38854
rect 5303 38820 5327 38854
rect 5366 38820 5372 38854
rect 5372 38820 5400 38854
rect 5439 38820 5441 38854
rect 5441 38820 5473 38854
rect 5512 38820 5544 38854
rect 5544 38820 5546 38854
rect 5584 38820 5613 38854
rect 5613 38820 5618 38854
rect 5656 38820 5682 38854
rect 5682 38820 5690 38854
rect 5728 38820 5751 38854
rect 5751 38820 5762 38854
rect 5800 38820 5820 38854
rect 5820 38820 5834 38854
rect 5872 38820 5889 38854
rect 5889 38820 5906 38854
rect 5944 38820 5958 38854
rect 5958 38820 5978 38854
rect 6016 38820 6027 38854
rect 6027 38820 6050 38854
rect 6088 38820 6096 38854
rect 6096 38820 6122 38854
rect 6160 38820 6165 38854
rect 6165 38820 6194 38854
rect 6232 38820 6234 38854
rect 6234 38820 6266 38854
rect 6304 38820 6336 38854
rect 6336 38820 6338 38854
rect 6376 38820 6404 38854
rect 6404 38820 6410 38854
rect 6448 38820 6472 38854
rect 6472 38820 6482 38854
rect 6520 38820 6540 38854
rect 6540 38820 6554 38854
rect 6592 38820 6608 38854
rect 6608 38820 6626 38854
rect 6664 38820 6676 38854
rect 6676 38820 6698 38854
rect 6736 38820 6744 38854
rect 6744 38820 6770 38854
rect 6808 38820 6812 38854
rect 6812 38820 6842 38854
rect 6880 38820 6914 38854
rect 6952 38820 6982 38854
rect 6982 38820 6986 38854
rect 7024 38820 7050 38854
rect 7050 38820 7058 38854
rect 7096 38820 7118 38854
rect 7118 38820 7130 38854
rect 7168 38820 7186 38854
rect 7186 38820 7202 38854
rect 7240 38820 7254 38854
rect 7254 38820 7274 38854
rect 7312 38820 7322 38854
rect 7322 38820 7346 38854
rect 7384 38820 7390 38854
rect 7390 38820 7418 38854
rect 7456 38820 7458 38854
rect 7458 38820 7490 38854
rect 7528 38820 7560 38854
rect 7560 38820 7562 38854
rect 7600 38820 7628 38854
rect 7628 38820 7634 38854
rect 7672 38820 7696 38854
rect 7696 38820 7706 38854
rect 7744 38820 7764 38854
rect 7764 38820 7778 38854
rect 7816 38820 7832 38854
rect 7832 38820 7850 38854
rect 7888 38820 7900 38854
rect 7900 38820 7922 38854
rect 7960 38820 7968 38854
rect 7968 38820 7994 38854
rect 8032 38820 8036 38854
rect 8036 38820 8066 38854
rect 8104 38820 8138 38854
rect 8176 38820 8206 38854
rect 8206 38820 8210 38854
rect 8248 38820 8274 38854
rect 8274 38820 8282 38854
rect 8320 38820 8342 38854
rect 8342 38820 8354 38854
rect 8392 38820 8410 38854
rect 8410 38820 8426 38854
rect 8464 38820 8478 38854
rect 8478 38820 8498 38854
rect 8536 38820 8546 38854
rect 8546 38820 8570 38854
rect 8608 38820 8614 38854
rect 8614 38820 8642 38854
rect 8680 38820 8682 38854
rect 8682 38820 8714 38854
rect 8752 38820 8784 38854
rect 8784 38820 8786 38854
rect 8824 38820 8852 38854
rect 8852 38820 8858 38854
rect 8896 38820 8920 38854
rect 8920 38820 8930 38854
rect 8968 38820 8988 38854
rect 8988 38820 9002 38854
rect 9040 38820 9056 38854
rect 9056 38820 9074 38854
rect 9112 38820 9124 38854
rect 9124 38820 9146 38854
rect 9184 38820 9192 38854
rect 9192 38820 9218 38854
rect 9256 38820 9260 38854
rect 9260 38820 9290 38854
rect 9328 38820 9362 38854
rect 9400 38820 9430 38854
rect 9430 38820 9434 38854
rect 9472 38820 9498 38854
rect 9498 38820 9506 38854
rect 9544 38820 9566 38854
rect 9566 38820 9578 38854
rect 9616 38820 9634 38854
rect 9634 38820 9650 38854
rect 9688 38820 9702 38854
rect 9702 38820 9722 38854
rect 9760 38820 9770 38854
rect 9770 38820 9794 38854
rect 9832 38820 9838 38854
rect 9838 38820 9866 38854
rect 9904 38820 9906 38854
rect 9906 38820 9938 38854
rect 9976 38820 10008 38854
rect 10008 38820 10010 38854
rect 10048 38820 10076 38854
rect 10076 38820 10082 38854
rect 10120 38820 10144 38854
rect 10144 38820 10154 38854
rect 10192 38820 10212 38854
rect 10212 38820 10226 38854
rect 10264 38820 10280 38854
rect 10280 38820 10298 38854
rect 10336 38820 10348 38854
rect 10348 38820 10370 38854
rect 10408 38820 10416 38854
rect 10416 38820 10442 38854
rect 10480 38820 10484 38854
rect 10484 38820 10514 38854
rect 10552 38820 10586 38854
rect 10624 38820 10654 38854
rect 10654 38820 10658 38854
rect 10696 38820 10722 38854
rect 10722 38820 10730 38854
rect 10768 38820 10790 38854
rect 10790 38820 10802 38854
rect 10840 38820 10858 38854
rect 10858 38820 10874 38854
rect 10912 38820 10926 38854
rect 10926 38820 10946 38854
rect 10984 38820 10994 38854
rect 10994 38820 11018 38854
rect 11056 38820 11062 38854
rect 11062 38820 11090 38854
rect 11128 38820 11130 38854
rect 11130 38820 11162 38854
rect 11200 38820 11232 38854
rect 11232 38820 11234 38854
rect 11272 38820 11300 38854
rect 11300 38820 11306 38854
rect 11344 38820 11368 38854
rect 11368 38820 11378 38854
rect 11416 38820 11436 38854
rect 11436 38820 11450 38854
rect 11488 38820 11504 38854
rect 11504 38820 11522 38854
rect 11560 38820 11572 38854
rect 11572 38820 11594 38854
rect 11632 38820 11640 38854
rect 11640 38820 11666 38854
rect 11704 38820 11708 38854
rect 11708 38820 11738 38854
rect 11776 38820 11810 38854
rect 11848 38820 11878 38854
rect 11878 38820 11882 38854
rect 11920 38820 11946 38854
rect 11946 38820 11954 38854
rect 11992 38820 12014 38854
rect 12014 38820 12026 38854
rect 12064 38820 12082 38854
rect 12082 38820 12098 38854
rect 12136 38820 12150 38854
rect 12150 38820 12170 38854
rect 12208 38820 12218 38854
rect 12218 38820 12242 38854
rect 12280 38820 12286 38854
rect 12286 38820 12314 38854
rect 12352 38820 12354 38854
rect 12354 38820 12386 38854
rect 12424 38820 12456 38854
rect 12456 38820 12458 38854
rect 12496 38820 12524 38854
rect 12524 38820 12530 38854
rect 12568 38820 12592 38854
rect 12592 38820 12602 38854
rect 12640 38820 12660 38854
rect 12660 38820 12674 38854
rect 12712 38820 12728 38854
rect 12728 38820 12746 38854
rect 12784 38820 12796 38854
rect 12796 38820 12818 38854
rect 12856 38820 12864 38854
rect 12864 38820 12890 38854
rect 12928 38820 12932 38854
rect 12932 38820 12962 38854
rect 13000 38820 13034 38854
rect 13072 38820 13102 38854
rect 13102 38820 13106 38854
rect 2219 38773 2253 38807
rect 2291 38773 2325 38807
rect 2363 38774 2397 38808
rect 2219 38700 2253 38734
rect 2291 38700 2325 38734
rect 2363 38701 2397 38735
rect 2219 38627 2253 38661
rect 2291 38627 2325 38661
rect 2363 38628 2397 38662
rect 2219 38554 2253 38588
rect 2291 38554 2325 38588
rect 2363 38555 2397 38589
rect 2219 38481 2253 38515
rect 2291 38481 2325 38515
rect 2363 38482 2397 38516
rect 2219 38408 2253 38442
rect 2291 38408 2325 38442
rect 2363 38409 2397 38443
rect 2219 38335 2253 38369
rect 2291 38335 2325 38369
rect 2363 38336 2397 38370
rect 2219 38262 2253 38296
rect 2291 38262 2325 38296
rect 2363 38263 2397 38297
rect 2219 38189 2253 38223
rect 2291 38189 2325 38223
rect 2363 38190 2397 38224
rect 2219 38116 2253 38150
rect 2291 38116 2325 38150
rect 2363 38117 2397 38151
rect 2219 38043 2253 38077
rect 2291 38043 2325 38077
rect 2363 38044 2397 38078
rect 2219 37970 2253 38004
rect 2291 37970 2325 38004
rect 2363 37971 2397 38005
rect 2219 37897 2253 37931
rect 2291 37897 2325 37931
rect 2363 37898 2397 37932
rect 2219 37824 2253 37858
rect 2291 37824 2325 37858
rect 2363 37825 2397 37859
rect 2219 37751 2253 37785
rect 2291 37751 2325 37785
rect 2363 37752 2397 37786
rect 2219 37678 2253 37712
rect 2291 37678 2325 37712
rect 2363 37679 2397 37713
rect 2219 37605 2253 37639
rect 2291 37605 2325 37639
rect 2363 37606 2397 37640
rect 2219 37532 2253 37566
rect 2291 37532 2325 37566
rect 2363 37533 2397 37567
rect 2219 37459 2253 37493
rect 2291 37459 2325 37493
rect 2363 37460 2397 37494
rect 2219 37386 2253 37420
rect 2291 37386 2325 37420
rect 2363 37387 2397 37421
rect 2679 38680 2713 38714
rect 2751 38680 2785 38714
rect 2679 38607 2713 38641
rect 2751 38607 2785 38641
rect 2679 38534 2713 38568
rect 2751 38534 2785 38568
rect 2679 38461 2713 38495
rect 2751 38461 2785 38495
rect 2679 37380 2785 38422
rect 2956 38680 2990 38714
rect 3028 38680 3062 38714
rect 2956 38607 2990 38641
rect 3028 38607 3062 38641
rect 2956 38534 2990 38568
rect 3028 38534 3062 38568
rect 2956 38461 2990 38495
rect 3028 38461 3062 38495
rect 2956 37380 3062 38422
rect 3233 38680 3267 38714
rect 3305 38680 3339 38714
rect 3233 38607 3267 38641
rect 3305 38607 3339 38641
rect 3233 38534 3267 38568
rect 3305 38534 3339 38568
rect 3233 38461 3267 38495
rect 3305 38461 3339 38495
rect 3233 37380 3339 38422
rect 3510 38680 3544 38714
rect 3582 38680 3616 38714
rect 3510 38607 3544 38641
rect 3582 38607 3616 38641
rect 3510 38534 3544 38568
rect 3582 38534 3616 38568
rect 3510 38461 3544 38495
rect 3582 38461 3616 38495
rect 3510 37380 3616 38422
rect 3787 38680 3821 38714
rect 3859 38680 3893 38714
rect 3787 38607 3821 38641
rect 3859 38607 3893 38641
rect 3787 38534 3821 38568
rect 3859 38534 3893 38568
rect 3787 38461 3821 38495
rect 3859 38461 3893 38495
rect 3787 37380 3893 38422
rect 4064 38680 4098 38714
rect 4136 38680 4170 38714
rect 4064 38607 4098 38641
rect 4136 38607 4170 38641
rect 4064 38534 4098 38568
rect 4136 38534 4170 38568
rect 4064 38461 4098 38495
rect 4136 38461 4170 38495
rect 4064 37380 4170 38422
rect 4341 38680 4375 38714
rect 4413 38680 4447 38714
rect 4341 38607 4375 38641
rect 4413 38607 4447 38641
rect 4341 38534 4375 38568
rect 4413 38534 4447 38568
rect 4341 38461 4375 38495
rect 4413 38461 4447 38495
rect 4341 37380 4447 38422
rect 4618 38680 4652 38714
rect 4690 38680 4724 38714
rect 4618 38607 4652 38641
rect 4690 38607 4724 38641
rect 4618 38534 4652 38568
rect 4690 38534 4724 38568
rect 4618 38461 4652 38495
rect 4690 38461 4724 38495
rect 4618 37380 4724 38422
rect 4895 38680 4929 38714
rect 4967 38680 5001 38714
rect 4895 38607 4929 38641
rect 4967 38607 5001 38641
rect 4895 38534 4929 38568
rect 4967 38534 5001 38568
rect 4895 38461 4929 38495
rect 4967 38461 5001 38495
rect 4895 37380 5001 38422
rect 5172 38680 5206 38714
rect 5244 38680 5278 38714
rect 5172 38607 5206 38641
rect 5244 38607 5278 38641
rect 5172 38534 5206 38568
rect 5244 38534 5278 38568
rect 5172 38461 5206 38495
rect 5244 38461 5278 38495
rect 5172 37380 5278 38422
rect 5449 38680 5483 38714
rect 5521 38680 5555 38714
rect 5449 38607 5483 38641
rect 5521 38607 5555 38641
rect 5449 38534 5483 38568
rect 5521 38534 5555 38568
rect 5449 38461 5483 38495
rect 5521 38461 5555 38495
rect 5449 37380 5555 38422
rect 5726 38680 5760 38714
rect 5798 38680 5832 38714
rect 5726 38607 5760 38641
rect 5798 38607 5832 38641
rect 5726 38534 5760 38568
rect 5798 38534 5832 38568
rect 5726 38461 5760 38495
rect 5798 38461 5832 38495
rect 5726 37380 5832 38422
rect 6003 38680 6037 38714
rect 6075 38680 6109 38714
rect 6003 38607 6037 38641
rect 6075 38607 6109 38641
rect 6003 38534 6037 38568
rect 6075 38534 6109 38568
rect 6003 38461 6037 38495
rect 6075 38461 6109 38495
rect 6003 37380 6109 38422
rect 6280 38680 6314 38714
rect 6352 38680 6386 38714
rect 6280 38607 6314 38641
rect 6352 38607 6386 38641
rect 6280 38534 6314 38568
rect 6352 38534 6386 38568
rect 6280 38461 6314 38495
rect 6352 38461 6386 38495
rect 6280 37380 6386 38422
rect 6557 38680 6591 38714
rect 6629 38680 6663 38714
rect 6557 38607 6591 38641
rect 6629 38607 6663 38641
rect 6557 38534 6591 38568
rect 6629 38534 6663 38568
rect 6557 38461 6591 38495
rect 6629 38461 6663 38495
rect 6557 37380 6663 38422
rect 6834 38680 6868 38714
rect 6906 38680 6940 38714
rect 6834 38607 6868 38641
rect 6906 38607 6940 38641
rect 6834 38534 6868 38568
rect 6906 38534 6940 38568
rect 6834 38461 6868 38495
rect 6906 38461 6940 38495
rect 6834 37380 6940 38422
rect 7111 38680 7145 38714
rect 7183 38680 7217 38714
rect 7111 38607 7145 38641
rect 7183 38607 7217 38641
rect 7111 38534 7145 38568
rect 7183 38534 7217 38568
rect 7111 38461 7145 38495
rect 7183 38461 7217 38495
rect 7111 37380 7217 38422
rect 7388 38680 7422 38714
rect 7460 38680 7494 38714
rect 7388 38607 7422 38641
rect 7460 38607 7494 38641
rect 7388 38534 7422 38568
rect 7460 38534 7494 38568
rect 7388 38461 7422 38495
rect 7460 38461 7494 38495
rect 7388 37380 7494 38422
rect 7665 38680 7699 38714
rect 7737 38680 7771 38714
rect 7665 38607 7699 38641
rect 7737 38607 7771 38641
rect 7665 38534 7699 38568
rect 7737 38534 7771 38568
rect 7665 38461 7699 38495
rect 7737 38461 7771 38495
rect 7665 37380 7771 38422
rect 7942 38680 7976 38714
rect 8014 38680 8048 38714
rect 7942 38607 7976 38641
rect 8014 38607 8048 38641
rect 7942 38534 7976 38568
rect 8014 38534 8048 38568
rect 7942 38461 7976 38495
rect 8014 38461 8048 38495
rect 7942 37380 8048 38422
rect 8219 38680 8253 38714
rect 8291 38680 8325 38714
rect 8219 38607 8253 38641
rect 8291 38607 8325 38641
rect 8219 38534 8253 38568
rect 8291 38534 8325 38568
rect 8219 38461 8253 38495
rect 8291 38461 8325 38495
rect 8219 37380 8325 38422
rect 8496 38680 8530 38714
rect 8568 38680 8602 38714
rect 8496 38607 8530 38641
rect 8568 38607 8602 38641
rect 8496 38534 8530 38568
rect 8568 38534 8602 38568
rect 8496 38461 8530 38495
rect 8568 38461 8602 38495
rect 8496 37380 8602 38422
rect 8773 38680 8807 38714
rect 8845 38680 8879 38714
rect 8773 38607 8807 38641
rect 8845 38607 8879 38641
rect 8773 38534 8807 38568
rect 8845 38534 8879 38568
rect 8773 38461 8807 38495
rect 8845 38461 8879 38495
rect 8773 37380 8879 38422
rect 9050 38680 9084 38714
rect 9122 38680 9156 38714
rect 9050 38607 9084 38641
rect 9122 38607 9156 38641
rect 9050 38534 9084 38568
rect 9122 38534 9156 38568
rect 9050 38461 9084 38495
rect 9122 38461 9156 38495
rect 9050 37380 9156 38422
rect 9327 38680 9361 38714
rect 9399 38680 9433 38714
rect 9327 38607 9361 38641
rect 9399 38607 9433 38641
rect 9327 38534 9361 38568
rect 9399 38534 9433 38568
rect 9327 38461 9361 38495
rect 9399 38461 9433 38495
rect 9327 37380 9433 38422
rect 9604 38680 9638 38714
rect 9676 38680 9710 38714
rect 9604 38607 9638 38641
rect 9676 38607 9710 38641
rect 9604 38534 9638 38568
rect 9676 38534 9710 38568
rect 9604 38461 9638 38495
rect 9676 38461 9710 38495
rect 9604 37380 9710 38422
rect 9881 38680 9915 38714
rect 9953 38680 9987 38714
rect 9881 38607 9915 38641
rect 9953 38607 9987 38641
rect 9881 38534 9915 38568
rect 9953 38534 9987 38568
rect 9881 38461 9915 38495
rect 9953 38461 9987 38495
rect 9881 37380 9987 38422
rect 10158 38680 10192 38714
rect 10230 38680 10264 38714
rect 10158 38607 10192 38641
rect 10230 38607 10264 38641
rect 10158 38534 10192 38568
rect 10230 38534 10264 38568
rect 10158 38461 10192 38495
rect 10230 38461 10264 38495
rect 10158 37380 10264 38422
rect 10435 38680 10469 38714
rect 10507 38680 10541 38714
rect 10435 38607 10469 38641
rect 10507 38607 10541 38641
rect 10435 38534 10469 38568
rect 10507 38534 10541 38568
rect 10435 38461 10469 38495
rect 10507 38461 10541 38495
rect 10435 37380 10541 38422
rect 10712 38680 10746 38714
rect 10784 38680 10818 38714
rect 10712 38607 10746 38641
rect 10784 38607 10818 38641
rect 10712 38534 10746 38568
rect 10784 38534 10818 38568
rect 10712 38461 10746 38495
rect 10784 38461 10818 38495
rect 10712 37380 10818 38422
rect 10989 38680 11023 38714
rect 11061 38680 11095 38714
rect 10989 38607 11023 38641
rect 11061 38607 11095 38641
rect 10989 38534 11023 38568
rect 11061 38534 11095 38568
rect 10989 38461 11023 38495
rect 11061 38461 11095 38495
rect 10989 37380 11095 38422
rect 11266 38680 11300 38714
rect 11338 38680 11372 38714
rect 11266 38607 11300 38641
rect 11338 38607 11372 38641
rect 11266 38534 11300 38568
rect 11338 38534 11372 38568
rect 11266 38461 11300 38495
rect 11338 38461 11372 38495
rect 11266 37380 11372 38422
rect 11543 38680 11577 38714
rect 11615 38680 11649 38714
rect 11543 38607 11577 38641
rect 11615 38607 11649 38641
rect 11543 38534 11577 38568
rect 11615 38534 11649 38568
rect 11543 38461 11577 38495
rect 11615 38461 11649 38495
rect 11543 37380 11649 38422
rect 11820 38680 11854 38714
rect 11892 38680 11926 38714
rect 11820 38607 11854 38641
rect 11892 38607 11926 38641
rect 11820 38534 11854 38568
rect 11892 38534 11926 38568
rect 11820 38461 11854 38495
rect 11892 38461 11926 38495
rect 11820 37380 11926 38422
rect 12097 38680 12131 38714
rect 12169 38680 12203 38714
rect 12097 38607 12131 38641
rect 12169 38607 12203 38641
rect 12097 38534 12131 38568
rect 12169 38534 12203 38568
rect 12097 38461 12131 38495
rect 12169 38461 12203 38495
rect 12097 37380 12203 38422
rect 12374 38680 12408 38714
rect 12446 38680 12480 38714
rect 12374 38607 12408 38641
rect 12446 38607 12480 38641
rect 12374 38534 12408 38568
rect 12446 38534 12480 38568
rect 12374 38461 12408 38495
rect 12446 38461 12480 38495
rect 12374 37380 12480 38422
rect 12651 38680 12685 38714
rect 12723 38680 12757 38714
rect 12651 38607 12685 38641
rect 12723 38607 12757 38641
rect 12651 38534 12685 38568
rect 12723 38534 12757 38568
rect 12651 38461 12685 38495
rect 12723 38461 12757 38495
rect 12651 37380 12757 38422
rect 12928 38680 12962 38714
rect 13000 38680 13034 38714
rect 12928 38607 12962 38641
rect 13000 38607 13034 38641
rect 12928 38534 12962 38568
rect 13000 38534 13034 38568
rect 12928 38461 12962 38495
rect 13000 38461 13034 38495
rect 12928 37380 13034 38422
rect 13205 38680 13239 38714
rect 13277 38680 13311 38714
rect 13205 38607 13239 38641
rect 13277 38607 13311 38641
rect 13205 38534 13239 38568
rect 13277 38534 13311 38568
rect 13205 38461 13239 38495
rect 13277 38461 13311 38495
rect 13205 37380 13311 38422
rect 2219 37313 2253 37347
rect 2291 37313 2325 37347
rect 2363 37314 2397 37348
rect 2219 37240 2253 37274
rect 2291 37240 2325 37274
rect 2363 37241 2397 37275
rect 2219 37167 2253 37201
rect 2291 37167 2325 37201
rect 2363 37168 2397 37202
rect 2219 37094 2253 37128
rect 2291 37094 2325 37128
rect 2363 37095 2397 37129
rect 2219 37021 2253 37055
rect 2291 37021 2325 37055
rect 2363 37022 2397 37056
rect 2219 36948 2253 36982
rect 2291 36948 2325 36982
rect 2363 36949 2397 36983
rect 2219 36875 2253 36909
rect 2291 36875 2325 36909
rect 2363 36876 2397 36910
rect 2219 36802 2253 36836
rect 2291 36802 2325 36836
rect 2363 36803 2397 36837
rect 2482 37290 2516 37324
rect 2568 37290 2602 37324
rect 2654 37290 2688 37324
rect 2740 37290 2774 37324
rect 2826 37290 2860 37324
rect 2482 37213 2516 37247
rect 2568 37213 2602 37247
rect 2654 37213 2688 37247
rect 2740 37213 2774 37247
rect 2826 37213 2860 37247
rect 2482 37136 2516 37170
rect 2568 37136 2602 37170
rect 2654 37136 2688 37170
rect 2740 37136 2774 37170
rect 2826 37136 2860 37170
rect 2482 37059 2516 37093
rect 2568 37059 2602 37093
rect 2654 37059 2688 37093
rect 2740 37059 2774 37093
rect 2826 37059 2860 37093
rect 2482 36982 2516 37016
rect 2568 36982 2602 37016
rect 2654 36982 2688 37016
rect 2740 36982 2774 37016
rect 2826 36982 2860 37016
rect 2482 36905 2516 36939
rect 2568 36905 2602 36939
rect 2654 36905 2688 36939
rect 2740 36905 2774 36939
rect 2826 36905 2860 36939
rect 2482 36828 2516 36862
rect 2568 36828 2602 36862
rect 2654 36828 2688 36862
rect 2740 36828 2774 36862
rect 2826 36828 2860 36862
rect 2219 36729 2253 36763
rect 2291 36729 2325 36763
rect 2363 36730 2397 36764
rect 2219 36656 2253 36690
rect 2291 36656 2325 36690
rect 2363 36657 2397 36691
rect 2219 36583 2253 36617
rect 2291 36583 2325 36617
rect 2363 36584 2397 36618
rect 2219 36510 2253 36544
rect 2291 36510 2325 36544
rect 2363 36511 2397 36545
rect 2219 36437 2253 36471
rect 2291 36437 2325 36471
rect 2363 36438 2397 36472
rect 2219 36364 2253 36398
rect 2291 36364 2325 36398
rect 2363 36365 2397 36399
rect 2219 36291 2253 36325
rect 2291 36291 2325 36325
rect 2363 36292 2397 36326
rect 2219 36218 2253 36252
rect 2291 36218 2325 36252
rect 2363 36219 2397 36253
rect 2219 36145 2253 36179
rect 2291 36145 2325 36179
rect 2363 36146 2397 36180
rect 2219 36072 2253 36106
rect 2291 36072 2325 36106
rect 2363 36073 2397 36107
rect 2219 35999 2253 36033
rect 2291 35999 2325 36033
rect 2363 36000 2397 36034
rect 2219 35926 2253 35960
rect 2291 35926 2325 35960
rect 2363 35927 2397 35961
rect 2219 35853 2253 35887
rect 2291 35853 2325 35887
rect 2363 35854 2397 35888
rect 2219 35780 2253 35814
rect 2291 35780 2325 35814
rect 2363 35781 2397 35815
rect 2219 35707 2253 35741
rect 2291 35707 2325 35741
rect 2363 35708 2397 35742
rect 2219 35634 2253 35668
rect 2291 35634 2325 35668
rect 2363 35635 2397 35669
rect 2219 35561 2253 35595
rect 2291 35561 2325 35595
rect 2363 35562 2397 35596
rect 2219 33688 2274 35522
rect 2274 35450 2325 35522
rect 2363 35489 2397 35523
rect 2274 33688 2397 35450
rect 3233 36680 3267 36714
rect 3305 36680 3339 36714
rect 3233 36607 3267 36641
rect 3305 36607 3339 36641
rect 3233 36534 3267 36568
rect 3305 36534 3339 36568
rect 3233 36461 3267 36495
rect 3305 36461 3339 36495
rect 3233 35380 3339 36422
rect 3510 36680 3544 36714
rect 3582 36680 3616 36714
rect 3510 36607 3544 36641
rect 3582 36607 3616 36641
rect 3510 36534 3544 36568
rect 3582 36534 3616 36568
rect 3510 36461 3544 36495
rect 3582 36461 3616 36495
rect 3510 35380 3616 36422
rect 3787 36680 3821 36714
rect 3859 36680 3893 36714
rect 3787 36607 3821 36641
rect 3859 36607 3893 36641
rect 3787 36534 3821 36568
rect 3859 36534 3893 36568
rect 3787 36461 3821 36495
rect 3859 36461 3893 36495
rect 3787 35380 3893 36422
rect 4064 36680 4098 36714
rect 4136 36680 4170 36714
rect 4064 36607 4098 36641
rect 4136 36607 4170 36641
rect 4064 36534 4098 36568
rect 4136 36534 4170 36568
rect 4064 36461 4098 36495
rect 4136 36461 4170 36495
rect 4064 35380 4170 36422
rect 4341 36680 4375 36714
rect 4413 36680 4447 36714
rect 4341 36607 4375 36641
rect 4413 36607 4447 36641
rect 4341 36534 4375 36568
rect 4413 36534 4447 36568
rect 4341 36461 4375 36495
rect 4413 36461 4447 36495
rect 4341 35380 4447 36422
rect 4618 36680 4652 36714
rect 4690 36680 4724 36714
rect 4618 36607 4652 36641
rect 4690 36607 4724 36641
rect 4618 36534 4652 36568
rect 4690 36534 4724 36568
rect 4618 36461 4652 36495
rect 4690 36461 4724 36495
rect 4618 35380 4724 36422
rect 4895 36680 4929 36714
rect 4967 36680 5001 36714
rect 4895 36607 4929 36641
rect 4967 36607 5001 36641
rect 4895 36534 4929 36568
rect 4967 36534 5001 36568
rect 4895 36461 4929 36495
rect 4967 36461 5001 36495
rect 4895 35380 5001 36422
rect 5172 36680 5206 36714
rect 5244 36680 5278 36714
rect 5172 36607 5206 36641
rect 5244 36607 5278 36641
rect 5172 36534 5206 36568
rect 5244 36534 5278 36568
rect 5172 36461 5206 36495
rect 5244 36461 5278 36495
rect 5172 35380 5278 36422
rect 5449 36680 5483 36714
rect 5521 36680 5555 36714
rect 5449 36607 5483 36641
rect 5521 36607 5555 36641
rect 5449 36534 5483 36568
rect 5521 36534 5555 36568
rect 5449 36461 5483 36495
rect 5521 36461 5555 36495
rect 5449 35380 5555 36422
rect 5726 36680 5760 36714
rect 5798 36680 5832 36714
rect 5726 36607 5760 36641
rect 5798 36607 5832 36641
rect 5726 36534 5760 36568
rect 5798 36534 5832 36568
rect 5726 36461 5760 36495
rect 5798 36461 5832 36495
rect 5726 35380 5832 36422
rect 6003 36680 6037 36714
rect 6075 36680 6109 36714
rect 6003 36607 6037 36641
rect 6075 36607 6109 36641
rect 6003 36534 6037 36568
rect 6075 36534 6109 36568
rect 6003 36461 6037 36495
rect 6075 36461 6109 36495
rect 6003 35380 6109 36422
rect 6280 36680 6314 36714
rect 6352 36680 6386 36714
rect 6280 36607 6314 36641
rect 6352 36607 6386 36641
rect 6280 36534 6314 36568
rect 6352 36534 6386 36568
rect 6280 36461 6314 36495
rect 6352 36461 6386 36495
rect 6280 35380 6386 36422
rect 6557 36680 6591 36714
rect 6629 36680 6663 36714
rect 6557 36607 6591 36641
rect 6629 36607 6663 36641
rect 6557 36534 6591 36568
rect 6629 36534 6663 36568
rect 6557 36461 6591 36495
rect 6629 36461 6663 36495
rect 6557 35380 6663 36422
rect 6834 36680 6868 36714
rect 6906 36680 6940 36714
rect 6834 36607 6868 36641
rect 6906 36607 6940 36641
rect 6834 36534 6868 36568
rect 6906 36534 6940 36568
rect 6834 36461 6868 36495
rect 6906 36461 6940 36495
rect 6834 35380 6940 36422
rect 7111 36680 7145 36714
rect 7183 36680 7217 36714
rect 7111 36607 7145 36641
rect 7183 36607 7217 36641
rect 7111 36534 7145 36568
rect 7183 36534 7217 36568
rect 7111 36461 7145 36495
rect 7183 36461 7217 36495
rect 7111 35380 7217 36422
rect 7388 36680 7422 36714
rect 7460 36680 7494 36714
rect 7388 36607 7422 36641
rect 7460 36607 7494 36641
rect 7388 36534 7422 36568
rect 7460 36534 7494 36568
rect 7388 36461 7422 36495
rect 7460 36461 7494 36495
rect 7388 35380 7494 36422
rect 7665 36680 7699 36714
rect 7737 36680 7771 36714
rect 7665 36607 7699 36641
rect 7737 36607 7771 36641
rect 7665 36534 7699 36568
rect 7737 36534 7771 36568
rect 7665 36461 7699 36495
rect 7737 36461 7771 36495
rect 7665 35380 7771 36422
rect 7942 36680 7976 36714
rect 8014 36680 8048 36714
rect 7942 36607 7976 36641
rect 8014 36607 8048 36641
rect 7942 36534 7976 36568
rect 8014 36534 8048 36568
rect 7942 36461 7976 36495
rect 8014 36461 8048 36495
rect 7942 35380 8048 36422
rect 8219 36680 8253 36714
rect 8291 36680 8325 36714
rect 8219 36607 8253 36641
rect 8291 36607 8325 36641
rect 8219 36534 8253 36568
rect 8291 36534 8325 36568
rect 8219 36461 8253 36495
rect 8291 36461 8325 36495
rect 8219 35380 8325 36422
rect 8496 36680 8530 36714
rect 8568 36680 8602 36714
rect 8496 36607 8530 36641
rect 8568 36607 8602 36641
rect 8496 36534 8530 36568
rect 8568 36534 8602 36568
rect 8496 36461 8530 36495
rect 8568 36461 8602 36495
rect 8496 35380 8602 36422
rect 8773 36680 8807 36714
rect 8845 36680 8879 36714
rect 8773 36607 8807 36641
rect 8845 36607 8879 36641
rect 8773 36534 8807 36568
rect 8845 36534 8879 36568
rect 8773 36461 8807 36495
rect 8845 36461 8879 36495
rect 8773 35380 8879 36422
rect 9050 36680 9084 36714
rect 9122 36680 9156 36714
rect 9050 36607 9084 36641
rect 9122 36607 9156 36641
rect 9050 36534 9084 36568
rect 9122 36534 9156 36568
rect 9050 36461 9084 36495
rect 9122 36461 9156 36495
rect 9050 35380 9156 36422
rect 9327 36680 9361 36714
rect 9399 36680 9433 36714
rect 9327 36607 9361 36641
rect 9399 36607 9433 36641
rect 9327 36534 9361 36568
rect 9399 36534 9433 36568
rect 9327 36461 9361 36495
rect 9399 36461 9433 36495
rect 9327 35380 9433 36422
rect 9604 36680 9638 36714
rect 9676 36680 9710 36714
rect 9604 36607 9638 36641
rect 9676 36607 9710 36641
rect 9604 36534 9638 36568
rect 9676 36534 9710 36568
rect 9604 36461 9638 36495
rect 9676 36461 9710 36495
rect 9604 35380 9710 36422
rect 9881 36680 9915 36714
rect 9953 36680 9987 36714
rect 9881 36607 9915 36641
rect 9953 36607 9987 36641
rect 9881 36534 9915 36568
rect 9953 36534 9987 36568
rect 9881 36461 9915 36495
rect 9953 36461 9987 36495
rect 9881 35380 9987 36422
rect 10158 36680 10192 36714
rect 10230 36680 10264 36714
rect 10158 36607 10192 36641
rect 10230 36607 10264 36641
rect 10158 36534 10192 36568
rect 10230 36534 10264 36568
rect 10158 36461 10192 36495
rect 10230 36461 10264 36495
rect 10158 35380 10264 36422
rect 10435 36680 10469 36714
rect 10507 36680 10541 36714
rect 10435 36607 10469 36641
rect 10507 36607 10541 36641
rect 10435 36534 10469 36568
rect 10507 36534 10541 36568
rect 10435 36461 10469 36495
rect 10507 36461 10541 36495
rect 10435 35380 10541 36422
rect 10712 36680 10746 36714
rect 10784 36680 10818 36714
rect 10712 36607 10746 36641
rect 10784 36607 10818 36641
rect 10712 36534 10746 36568
rect 10784 36534 10818 36568
rect 10712 36461 10746 36495
rect 10784 36461 10818 36495
rect 10712 35380 10818 36422
rect 10989 36680 11023 36714
rect 11061 36680 11095 36714
rect 10989 36607 11023 36641
rect 11061 36607 11095 36641
rect 10989 36534 11023 36568
rect 11061 36534 11095 36568
rect 10989 36461 11023 36495
rect 11061 36461 11095 36495
rect 10989 35380 11095 36422
rect 11266 36680 11300 36714
rect 11338 36680 11372 36714
rect 11266 36607 11300 36641
rect 11338 36607 11372 36641
rect 11266 36534 11300 36568
rect 11338 36534 11372 36568
rect 11266 36461 11300 36495
rect 11338 36461 11372 36495
rect 11266 35380 11372 36422
rect 11543 36680 11577 36714
rect 11615 36680 11649 36714
rect 11543 36607 11577 36641
rect 11615 36607 11649 36641
rect 11543 36534 11577 36568
rect 11615 36534 11649 36568
rect 11543 36461 11577 36495
rect 11615 36461 11649 36495
rect 11543 35380 11649 36422
rect 11820 36680 11854 36714
rect 11892 36680 11926 36714
rect 11820 36607 11854 36641
rect 11892 36607 11926 36641
rect 11820 36534 11854 36568
rect 11892 36534 11926 36568
rect 11820 36461 11854 36495
rect 11892 36461 11926 36495
rect 11820 35380 11926 36422
rect 12097 36680 12131 36714
rect 12169 36680 12203 36714
rect 12097 36607 12131 36641
rect 12169 36607 12203 36641
rect 12097 36534 12131 36568
rect 12169 36534 12203 36568
rect 12097 36461 12131 36495
rect 12169 36461 12203 36495
rect 12097 35380 12203 36422
rect 12374 36680 12408 36714
rect 12446 36680 12480 36714
rect 12374 36607 12408 36641
rect 12446 36607 12480 36641
rect 12374 36534 12408 36568
rect 12446 36534 12480 36568
rect 12374 36461 12408 36495
rect 12446 36461 12480 36495
rect 12374 35380 12480 36422
rect 12651 36680 12685 36714
rect 12723 36680 12757 36714
rect 12651 36607 12685 36641
rect 12723 36607 12757 36641
rect 12651 36534 12685 36568
rect 12723 36534 12757 36568
rect 12651 36461 12685 36495
rect 12723 36461 12757 36495
rect 12651 35380 12757 36422
rect 12928 36680 12962 36714
rect 13000 36680 13034 36714
rect 12928 36607 12962 36641
rect 13000 36607 13034 36641
rect 12928 36534 12962 36568
rect 13000 36534 13034 36568
rect 12928 36461 12962 36495
rect 13000 36461 13034 36495
rect 12928 35380 13034 36422
rect 13205 36680 13239 36714
rect 13277 36680 13311 36714
rect 13205 36607 13239 36641
rect 13277 36607 13311 36641
rect 13205 36534 13239 36568
rect 13277 36534 13311 36568
rect 13205 36461 13239 36495
rect 13277 36461 13311 36495
rect 13205 35380 13311 36422
rect 2674 35287 2708 35321
rect 2750 35287 2784 35321
rect 2826 35287 2860 35321
rect 2674 35210 2708 35244
rect 2750 35210 2784 35244
rect 2826 35210 2860 35244
rect 2674 35133 2708 35167
rect 2750 35133 2784 35167
rect 2826 35133 2860 35167
rect 2674 35055 2708 35089
rect 2750 35055 2784 35089
rect 2826 35055 2860 35089
rect 2674 34977 2708 35011
rect 2750 34977 2784 35011
rect 2826 34977 2860 35011
rect 2674 34899 2708 34933
rect 2750 34899 2784 34933
rect 2826 34899 2860 34933
rect 2674 34821 2708 34855
rect 2750 34821 2784 34855
rect 2826 34821 2860 34855
rect 2219 33610 2253 33644
rect 2325 33610 2359 33644
rect 2219 33537 2253 33571
rect 2325 33537 2359 33571
rect 2219 33464 2253 33498
rect 2325 33464 2359 33498
rect 2219 33391 2253 33425
rect 2325 33391 2359 33425
rect 3173 34680 3207 34714
rect 3245 34680 3279 34714
rect 3173 34607 3207 34641
rect 3245 34607 3279 34641
rect 3173 34534 3207 34568
rect 3245 34534 3279 34568
rect 3173 34461 3207 34495
rect 3245 34461 3279 34495
rect 3173 33380 3279 34422
rect 3591 34680 3625 34714
rect 3663 34680 3697 34714
rect 3591 34607 3625 34641
rect 3663 34607 3697 34641
rect 3591 34534 3625 34568
rect 3663 34534 3697 34568
rect 3591 34461 3625 34495
rect 3663 34461 3697 34495
rect 3591 33380 3697 34422
rect 4009 34680 4043 34714
rect 4081 34680 4115 34714
rect 4009 34607 4043 34641
rect 4081 34607 4115 34641
rect 4009 34534 4043 34568
rect 4081 34534 4115 34568
rect 4009 34461 4043 34495
rect 4081 34461 4115 34495
rect 4009 33380 4115 34422
rect 4427 34680 4461 34714
rect 4499 34680 4533 34714
rect 4427 34607 4461 34641
rect 4499 34607 4533 34641
rect 4427 34534 4461 34568
rect 4499 34534 4533 34568
rect 4427 34461 4461 34495
rect 4499 34461 4533 34495
rect 4427 33380 4533 34422
rect 4845 34680 4879 34714
rect 4917 34680 4951 34714
rect 4845 34607 4879 34641
rect 4917 34607 4951 34641
rect 4845 34534 4879 34568
rect 4917 34534 4951 34568
rect 4845 34461 4879 34495
rect 4917 34461 4951 34495
rect 4845 33380 4951 34422
rect 5263 34680 5297 34714
rect 5335 34680 5369 34714
rect 5263 34607 5297 34641
rect 5335 34607 5369 34641
rect 5263 34534 5297 34568
rect 5335 34534 5369 34568
rect 5263 34461 5297 34495
rect 5335 34461 5369 34495
rect 5263 33380 5369 34422
rect 5681 34680 5715 34714
rect 5753 34680 5787 34714
rect 5681 34607 5715 34641
rect 5753 34607 5787 34641
rect 5681 34534 5715 34568
rect 5753 34534 5787 34568
rect 5681 34461 5715 34495
rect 5753 34461 5787 34495
rect 5681 33380 5787 34422
rect 6099 34680 6133 34714
rect 6171 34680 6205 34714
rect 6099 34607 6133 34641
rect 6171 34607 6205 34641
rect 6099 34534 6133 34568
rect 6171 34534 6205 34568
rect 6099 34461 6133 34495
rect 6171 34461 6205 34495
rect 6099 33380 6205 34422
rect 6517 34680 6551 34714
rect 6589 34680 6623 34714
rect 6517 34607 6551 34641
rect 6589 34607 6623 34641
rect 6517 34534 6551 34568
rect 6589 34534 6623 34568
rect 6517 34461 6551 34495
rect 6589 34461 6623 34495
rect 6517 33380 6623 34422
rect 6935 34680 6969 34714
rect 7007 34680 7041 34714
rect 6935 34607 6969 34641
rect 7007 34607 7041 34641
rect 6935 34534 6969 34568
rect 7007 34534 7041 34568
rect 6935 34461 6969 34495
rect 7007 34461 7041 34495
rect 6935 33380 7041 34422
rect 7353 34680 7387 34714
rect 7425 34680 7459 34714
rect 7353 34607 7387 34641
rect 7425 34607 7459 34641
rect 7353 34534 7387 34568
rect 7425 34534 7459 34568
rect 7353 34461 7387 34495
rect 7425 34461 7459 34495
rect 7353 33380 7459 34422
rect 7771 34680 7805 34714
rect 7843 34680 7877 34714
rect 7771 34607 7805 34641
rect 7843 34607 7877 34641
rect 7771 34534 7805 34568
rect 7843 34534 7877 34568
rect 7771 34461 7805 34495
rect 7843 34461 7877 34495
rect 7771 33380 7877 34422
rect 8189 34680 8223 34714
rect 8261 34680 8295 34714
rect 8189 34607 8223 34641
rect 8261 34607 8295 34641
rect 8189 34534 8223 34568
rect 8261 34534 8295 34568
rect 8189 34461 8223 34495
rect 8261 34461 8295 34495
rect 8189 33380 8295 34422
rect 8607 34680 8641 34714
rect 8679 34680 8713 34714
rect 8607 34607 8641 34641
rect 8679 34607 8713 34641
rect 8607 34534 8641 34568
rect 8679 34534 8713 34568
rect 8607 34461 8641 34495
rect 8679 34461 8713 34495
rect 8607 33380 8713 34422
rect 9025 34680 9059 34714
rect 9097 34680 9131 34714
rect 9025 34607 9059 34641
rect 9097 34607 9131 34641
rect 9025 34534 9059 34568
rect 9097 34534 9131 34568
rect 9025 34461 9059 34495
rect 9097 34461 9131 34495
rect 9025 33380 9131 34422
rect 9443 34680 9477 34714
rect 9515 34680 9549 34714
rect 9443 34607 9477 34641
rect 9515 34607 9549 34641
rect 9443 34534 9477 34568
rect 9515 34534 9549 34568
rect 9443 34461 9477 34495
rect 9515 34461 9549 34495
rect 9443 33380 9549 34422
rect 9861 34680 9895 34714
rect 9933 34680 9967 34714
rect 9861 34607 9895 34641
rect 9933 34607 9967 34641
rect 9861 34534 9895 34568
rect 9933 34534 9967 34568
rect 9861 34461 9895 34495
rect 9933 34461 9967 34495
rect 9861 33380 9967 34422
rect 10279 34680 10313 34714
rect 10351 34680 10385 34714
rect 10279 34607 10313 34641
rect 10351 34607 10385 34641
rect 10279 34534 10313 34568
rect 10351 34534 10385 34568
rect 10279 34461 10313 34495
rect 10351 34461 10385 34495
rect 10279 33380 10385 34422
rect 10697 34680 10731 34714
rect 10769 34680 10803 34714
rect 10697 34607 10731 34641
rect 10769 34607 10803 34641
rect 10697 34534 10731 34568
rect 10769 34534 10803 34568
rect 10697 34461 10731 34495
rect 10769 34461 10803 34495
rect 10697 33380 10803 34422
rect 11115 34680 11149 34714
rect 11187 34680 11221 34714
rect 11115 34607 11149 34641
rect 11187 34607 11221 34641
rect 11115 34534 11149 34568
rect 11187 34534 11221 34568
rect 11115 34461 11149 34495
rect 11187 34461 11221 34495
rect 11115 33380 11221 34422
rect 11533 34680 11567 34714
rect 11605 34680 11639 34714
rect 11533 34607 11567 34641
rect 11605 34607 11639 34641
rect 11533 34534 11567 34568
rect 11605 34534 11639 34568
rect 11533 34461 11567 34495
rect 11605 34461 11639 34495
rect 11533 33380 11639 34422
rect 11951 34680 11985 34714
rect 12023 34680 12057 34714
rect 11951 34607 11985 34641
rect 12023 34607 12057 34641
rect 11951 34534 11985 34568
rect 12023 34534 12057 34568
rect 11951 34461 11985 34495
rect 12023 34461 12057 34495
rect 11951 33380 12057 34422
rect 12369 34680 12403 34714
rect 12441 34680 12475 34714
rect 12369 34607 12403 34641
rect 12441 34607 12475 34641
rect 12369 34534 12403 34568
rect 12441 34534 12475 34568
rect 12369 34461 12403 34495
rect 12441 34461 12475 34495
rect 12369 33380 12475 34422
rect 12787 34680 12821 34714
rect 12859 34680 12893 34714
rect 12787 34607 12821 34641
rect 12859 34607 12893 34641
rect 12787 34534 12821 34568
rect 12859 34534 12893 34568
rect 12787 34461 12821 34495
rect 12859 34461 12893 34495
rect 12787 33380 12893 34422
rect 13205 34680 13239 34714
rect 13277 34680 13311 34714
rect 13205 34607 13239 34641
rect 13277 34607 13311 34641
rect 13205 34534 13239 34568
rect 13277 34534 13311 34568
rect 13205 34461 13239 34495
rect 13277 34461 13311 34495
rect 13205 33380 13311 34422
rect 2219 33318 2253 33352
rect 2325 33318 2359 33352
rect 2219 33245 2253 33279
rect 2325 33245 2359 33279
rect 2219 33172 2253 33206
rect 2325 33172 2359 33206
rect 2219 33099 2253 33133
rect 2325 33099 2359 33133
rect 2219 33026 2253 33060
rect 2325 33026 2359 33060
rect 2219 32953 2253 32987
rect 2325 32953 2359 32987
rect 2219 32880 2253 32914
rect 2325 32880 2359 32914
rect 2219 32807 2253 32841
rect 2325 32807 2359 32841
rect 2674 33288 2708 33322
rect 2750 33288 2784 33322
rect 2826 33288 2860 33322
rect 2674 33211 2708 33245
rect 2750 33211 2784 33245
rect 2826 33211 2860 33245
rect 2674 33134 2708 33168
rect 2750 33134 2784 33168
rect 2826 33134 2860 33168
rect 2674 33056 2708 33090
rect 2750 33056 2784 33090
rect 2826 33056 2860 33090
rect 2674 32978 2708 33012
rect 2750 32978 2784 33012
rect 2826 32978 2860 33012
rect 2674 32900 2708 32934
rect 2750 32900 2784 32934
rect 2826 32900 2860 32934
rect 2674 32822 2708 32856
rect 2750 32822 2784 32856
rect 2826 32822 2860 32856
rect 2219 32734 2253 32768
rect 2325 32734 2359 32768
rect 2219 32661 2253 32695
rect 2325 32661 2359 32695
rect 2219 32588 2253 32622
rect 2325 32588 2359 32622
rect 2219 32515 2253 32549
rect 2325 32515 2359 32549
rect 2219 32442 2253 32476
rect 2325 32442 2359 32476
rect 2219 32369 2253 32403
rect 2325 32369 2359 32403
rect 2219 32296 2253 32330
rect 2325 32296 2359 32330
rect 2219 32223 2253 32257
rect 2325 32223 2359 32257
rect 2219 32150 2253 32184
rect 2325 32150 2359 32184
rect 2219 32077 2253 32111
rect 2325 32077 2359 32111
rect 2219 32004 2253 32038
rect 2325 32004 2359 32038
rect 2219 31931 2253 31965
rect 2325 31931 2359 31965
rect 2219 31858 2253 31892
rect 2325 31858 2359 31892
rect 2219 31785 2253 31819
rect 2325 31785 2359 31819
rect 2219 31712 2253 31746
rect 2325 31712 2359 31746
rect 2219 31639 2253 31673
rect 2325 31639 2359 31673
rect 2219 31566 2253 31600
rect 2325 31566 2359 31600
rect 2219 31493 2253 31527
rect 2325 31493 2359 31527
rect 2219 31420 2253 31454
rect 2325 31420 2359 31454
rect 2219 31347 2253 31381
rect 2325 31347 2359 31381
rect 3173 32680 3207 32714
rect 3245 32680 3279 32714
rect 3173 32607 3207 32641
rect 3245 32607 3279 32641
rect 3173 32534 3207 32568
rect 3245 32534 3279 32568
rect 3173 32461 3207 32495
rect 3245 32461 3279 32495
rect 3173 31380 3279 32422
rect 3591 32680 3625 32714
rect 3663 32680 3697 32714
rect 3591 32607 3625 32641
rect 3663 32607 3697 32641
rect 3591 32534 3625 32568
rect 3663 32534 3697 32568
rect 3591 32461 3625 32495
rect 3663 32461 3697 32495
rect 3591 31380 3697 32422
rect 4009 32680 4043 32714
rect 4081 32680 4115 32714
rect 4009 32607 4043 32641
rect 4081 32607 4115 32641
rect 4009 32534 4043 32568
rect 4081 32534 4115 32568
rect 4009 32461 4043 32495
rect 4081 32461 4115 32495
rect 4009 31380 4115 32422
rect 4427 32680 4461 32714
rect 4499 32680 4533 32714
rect 4427 32607 4461 32641
rect 4499 32607 4533 32641
rect 4427 32534 4461 32568
rect 4499 32534 4533 32568
rect 4427 32461 4461 32495
rect 4499 32461 4533 32495
rect 4427 31380 4533 32422
rect 4845 32680 4879 32714
rect 4917 32680 4951 32714
rect 4845 32607 4879 32641
rect 4917 32607 4951 32641
rect 4845 32534 4879 32568
rect 4917 32534 4951 32568
rect 4845 32461 4879 32495
rect 4917 32461 4951 32495
rect 4845 31380 4951 32422
rect 5263 32680 5297 32714
rect 5335 32680 5369 32714
rect 5263 32607 5297 32641
rect 5335 32607 5369 32641
rect 5263 32534 5297 32568
rect 5335 32534 5369 32568
rect 5263 32461 5297 32495
rect 5335 32461 5369 32495
rect 5263 31380 5369 32422
rect 5681 32680 5715 32714
rect 5753 32680 5787 32714
rect 5681 32607 5715 32641
rect 5753 32607 5787 32641
rect 5681 32534 5715 32568
rect 5753 32534 5787 32568
rect 5681 32461 5715 32495
rect 5753 32461 5787 32495
rect 5681 31380 5787 32422
rect 6099 32680 6133 32714
rect 6171 32680 6205 32714
rect 6099 32607 6133 32641
rect 6171 32607 6205 32641
rect 6099 32534 6133 32568
rect 6171 32534 6205 32568
rect 6099 32461 6133 32495
rect 6171 32461 6205 32495
rect 6099 31380 6205 32422
rect 6517 32680 6551 32714
rect 6589 32680 6623 32714
rect 6517 32607 6551 32641
rect 6589 32607 6623 32641
rect 6517 32534 6551 32568
rect 6589 32534 6623 32568
rect 6517 32461 6551 32495
rect 6589 32461 6623 32495
rect 6517 31380 6623 32422
rect 6935 32680 6969 32714
rect 7007 32680 7041 32714
rect 6935 32607 6969 32641
rect 7007 32607 7041 32641
rect 6935 32534 6969 32568
rect 7007 32534 7041 32568
rect 6935 32461 6969 32495
rect 7007 32461 7041 32495
rect 6935 31380 7041 32422
rect 7353 32680 7387 32714
rect 7425 32680 7459 32714
rect 7353 32607 7387 32641
rect 7425 32607 7459 32641
rect 7353 32534 7387 32568
rect 7425 32534 7459 32568
rect 7353 32461 7387 32495
rect 7425 32461 7459 32495
rect 7353 31380 7459 32422
rect 7771 32680 7805 32714
rect 7843 32680 7877 32714
rect 7771 32607 7805 32641
rect 7843 32607 7877 32641
rect 7771 32534 7805 32568
rect 7843 32534 7877 32568
rect 7771 32461 7805 32495
rect 7843 32461 7877 32495
rect 7771 31380 7877 32422
rect 8189 32680 8223 32714
rect 8261 32680 8295 32714
rect 8189 32607 8223 32641
rect 8261 32607 8295 32641
rect 8189 32534 8223 32568
rect 8261 32534 8295 32568
rect 8189 32461 8223 32495
rect 8261 32461 8295 32495
rect 8189 31380 8295 32422
rect 8607 32680 8641 32714
rect 8679 32680 8713 32714
rect 8607 32607 8641 32641
rect 8679 32607 8713 32641
rect 8607 32534 8641 32568
rect 8679 32534 8713 32568
rect 8607 32461 8641 32495
rect 8679 32461 8713 32495
rect 8607 31380 8713 32422
rect 9025 32680 9059 32714
rect 9097 32680 9131 32714
rect 9025 32607 9059 32641
rect 9097 32607 9131 32641
rect 9025 32534 9059 32568
rect 9097 32534 9131 32568
rect 9025 32461 9059 32495
rect 9097 32461 9131 32495
rect 9025 31380 9131 32422
rect 9443 32680 9477 32714
rect 9515 32680 9549 32714
rect 9443 32607 9477 32641
rect 9515 32607 9549 32641
rect 9443 32534 9477 32568
rect 9515 32534 9549 32568
rect 9443 32461 9477 32495
rect 9515 32461 9549 32495
rect 9443 31380 9549 32422
rect 9861 32680 9895 32714
rect 9933 32680 9967 32714
rect 9861 32607 9895 32641
rect 9933 32607 9967 32641
rect 9861 32534 9895 32568
rect 9933 32534 9967 32568
rect 9861 32461 9895 32495
rect 9933 32461 9967 32495
rect 9861 31380 9967 32422
rect 10279 32680 10313 32714
rect 10351 32680 10385 32714
rect 10279 32607 10313 32641
rect 10351 32607 10385 32641
rect 10279 32534 10313 32568
rect 10351 32534 10385 32568
rect 10279 32461 10313 32495
rect 10351 32461 10385 32495
rect 10279 31380 10385 32422
rect 10697 32680 10731 32714
rect 10769 32680 10803 32714
rect 10697 32607 10731 32641
rect 10769 32607 10803 32641
rect 10697 32534 10731 32568
rect 10769 32534 10803 32568
rect 10697 32461 10731 32495
rect 10769 32461 10803 32495
rect 10697 31380 10803 32422
rect 11115 32680 11149 32714
rect 11187 32680 11221 32714
rect 11115 32607 11149 32641
rect 11187 32607 11221 32641
rect 11115 32534 11149 32568
rect 11187 32534 11221 32568
rect 11115 32461 11149 32495
rect 11187 32461 11221 32495
rect 11115 31380 11221 32422
rect 11533 32680 11567 32714
rect 11605 32680 11639 32714
rect 11533 32607 11567 32641
rect 11605 32607 11639 32641
rect 11533 32534 11567 32568
rect 11605 32534 11639 32568
rect 11533 32461 11567 32495
rect 11605 32461 11639 32495
rect 11533 31380 11639 32422
rect 11951 32680 11985 32714
rect 12023 32680 12057 32714
rect 11951 32607 11985 32641
rect 12023 32607 12057 32641
rect 11951 32534 11985 32568
rect 12023 32534 12057 32568
rect 11951 32461 11985 32495
rect 12023 32461 12057 32495
rect 11951 31380 12057 32422
rect 12369 32680 12403 32714
rect 12441 32680 12475 32714
rect 12369 32607 12403 32641
rect 12441 32607 12475 32641
rect 12369 32534 12403 32568
rect 12441 32534 12475 32568
rect 12369 32461 12403 32495
rect 12441 32461 12475 32495
rect 12369 31380 12475 32422
rect 12787 32680 12821 32714
rect 12859 32680 12893 32714
rect 12787 32607 12821 32641
rect 12859 32607 12893 32641
rect 12787 32534 12821 32568
rect 12859 32534 12893 32568
rect 12787 32461 12821 32495
rect 12859 32461 12893 32495
rect 12787 31380 12893 32422
rect 13205 32680 13239 32714
rect 13277 32680 13311 32714
rect 13205 32607 13239 32641
rect 13277 32607 13311 32641
rect 13205 32534 13239 32568
rect 13277 32534 13311 32568
rect 13205 32461 13239 32495
rect 13277 32461 13311 32495
rect 13205 31380 13311 32422
rect 2219 31274 2253 31308
rect 2325 31274 2359 31308
rect 2219 31201 2253 31235
rect 2325 31201 2359 31235
rect 2219 31128 2253 31162
rect 2325 31128 2359 31162
rect 2219 31055 2253 31089
rect 2325 31055 2359 31089
rect 2219 30982 2253 31016
rect 2325 30982 2359 31016
rect 2219 30909 2253 30943
rect 2325 30909 2359 30943
rect 2219 30837 2253 30871
rect 2325 30837 2359 30871
rect 2674 31289 2708 31323
rect 2750 31289 2784 31323
rect 2826 31289 2860 31323
rect 2674 31212 2708 31246
rect 2750 31212 2784 31246
rect 2826 31212 2860 31246
rect 2674 31135 2708 31169
rect 2750 31135 2784 31169
rect 2826 31135 2860 31169
rect 2674 31057 2708 31091
rect 2750 31057 2784 31091
rect 2826 31057 2860 31091
rect 2674 30979 2708 31013
rect 2750 30979 2784 31013
rect 2826 30979 2860 31013
rect 2674 30901 2708 30935
rect 2750 30901 2784 30935
rect 2826 30901 2860 30935
rect 2674 30823 2708 30857
rect 2750 30823 2784 30857
rect 2826 30823 2860 30857
rect 2219 30765 2253 30799
rect 2325 30765 2359 30799
rect 2219 30693 2253 30727
rect 2325 30693 2359 30727
rect 2219 30621 2253 30655
rect 2325 30621 2359 30655
rect 2219 30549 2253 30583
rect 2325 30549 2359 30583
rect 2219 30477 2253 30511
rect 2325 30477 2359 30511
rect 2219 30405 2253 30439
rect 2325 30405 2359 30439
rect 2219 30333 2253 30367
rect 2325 30333 2359 30367
rect 2219 30261 2253 30295
rect 2325 30261 2359 30295
rect 2219 30189 2253 30223
rect 2325 30189 2359 30223
rect 2219 30117 2253 30151
rect 2325 30117 2359 30151
rect 2219 30045 2253 30079
rect 2325 30045 2359 30079
rect 2219 29973 2253 30007
rect 2325 29973 2359 30007
rect 2219 29901 2253 29935
rect 2325 29901 2359 29935
rect 2219 29829 2253 29863
rect 2325 29829 2359 29863
rect 2219 29757 2253 29791
rect 2325 29757 2359 29791
rect 2219 29685 2253 29719
rect 2325 29685 2359 29719
rect 2219 29613 2253 29647
rect 2325 29613 2359 29647
rect 2219 29541 2253 29575
rect 2325 29541 2359 29575
rect 2219 29469 2253 29503
rect 2325 29469 2359 29503
rect 2219 29397 2253 29431
rect 2325 29397 2359 29431
rect 3173 30680 3207 30714
rect 3245 30680 3279 30714
rect 3173 30607 3207 30641
rect 3245 30607 3279 30641
rect 3173 30534 3207 30568
rect 3245 30534 3279 30568
rect 3173 30461 3207 30495
rect 3245 30461 3279 30495
rect 3173 29380 3279 30422
rect 3591 30680 3625 30714
rect 3663 30680 3697 30714
rect 3591 30607 3625 30641
rect 3663 30607 3697 30641
rect 3591 30534 3625 30568
rect 3663 30534 3697 30568
rect 3591 30461 3625 30495
rect 3663 30461 3697 30495
rect 3591 29380 3697 30422
rect 4009 30680 4043 30714
rect 4081 30680 4115 30714
rect 4009 30607 4043 30641
rect 4081 30607 4115 30641
rect 4009 30534 4043 30568
rect 4081 30534 4115 30568
rect 4009 30461 4043 30495
rect 4081 30461 4115 30495
rect 4009 29380 4115 30422
rect 4427 30680 4461 30714
rect 4499 30680 4533 30714
rect 4427 30607 4461 30641
rect 4499 30607 4533 30641
rect 4427 30534 4461 30568
rect 4499 30534 4533 30568
rect 4427 30461 4461 30495
rect 4499 30461 4533 30495
rect 4427 29380 4533 30422
rect 4845 30680 4879 30714
rect 4917 30680 4951 30714
rect 4845 30607 4879 30641
rect 4917 30607 4951 30641
rect 4845 30534 4879 30568
rect 4917 30534 4951 30568
rect 4845 30461 4879 30495
rect 4917 30461 4951 30495
rect 4845 29380 4951 30422
rect 5263 30680 5297 30714
rect 5335 30680 5369 30714
rect 5263 30607 5297 30641
rect 5335 30607 5369 30641
rect 5263 30534 5297 30568
rect 5335 30534 5369 30568
rect 5263 30461 5297 30495
rect 5335 30461 5369 30495
rect 5263 29380 5369 30422
rect 5681 30680 5715 30714
rect 5753 30680 5787 30714
rect 5681 30607 5715 30641
rect 5753 30607 5787 30641
rect 5681 30534 5715 30568
rect 5753 30534 5787 30568
rect 5681 30461 5715 30495
rect 5753 30461 5787 30495
rect 5681 29380 5787 30422
rect 6099 30680 6133 30714
rect 6171 30680 6205 30714
rect 6099 30607 6133 30641
rect 6171 30607 6205 30641
rect 6099 30534 6133 30568
rect 6171 30534 6205 30568
rect 6099 30461 6133 30495
rect 6171 30461 6205 30495
rect 6099 29380 6205 30422
rect 6517 30680 6551 30714
rect 6589 30680 6623 30714
rect 6517 30607 6551 30641
rect 6589 30607 6623 30641
rect 6517 30534 6551 30568
rect 6589 30534 6623 30568
rect 6517 30461 6551 30495
rect 6589 30461 6623 30495
rect 6517 29380 6623 30422
rect 6935 30680 6969 30714
rect 7007 30680 7041 30714
rect 6935 30607 6969 30641
rect 7007 30607 7041 30641
rect 6935 30534 6969 30568
rect 7007 30534 7041 30568
rect 6935 30461 6969 30495
rect 7007 30461 7041 30495
rect 6935 29380 7041 30422
rect 7353 30680 7387 30714
rect 7425 30680 7459 30714
rect 7353 30607 7387 30641
rect 7425 30607 7459 30641
rect 7353 30534 7387 30568
rect 7425 30534 7459 30568
rect 7353 30461 7387 30495
rect 7425 30461 7459 30495
rect 7353 29380 7459 30422
rect 7771 30680 7805 30714
rect 7843 30680 7877 30714
rect 7771 30607 7805 30641
rect 7843 30607 7877 30641
rect 7771 30534 7805 30568
rect 7843 30534 7877 30568
rect 7771 30461 7805 30495
rect 7843 30461 7877 30495
rect 7771 29380 7877 30422
rect 8189 30680 8223 30714
rect 8261 30680 8295 30714
rect 8189 30607 8223 30641
rect 8261 30607 8295 30641
rect 8189 30534 8223 30568
rect 8261 30534 8295 30568
rect 8189 30461 8223 30495
rect 8261 30461 8295 30495
rect 8189 29380 8295 30422
rect 8607 30680 8641 30714
rect 8679 30680 8713 30714
rect 8607 30607 8641 30641
rect 8679 30607 8713 30641
rect 8607 30534 8641 30568
rect 8679 30534 8713 30568
rect 8607 30461 8641 30495
rect 8679 30461 8713 30495
rect 8607 29380 8713 30422
rect 9025 30680 9059 30714
rect 9097 30680 9131 30714
rect 9025 30607 9059 30641
rect 9097 30607 9131 30641
rect 9025 30534 9059 30568
rect 9097 30534 9131 30568
rect 9025 30461 9059 30495
rect 9097 30461 9131 30495
rect 9025 29380 9131 30422
rect 9443 30680 9477 30714
rect 9515 30680 9549 30714
rect 9443 30607 9477 30641
rect 9515 30607 9549 30641
rect 9443 30534 9477 30568
rect 9515 30534 9549 30568
rect 9443 30461 9477 30495
rect 9515 30461 9549 30495
rect 9443 29380 9549 30422
rect 9861 30680 9895 30714
rect 9933 30680 9967 30714
rect 9861 30607 9895 30641
rect 9933 30607 9967 30641
rect 9861 30534 9895 30568
rect 9933 30534 9967 30568
rect 9861 30461 9895 30495
rect 9933 30461 9967 30495
rect 9861 29380 9967 30422
rect 10279 30680 10313 30714
rect 10351 30680 10385 30714
rect 10279 30607 10313 30641
rect 10351 30607 10385 30641
rect 10279 30534 10313 30568
rect 10351 30534 10385 30568
rect 10279 30461 10313 30495
rect 10351 30461 10385 30495
rect 10279 29380 10385 30422
rect 10697 30680 10731 30714
rect 10769 30680 10803 30714
rect 10697 30607 10731 30641
rect 10769 30607 10803 30641
rect 10697 30534 10731 30568
rect 10769 30534 10803 30568
rect 10697 30461 10731 30495
rect 10769 30461 10803 30495
rect 10697 29380 10803 30422
rect 11115 30680 11149 30714
rect 11187 30680 11221 30714
rect 11115 30607 11149 30641
rect 11187 30607 11221 30641
rect 11115 30534 11149 30568
rect 11187 30534 11221 30568
rect 11115 30461 11149 30495
rect 11187 30461 11221 30495
rect 11115 29380 11221 30422
rect 11533 30680 11567 30714
rect 11605 30680 11639 30714
rect 11533 30607 11567 30641
rect 11605 30607 11639 30641
rect 11533 30534 11567 30568
rect 11605 30534 11639 30568
rect 11533 30461 11567 30495
rect 11605 30461 11639 30495
rect 11533 29380 11639 30422
rect 11951 30680 11985 30714
rect 12023 30680 12057 30714
rect 11951 30607 11985 30641
rect 12023 30607 12057 30641
rect 11951 30534 11985 30568
rect 12023 30534 12057 30568
rect 11951 30461 11985 30495
rect 12023 30461 12057 30495
rect 11951 29380 12057 30422
rect 12369 30680 12403 30714
rect 12441 30680 12475 30714
rect 12369 30607 12403 30641
rect 12441 30607 12475 30641
rect 12369 30534 12403 30568
rect 12441 30534 12475 30568
rect 12369 30461 12403 30495
rect 12441 30461 12475 30495
rect 12369 29380 12475 30422
rect 12787 30680 12821 30714
rect 12859 30680 12893 30714
rect 12787 30607 12821 30641
rect 12859 30607 12893 30641
rect 12787 30534 12821 30568
rect 12859 30534 12893 30568
rect 12787 30461 12821 30495
rect 12859 30461 12893 30495
rect 12787 29380 12893 30422
rect 13205 30680 13239 30714
rect 13277 30680 13311 30714
rect 13205 30607 13239 30641
rect 13277 30607 13311 30641
rect 13205 30534 13239 30568
rect 13277 30534 13311 30568
rect 13205 30461 13239 30495
rect 13277 30461 13311 30495
rect 13205 29380 13311 30422
rect 2219 29325 2253 29359
rect 2325 29325 2359 29359
rect 2219 29253 2253 29287
rect 2325 29253 2359 29287
rect 2219 29181 2253 29215
rect 2325 29181 2359 29215
rect 2219 29109 2253 29143
rect 2325 29109 2359 29143
rect 2674 29286 2708 29320
rect 2750 29286 2784 29320
rect 2826 29286 2860 29320
rect 2674 29205 2708 29239
rect 2750 29205 2784 29239
rect 2826 29205 2860 29239
rect 2674 29123 2708 29157
rect 2750 29123 2784 29157
rect 2826 29123 2860 29157
rect 2219 29037 2253 29071
rect 2325 29037 2359 29071
rect 2219 28965 2253 28999
rect 2325 28995 2359 28999
rect 2325 28965 2342 28995
rect 2342 28965 2359 28995
rect 2219 28893 2253 28927
rect 2325 28893 2342 28927
rect 2342 28893 2359 28927
rect 4845 28680 4879 28714
rect 4917 28680 4951 28714
rect 4845 28607 4879 28641
rect 4917 28607 4951 28641
rect 4845 28534 4879 28568
rect 4917 28534 4951 28568
rect 4845 28461 4879 28495
rect 4917 28461 4951 28495
rect 4845 27380 4951 28422
rect 5263 28680 5297 28714
rect 5335 28680 5369 28714
rect 5263 28607 5297 28641
rect 5335 28607 5369 28641
rect 5263 28534 5297 28568
rect 5335 28534 5369 28568
rect 5263 28461 5297 28495
rect 5335 28461 5369 28495
rect 5263 27380 5369 28422
rect 5681 28680 5715 28714
rect 5753 28680 5787 28714
rect 5681 28607 5715 28641
rect 5753 28607 5787 28641
rect 5681 28534 5715 28568
rect 5753 28534 5787 28568
rect 5681 28461 5715 28495
rect 5753 28461 5787 28495
rect 5681 27380 5787 28422
rect 6099 28680 6133 28714
rect 6171 28680 6205 28714
rect 6099 28607 6133 28641
rect 6171 28607 6205 28641
rect 6099 28534 6133 28568
rect 6171 28534 6205 28568
rect 6099 28461 6133 28495
rect 6171 28461 6205 28495
rect 6099 27380 6205 28422
rect 6517 28680 6551 28714
rect 6589 28680 6623 28714
rect 6517 28607 6551 28641
rect 6589 28607 6623 28641
rect 6517 28534 6551 28568
rect 6589 28534 6623 28568
rect 6517 28461 6551 28495
rect 6589 28461 6623 28495
rect 6517 27380 6623 28422
rect 6935 28680 6969 28714
rect 7007 28680 7041 28714
rect 6935 28607 6969 28641
rect 7007 28607 7041 28641
rect 6935 28534 6969 28568
rect 7007 28534 7041 28568
rect 6935 28461 6969 28495
rect 7007 28461 7041 28495
rect 6935 27380 7041 28422
rect 7353 28680 7387 28714
rect 7425 28680 7459 28714
rect 7353 28607 7387 28641
rect 7425 28607 7459 28641
rect 7353 28534 7387 28568
rect 7425 28534 7459 28568
rect 7353 28461 7387 28495
rect 7425 28461 7459 28495
rect 7353 27380 7459 28422
rect 7771 28680 7805 28714
rect 7843 28680 7877 28714
rect 7771 28607 7805 28641
rect 7843 28607 7877 28641
rect 7771 28534 7805 28568
rect 7843 28534 7877 28568
rect 7771 28461 7805 28495
rect 7843 28461 7877 28495
rect 7771 27380 7877 28422
rect 8189 28680 8223 28714
rect 8261 28680 8295 28714
rect 8189 28607 8223 28641
rect 8261 28607 8295 28641
rect 8189 28534 8223 28568
rect 8261 28534 8295 28568
rect 8189 28461 8223 28495
rect 8261 28461 8295 28495
rect 8189 27380 8295 28422
rect 8607 28680 8641 28714
rect 8679 28680 8713 28714
rect 8607 28607 8641 28641
rect 8679 28607 8713 28641
rect 8607 28534 8641 28568
rect 8679 28534 8713 28568
rect 8607 28461 8641 28495
rect 8679 28461 8713 28495
rect 8607 27380 8713 28422
rect 9025 28680 9059 28714
rect 9097 28680 9131 28714
rect 9025 28607 9059 28641
rect 9097 28607 9131 28641
rect 9025 28534 9059 28568
rect 9097 28534 9131 28568
rect 9025 28461 9059 28495
rect 9097 28461 9131 28495
rect 9025 27380 9131 28422
rect 9443 28680 9477 28714
rect 9515 28680 9549 28714
rect 9443 28607 9477 28641
rect 9515 28607 9549 28641
rect 9443 28534 9477 28568
rect 9515 28534 9549 28568
rect 9443 28461 9477 28495
rect 9515 28461 9549 28495
rect 9443 27380 9549 28422
rect 9861 28680 9895 28714
rect 9933 28680 9967 28714
rect 9861 28607 9895 28641
rect 9933 28607 9967 28641
rect 9861 28534 9895 28568
rect 9933 28534 9967 28568
rect 9861 28461 9895 28495
rect 9933 28461 9967 28495
rect 9861 27380 9967 28422
rect 10279 28680 10313 28714
rect 10351 28680 10385 28714
rect 10279 28607 10313 28641
rect 10351 28607 10385 28641
rect 10279 28534 10313 28568
rect 10351 28534 10385 28568
rect 10279 28461 10313 28495
rect 10351 28461 10385 28495
rect 10279 27380 10385 28422
rect 10697 28680 10731 28714
rect 10769 28680 10803 28714
rect 10697 28607 10731 28641
rect 10769 28607 10803 28641
rect 10697 28534 10731 28568
rect 10769 28534 10803 28568
rect 10697 28461 10731 28495
rect 10769 28461 10803 28495
rect 10697 27380 10803 28422
rect 11115 28680 11149 28714
rect 11187 28680 11221 28714
rect 11115 28607 11149 28641
rect 11187 28607 11221 28641
rect 11115 28534 11149 28568
rect 11187 28534 11221 28568
rect 11115 28461 11149 28495
rect 11187 28461 11221 28495
rect 11115 27380 11221 28422
rect 11533 28680 11567 28714
rect 11605 28680 11639 28714
rect 11533 28607 11567 28641
rect 11605 28607 11639 28641
rect 11533 28534 11567 28568
rect 11605 28534 11639 28568
rect 11533 28461 11567 28495
rect 11605 28461 11639 28495
rect 11533 27380 11639 28422
rect 11951 28680 11985 28714
rect 12023 28680 12057 28714
rect 11951 28607 11985 28641
rect 12023 28607 12057 28641
rect 11951 28534 11985 28568
rect 12023 28534 12057 28568
rect 11951 28461 11985 28495
rect 12023 28461 12057 28495
rect 11951 27380 12057 28422
rect 12369 28680 12403 28714
rect 12441 28680 12475 28714
rect 12369 28607 12403 28641
rect 12441 28607 12475 28641
rect 12369 28534 12403 28568
rect 12441 28534 12475 28568
rect 12369 28461 12403 28495
rect 12441 28461 12475 28495
rect 12369 27380 12475 28422
rect 12787 28680 12821 28714
rect 12859 28680 12893 28714
rect 12787 28607 12821 28641
rect 12859 28607 12893 28641
rect 12787 28534 12821 28568
rect 12859 28534 12893 28568
rect 12787 28461 12821 28495
rect 12859 28461 12893 28495
rect 12787 27380 12893 28422
rect 13205 28680 13239 28714
rect 13277 28680 13311 28714
rect 13205 28607 13239 28641
rect 13277 28607 13311 28641
rect 13205 28534 13239 28568
rect 13277 28534 13311 28568
rect 13205 28461 13239 28495
rect 13277 28461 13311 28495
rect 13205 27380 13311 28422
rect 4339 27287 4373 27321
rect 4415 27287 4449 27321
rect 4491 27287 4525 27321
rect 4339 27210 4373 27244
rect 4415 27210 4449 27244
rect 4491 27210 4525 27244
rect 4339 27133 4373 27167
rect 4415 27133 4449 27167
rect 4491 27133 4525 27167
rect 4339 27055 4373 27089
rect 4415 27055 4449 27089
rect 4491 27055 4525 27089
rect 4339 26977 4373 27011
rect 4415 26977 4449 27011
rect 4491 26977 4525 27011
rect 4339 26899 4373 26933
rect 4415 26899 4449 26933
rect 4491 26899 4525 26933
rect 4339 26821 4373 26855
rect 4415 26821 4449 26855
rect 4491 26821 4525 26855
rect 4845 26718 4879 26752
rect 4917 26718 4951 26752
rect 4845 26643 4879 26677
rect 4917 26643 4951 26677
rect 4845 26568 4879 26602
rect 4917 26568 4951 26602
rect 4845 26493 4879 26527
rect 4917 26493 4951 26527
rect 4845 26418 4879 26452
rect 4917 26418 4951 26452
rect 4845 26343 4879 26377
rect 4917 26343 4951 26377
rect 4845 26268 4879 26302
rect 4917 26268 4951 26302
rect 4845 26193 4879 26227
rect 4917 26193 4951 26227
rect 4845 26118 4879 26152
rect 4917 26118 4951 26152
rect 4845 26043 4879 26077
rect 4917 26043 4951 26077
rect 4845 25968 4879 26002
rect 4917 25968 4951 26002
rect 4845 25894 4879 25928
rect 4917 25894 4951 25928
rect 4845 25820 4879 25854
rect 4917 25820 4951 25854
rect 4845 25746 4879 25780
rect 4917 25746 4951 25780
rect 5263 26709 5297 26743
rect 5335 26709 5369 26743
rect 5263 26634 5297 26668
rect 5335 26634 5369 26668
rect 5263 26560 5297 26594
rect 5335 26560 5369 26594
rect 5263 26486 5297 26520
rect 5335 26486 5369 26520
rect 5263 26412 5297 26446
rect 5335 26412 5369 26446
rect 5263 26338 5297 26372
rect 5335 26338 5369 26372
rect 5263 26264 5297 26298
rect 5335 26264 5369 26298
rect 5263 26190 5297 26224
rect 5335 26190 5369 26224
rect 5263 26116 5297 26150
rect 5335 26116 5369 26150
rect 5263 26042 5297 26076
rect 5335 26042 5369 26076
rect 5263 25968 5297 26002
rect 5335 25968 5369 26002
rect 5263 25894 5297 25928
rect 5335 25894 5369 25928
rect 5263 25820 5297 25854
rect 5335 25820 5369 25854
rect 5263 25746 5297 25780
rect 5335 25746 5369 25780
rect 5681 26718 5715 26752
rect 5753 26718 5787 26752
rect 5681 26645 5715 26679
rect 5753 26645 5787 26679
rect 5681 26572 5715 26606
rect 5753 26572 5787 26606
rect 5681 26499 5715 26533
rect 5753 26499 5787 26533
rect 5681 26426 5715 26460
rect 5753 26426 5787 26460
rect 5681 26353 5715 26387
rect 5753 26353 5787 26387
rect 5681 26280 5715 26314
rect 5753 26280 5787 26314
rect 5681 26207 5715 26241
rect 5753 26207 5787 26241
rect 5681 26134 5715 26168
rect 5753 26134 5787 26168
rect 5681 26061 5715 26095
rect 5753 26061 5787 26095
rect 5681 25772 5787 26022
rect 6099 26709 6133 26743
rect 6171 26709 6205 26743
rect 6099 26634 6133 26668
rect 6171 26634 6205 26668
rect 6099 26560 6133 26594
rect 6171 26560 6205 26594
rect 6099 26486 6133 26520
rect 6171 26486 6205 26520
rect 6099 26412 6133 26446
rect 6171 26412 6205 26446
rect 6099 26338 6133 26372
rect 6171 26338 6205 26372
rect 6099 26264 6133 26298
rect 6171 26264 6205 26298
rect 6099 26190 6133 26224
rect 6171 26190 6205 26224
rect 6099 26116 6133 26150
rect 6171 26116 6205 26150
rect 6099 26042 6133 26076
rect 6171 26042 6205 26076
rect 6099 25968 6133 26002
rect 6171 25968 6205 26002
rect 6099 25894 6133 25928
rect 6171 25894 6205 25928
rect 6099 25820 6133 25854
rect 6171 25820 6205 25854
rect 6099 25746 6133 25780
rect 6171 25746 6205 25780
rect 6517 26717 6551 26751
rect 6589 26717 6623 26751
rect 6517 26642 6551 26676
rect 6589 26642 6623 26676
rect 6517 26567 6551 26601
rect 6589 26567 6623 26601
rect 6517 26492 6551 26526
rect 6589 26492 6623 26526
rect 6517 26417 6551 26451
rect 6589 26417 6623 26451
rect 6517 26342 6551 26376
rect 6589 26342 6623 26376
rect 6517 26267 6551 26301
rect 6589 26267 6623 26301
rect 6517 26192 6551 26226
rect 6589 26192 6623 26226
rect 6517 26117 6551 26151
rect 6589 26117 6623 26151
rect 6517 26042 6551 26076
rect 6589 26042 6623 26076
rect 6517 25968 6551 26002
rect 6589 25968 6623 26002
rect 6517 25894 6551 25928
rect 6589 25894 6623 25928
rect 6517 25820 6551 25854
rect 6589 25820 6623 25854
rect 6517 25746 6551 25780
rect 6589 25746 6623 25780
rect 6935 26734 6969 26768
rect 7007 26734 7041 26768
rect 7771 26751 7805 26785
rect 7843 26751 7877 26785
rect 8607 26751 8641 26785
rect 8679 26751 8713 26785
rect 9443 26751 9477 26785
rect 9515 26751 9549 26785
rect 10279 26751 10313 26785
rect 10351 26751 10385 26785
rect 11115 26751 11149 26785
rect 11187 26751 11221 26785
rect 11951 26751 11985 26785
rect 12023 26751 12057 26785
rect 12787 26751 12821 26785
rect 12859 26751 12893 26785
rect 6935 26658 6969 26692
rect 7007 26658 7041 26692
rect 6935 26582 6969 26616
rect 7007 26582 7041 26616
rect 6935 26506 6969 26540
rect 7007 26506 7041 26540
rect 6935 26430 6969 26464
rect 7007 26430 7041 26464
rect 6935 26354 6969 26388
rect 7007 26354 7041 26388
rect 6935 26278 6969 26312
rect 7007 26278 7041 26312
rect 6935 26202 6969 26236
rect 7007 26202 7041 26236
rect 6935 26126 6969 26160
rect 7007 26126 7041 26160
rect 6935 26050 6969 26084
rect 7007 26050 7041 26084
rect 6935 25974 6969 26008
rect 7007 25974 7041 26008
rect 6935 25898 6969 25932
rect 7007 25898 7041 25932
rect 6935 25822 6969 25856
rect 7007 25822 7041 25856
rect 6935 25746 6969 25780
rect 7007 25746 7041 25780
rect 7353 26717 7387 26751
rect 7425 26717 7459 26751
rect 7353 26642 7387 26676
rect 7425 26642 7459 26676
rect 7353 26567 7387 26601
rect 7425 26567 7459 26601
rect 7353 26492 7387 26526
rect 7425 26492 7459 26526
rect 7353 26417 7387 26451
rect 7425 26417 7459 26451
rect 7353 26342 7387 26376
rect 7425 26342 7459 26376
rect 7353 26267 7387 26301
rect 7425 26267 7459 26301
rect 7353 26192 7387 26226
rect 7425 26192 7459 26226
rect 7353 26117 7387 26151
rect 7425 26117 7459 26151
rect 7353 26042 7387 26076
rect 7425 26042 7459 26076
rect 7353 25968 7387 26002
rect 7425 25968 7459 26002
rect 7353 25894 7387 25928
rect 7425 25894 7459 25928
rect 7353 25820 7387 25854
rect 7425 25820 7459 25854
rect 7353 25746 7387 25780
rect 7425 25746 7459 25780
rect 7771 26673 7805 26707
rect 7843 26673 7877 26707
rect 7771 26595 7805 26629
rect 7843 26595 7877 26629
rect 7771 26517 7805 26551
rect 7843 26517 7877 26551
rect 7771 26439 7805 26473
rect 7843 26439 7877 26473
rect 7771 26362 7805 26396
rect 7843 26362 7877 26396
rect 7771 26285 7805 26319
rect 7843 26285 7877 26319
rect 7771 26208 7805 26242
rect 7843 26208 7877 26242
rect 7771 26131 7805 26165
rect 7843 26131 7877 26165
rect 7771 26054 7805 26088
rect 7843 26054 7877 26088
rect 7771 25977 7805 26011
rect 7843 25977 7877 26011
rect 7771 25900 7805 25934
rect 7843 25900 7877 25934
rect 7771 25823 7805 25857
rect 7843 25823 7877 25857
rect 7771 25746 7805 25780
rect 7843 25746 7877 25780
rect 8189 26717 8223 26751
rect 8261 26717 8295 26751
rect 8189 26642 8223 26676
rect 8261 26642 8295 26676
rect 8189 26567 8223 26601
rect 8261 26567 8295 26601
rect 8189 26492 8223 26526
rect 8261 26492 8295 26526
rect 8189 26417 8223 26451
rect 8261 26417 8295 26451
rect 8189 26342 8223 26376
rect 8261 26342 8295 26376
rect 8189 26267 8223 26301
rect 8261 26267 8295 26301
rect 8189 26192 8223 26226
rect 8261 26192 8295 26226
rect 8189 26117 8223 26151
rect 8261 26117 8295 26151
rect 8189 26042 8223 26076
rect 8261 26042 8295 26076
rect 8189 25968 8223 26002
rect 8261 25968 8295 26002
rect 8189 25894 8223 25928
rect 8261 25894 8295 25928
rect 8189 25820 8223 25854
rect 8261 25820 8295 25854
rect 8189 25746 8223 25780
rect 8261 25746 8295 25780
rect 8607 26673 8641 26707
rect 8679 26673 8713 26707
rect 8607 26595 8641 26629
rect 8679 26595 8713 26629
rect 8607 26517 8641 26551
rect 8679 26517 8713 26551
rect 8607 26439 8641 26473
rect 8679 26439 8713 26473
rect 8607 26362 8641 26396
rect 8679 26362 8713 26396
rect 8607 26285 8641 26319
rect 8679 26285 8713 26319
rect 8607 26208 8641 26242
rect 8679 26208 8713 26242
rect 8607 26131 8641 26165
rect 8679 26131 8713 26165
rect 8607 26054 8641 26088
rect 8679 26054 8713 26088
rect 8607 25977 8641 26011
rect 8679 25977 8713 26011
rect 8607 25900 8641 25934
rect 8679 25900 8713 25934
rect 8607 25823 8641 25857
rect 8679 25823 8713 25857
rect 8607 25746 8641 25780
rect 8679 25746 8713 25780
rect 9025 26717 9059 26751
rect 9097 26717 9131 26751
rect 9025 26642 9059 26676
rect 9097 26642 9131 26676
rect 9025 26567 9059 26601
rect 9097 26567 9131 26601
rect 9025 26492 9059 26526
rect 9097 26492 9131 26526
rect 9025 26417 9059 26451
rect 9097 26417 9131 26451
rect 9025 26342 9059 26376
rect 9097 26342 9131 26376
rect 9025 26267 9059 26301
rect 9097 26267 9131 26301
rect 9025 26192 9059 26226
rect 9097 26192 9131 26226
rect 9025 26117 9059 26151
rect 9097 26117 9131 26151
rect 9025 26042 9059 26076
rect 9097 26042 9131 26076
rect 9025 25968 9059 26002
rect 9097 25968 9131 26002
rect 9025 25894 9059 25928
rect 9097 25894 9131 25928
rect 9025 25820 9059 25854
rect 9097 25820 9131 25854
rect 9025 25746 9059 25780
rect 9097 25746 9131 25780
rect 9443 26673 9477 26707
rect 9515 26673 9549 26707
rect 9443 26595 9477 26629
rect 9515 26595 9549 26629
rect 9443 26517 9477 26551
rect 9515 26517 9549 26551
rect 9443 26439 9477 26473
rect 9515 26439 9549 26473
rect 9443 26362 9477 26396
rect 9515 26362 9549 26396
rect 9443 26285 9477 26319
rect 9515 26285 9549 26319
rect 9443 26208 9477 26242
rect 9515 26208 9549 26242
rect 9443 26131 9477 26165
rect 9515 26131 9549 26165
rect 9443 26054 9477 26088
rect 9515 26054 9549 26088
rect 9443 25977 9477 26011
rect 9515 25977 9549 26011
rect 9443 25900 9477 25934
rect 9515 25900 9549 25934
rect 9443 25823 9477 25857
rect 9515 25823 9549 25857
rect 9443 25746 9477 25780
rect 9515 25746 9549 25780
rect 9861 26717 9895 26751
rect 9933 26717 9967 26751
rect 9861 26642 9895 26676
rect 9933 26642 9967 26676
rect 9861 26567 9895 26601
rect 9933 26567 9967 26601
rect 9861 26492 9895 26526
rect 9933 26492 9967 26526
rect 9861 26417 9895 26451
rect 9933 26417 9967 26451
rect 9861 26342 9895 26376
rect 9933 26342 9967 26376
rect 9861 26267 9895 26301
rect 9933 26267 9967 26301
rect 9861 26192 9895 26226
rect 9933 26192 9967 26226
rect 9861 26117 9895 26151
rect 9933 26117 9967 26151
rect 9861 26042 9895 26076
rect 9933 26042 9967 26076
rect 9861 25968 9895 26002
rect 9933 25968 9967 26002
rect 9861 25894 9895 25928
rect 9933 25894 9967 25928
rect 9861 25820 9895 25854
rect 9933 25820 9967 25854
rect 9861 25746 9895 25780
rect 9933 25746 9967 25780
rect 10279 26673 10313 26707
rect 10351 26673 10385 26707
rect 10279 26595 10313 26629
rect 10351 26595 10385 26629
rect 10279 26517 10313 26551
rect 10351 26517 10385 26551
rect 10279 26439 10313 26473
rect 10351 26439 10385 26473
rect 10279 26362 10313 26396
rect 10351 26362 10385 26396
rect 10279 26285 10313 26319
rect 10351 26285 10385 26319
rect 10279 26208 10313 26242
rect 10351 26208 10385 26242
rect 10279 26131 10313 26165
rect 10351 26131 10385 26165
rect 10279 26054 10313 26088
rect 10351 26054 10385 26088
rect 10279 25977 10313 26011
rect 10351 25977 10385 26011
rect 10279 25900 10313 25934
rect 10351 25900 10385 25934
rect 10279 25823 10313 25857
rect 10351 25823 10385 25857
rect 10279 25746 10313 25780
rect 10351 25746 10385 25780
rect 10697 26717 10731 26751
rect 10769 26717 10803 26751
rect 10697 26642 10731 26676
rect 10769 26642 10803 26676
rect 10697 26567 10731 26601
rect 10769 26567 10803 26601
rect 10697 26492 10731 26526
rect 10769 26492 10803 26526
rect 10697 26417 10731 26451
rect 10769 26417 10803 26451
rect 10697 26342 10731 26376
rect 10769 26342 10803 26376
rect 10697 26267 10731 26301
rect 10769 26267 10803 26301
rect 10697 26192 10731 26226
rect 10769 26192 10803 26226
rect 10697 26117 10731 26151
rect 10769 26117 10803 26151
rect 10697 26042 10731 26076
rect 10769 26042 10803 26076
rect 10697 25968 10731 26002
rect 10769 25968 10803 26002
rect 10697 25894 10731 25928
rect 10769 25894 10803 25928
rect 10697 25820 10731 25854
rect 10769 25820 10803 25854
rect 10697 25746 10731 25780
rect 10769 25746 10803 25780
rect 11115 26673 11149 26707
rect 11187 26673 11221 26707
rect 11115 26595 11149 26629
rect 11187 26595 11221 26629
rect 11115 26517 11149 26551
rect 11187 26517 11221 26551
rect 11115 26439 11149 26473
rect 11187 26439 11221 26473
rect 11115 26362 11149 26396
rect 11187 26362 11221 26396
rect 11115 26285 11149 26319
rect 11187 26285 11221 26319
rect 11115 26208 11149 26242
rect 11187 26208 11221 26242
rect 11115 26131 11149 26165
rect 11187 26131 11221 26165
rect 11115 26054 11149 26088
rect 11187 26054 11221 26088
rect 11115 25977 11149 26011
rect 11187 25977 11221 26011
rect 11115 25900 11149 25934
rect 11187 25900 11221 25934
rect 11115 25823 11149 25857
rect 11187 25823 11221 25857
rect 11115 25746 11149 25780
rect 11187 25746 11221 25780
rect 11533 26717 11567 26751
rect 11605 26717 11639 26751
rect 11533 26642 11567 26676
rect 11605 26642 11639 26676
rect 11533 26567 11567 26601
rect 11605 26567 11639 26601
rect 11533 26492 11567 26526
rect 11605 26492 11639 26526
rect 11533 26417 11567 26451
rect 11605 26417 11639 26451
rect 11533 26342 11567 26376
rect 11605 26342 11639 26376
rect 11533 26267 11567 26301
rect 11605 26267 11639 26301
rect 11533 26192 11567 26226
rect 11605 26192 11639 26226
rect 11533 26117 11567 26151
rect 11605 26117 11639 26151
rect 11533 26042 11567 26076
rect 11605 26042 11639 26076
rect 11533 25968 11567 26002
rect 11605 25968 11639 26002
rect 11533 25894 11567 25928
rect 11605 25894 11639 25928
rect 11533 25820 11567 25854
rect 11605 25820 11639 25854
rect 11533 25746 11567 25780
rect 11605 25746 11639 25780
rect 11951 26673 11985 26707
rect 12023 26673 12057 26707
rect 11951 26595 11985 26629
rect 12023 26595 12057 26629
rect 11951 26517 11985 26551
rect 12023 26517 12057 26551
rect 11951 26439 11985 26473
rect 12023 26439 12057 26473
rect 11951 26362 11985 26396
rect 12023 26362 12057 26396
rect 11951 26285 11985 26319
rect 12023 26285 12057 26319
rect 11951 26208 11985 26242
rect 12023 26208 12057 26242
rect 11951 26131 11985 26165
rect 12023 26131 12057 26165
rect 11951 26054 11985 26088
rect 12023 26054 12057 26088
rect 11951 25977 11985 26011
rect 12023 25977 12057 26011
rect 11951 25900 11985 25934
rect 12023 25900 12057 25934
rect 11951 25823 11985 25857
rect 12023 25823 12057 25857
rect 11951 25746 11985 25780
rect 12023 25746 12057 25780
rect 12369 26717 12403 26751
rect 12441 26717 12475 26751
rect 12369 26642 12403 26676
rect 12441 26642 12475 26676
rect 12369 26567 12403 26601
rect 12441 26567 12475 26601
rect 12369 26492 12403 26526
rect 12441 26492 12475 26526
rect 12369 26417 12403 26451
rect 12441 26417 12475 26451
rect 12369 26342 12403 26376
rect 12441 26342 12475 26376
rect 12369 26267 12403 26301
rect 12441 26267 12475 26301
rect 12369 26192 12403 26226
rect 12441 26192 12475 26226
rect 12369 26117 12403 26151
rect 12441 26117 12475 26151
rect 12369 26042 12403 26076
rect 12441 26042 12475 26076
rect 12369 25968 12403 26002
rect 12441 25968 12475 26002
rect 12369 25894 12403 25928
rect 12441 25894 12475 25928
rect 12369 25820 12403 25854
rect 12441 25820 12475 25854
rect 12369 25746 12403 25780
rect 12441 25746 12475 25780
rect 12787 26673 12821 26707
rect 12859 26673 12893 26707
rect 12787 26595 12821 26629
rect 12859 26595 12893 26629
rect 12787 26517 12821 26551
rect 12859 26517 12893 26551
rect 12787 26439 12821 26473
rect 12859 26439 12893 26473
rect 12787 26362 12821 26396
rect 12859 26362 12893 26396
rect 12787 26285 12821 26319
rect 12859 26285 12893 26319
rect 12787 26208 12821 26242
rect 12859 26208 12893 26242
rect 12787 26131 12821 26165
rect 12859 26131 12893 26165
rect 12787 26054 12821 26088
rect 12859 26054 12893 26088
rect 12787 25977 12821 26011
rect 12859 25977 12893 26011
rect 12787 25900 12821 25934
rect 12859 25900 12893 25934
rect 12787 25823 12821 25857
rect 12859 25823 12893 25857
rect 12787 25746 12821 25780
rect 12859 25746 12893 25780
rect 13205 26717 13239 26751
rect 13277 26717 13311 26751
rect 13205 26642 13239 26676
rect 13277 26642 13311 26676
rect 13205 26567 13239 26601
rect 13277 26567 13311 26601
rect 13205 26492 13239 26526
rect 13277 26492 13311 26526
rect 13205 26417 13239 26451
rect 13277 26417 13311 26451
rect 13205 26342 13239 26376
rect 13277 26342 13311 26376
rect 13205 26267 13239 26301
rect 13277 26267 13311 26301
rect 13205 26192 13239 26226
rect 13277 26192 13311 26226
rect 13205 26117 13239 26151
rect 13277 26117 13311 26151
rect 13205 26042 13239 26076
rect 13277 26042 13311 26076
rect 13205 25968 13239 26002
rect 13277 25968 13311 26002
rect 13205 25894 13239 25928
rect 13277 25894 13311 25928
rect 13205 25820 13239 25854
rect 13277 25820 13311 25854
rect 13205 25746 13239 25780
rect 13277 25746 13311 25780
rect 4344 25636 4378 25670
rect 4486 25636 4520 25670
rect 4727 25025 4761 25059
rect 4727 24952 4761 24986
rect 4727 24880 4761 24914
rect 4727 24808 4761 24842
rect 4727 24736 4761 24770
rect 4727 24664 4761 24698
rect 4727 24592 4761 24626
rect 4727 24520 4761 24554
rect 4727 24448 4761 24482
rect 4727 24376 4761 24410
rect 4727 24304 4761 24338
rect 4727 24232 4761 24266
rect 4727 24160 4761 24194
rect 4727 24088 4761 24122
rect 4727 24016 4761 24050
rect 5073 24938 5107 24972
rect 5073 24861 5107 24895
rect 5073 24784 5107 24818
rect 5073 24707 5107 24741
rect 5073 24630 5107 24664
rect 5073 24553 5107 24587
rect 5073 24476 5107 24510
rect 5073 24399 5107 24433
rect 5073 24322 5107 24356
rect 5073 24245 5107 24279
rect 5073 24168 5107 24202
rect 5073 24092 5107 24126
rect 5073 24016 5107 24050
rect 6719 24938 6753 24972
rect 6719 24861 6753 24895
rect 6719 24784 6753 24818
rect 6719 24707 6753 24741
rect 6719 24630 6753 24664
rect 6719 24553 6753 24587
rect 6719 24476 6753 24510
rect 6719 24399 6753 24433
rect 6719 24322 6753 24356
rect 6719 24245 6753 24279
rect 6719 24168 6753 24202
rect 6719 24092 6753 24126
rect 6719 24016 6753 24050
rect 8374 24938 8408 24972
rect 8374 24861 8408 24895
rect 8374 24784 8408 24818
rect 8374 24707 8408 24741
rect 8374 24630 8408 24664
rect 8374 24553 8408 24587
rect 8374 24476 8408 24510
rect 8374 24399 8408 24433
rect 8374 24322 8408 24356
rect 8374 24245 8408 24279
rect 8374 24168 8408 24202
rect 8374 24092 8408 24126
rect 8374 24016 8408 24050
rect 10030 24938 10064 24972
rect 10030 24861 10064 24895
rect 10030 24784 10064 24818
rect 10030 24707 10064 24741
rect 10030 24630 10064 24664
rect 10030 24553 10064 24587
rect 10030 24476 10064 24510
rect 10030 24399 10064 24433
rect 10030 24322 10064 24356
rect 10030 24245 10064 24279
rect 10030 24168 10064 24202
rect 10030 24092 10064 24126
rect 10030 24016 10064 24050
rect 11686 24938 11720 24972
rect 11686 24861 11720 24895
rect 11686 24784 11720 24818
rect 11686 24707 11720 24741
rect 11686 24630 11720 24664
rect 11686 24553 11720 24587
rect 11686 24476 11720 24510
rect 11686 24399 11720 24433
rect 11686 24322 11720 24356
rect 11686 24245 11720 24279
rect 11686 24168 11720 24202
rect 11686 24092 11720 24126
rect 11686 24016 11720 24050
rect 13342 24938 13376 24972
rect 13342 24861 13376 24895
rect 13342 24784 13376 24818
rect 13342 24707 13376 24741
rect 13342 24630 13376 24664
rect 13342 24553 13376 24587
rect 13342 24476 13376 24510
rect 13342 24399 13376 24433
rect 13342 24322 13376 24356
rect 13342 24245 13376 24279
rect 13342 24168 13376 24202
rect 13342 24092 13376 24126
rect 13342 24016 13376 24050
rect 5081 23663 5090 23697
rect 5090 23663 5115 23697
rect 5154 23663 5158 23697
rect 5158 23663 5188 23697
rect 5227 23663 5260 23697
rect 5260 23663 5261 23697
rect 5300 23663 5328 23697
rect 5328 23663 5334 23697
rect 5373 23663 5396 23697
rect 5396 23663 5407 23697
rect 5446 23663 5464 23697
rect 5464 23663 5480 23697
rect 5519 23663 5532 23697
rect 5532 23663 5553 23697
rect 5592 23663 5600 23697
rect 5600 23663 5626 23697
rect 5665 23663 5668 23697
rect 5668 23663 5699 23697
rect 5737 23663 5770 23697
rect 5770 23663 5771 23697
rect 5809 23663 5838 23697
rect 5838 23663 5843 23697
rect 5881 23663 5906 23697
rect 5906 23663 5915 23697
rect 5953 23663 5974 23697
rect 5974 23663 5987 23697
rect 6025 23663 6042 23697
rect 6042 23663 6059 23697
rect 6097 23663 6110 23697
rect 6110 23663 6131 23697
rect 6169 23663 6178 23697
rect 6178 23663 6203 23697
rect 6241 23663 6246 23697
rect 6246 23663 6275 23697
rect 6313 23663 6314 23697
rect 6314 23663 6347 23697
rect 6385 23663 6416 23697
rect 6416 23663 6419 23697
rect 6457 23663 6484 23697
rect 6484 23663 6491 23697
rect 6529 23663 6552 23697
rect 6552 23663 6563 23697
rect 6601 23663 6620 23697
rect 6620 23663 6635 23697
rect 6673 23663 6688 23697
rect 6688 23663 6707 23697
rect 6745 23663 6756 23697
rect 6756 23663 6779 23697
rect 6817 23663 6824 23697
rect 6824 23663 6851 23697
rect 6889 23663 6892 23697
rect 6892 23663 6923 23697
rect 6961 23663 6994 23697
rect 6994 23663 6995 23697
rect 7033 23663 7062 23697
rect 7062 23663 7067 23697
rect 7105 23663 7130 23697
rect 7130 23663 7139 23697
rect 7177 23663 7198 23697
rect 7198 23663 7211 23697
rect 7249 23663 7266 23697
rect 7266 23663 7283 23697
rect 7321 23663 7334 23697
rect 7334 23663 7355 23697
rect 7393 23663 7402 23697
rect 7402 23663 7427 23697
rect 7465 23663 7470 23697
rect 7470 23663 7499 23697
rect 7537 23663 7538 23697
rect 7538 23663 7571 23697
rect 7609 23663 7640 23697
rect 7640 23663 7643 23697
rect 7681 23663 7708 23697
rect 7708 23663 7715 23697
rect 7753 23663 7776 23697
rect 7776 23663 7787 23697
rect 7825 23663 7844 23697
rect 7844 23663 7859 23697
rect 7897 23663 7912 23697
rect 7912 23663 7931 23697
rect 7969 23663 7980 23697
rect 7980 23663 8003 23697
rect 8041 23663 8048 23697
rect 8048 23663 8075 23697
rect 8113 23663 8116 23697
rect 8116 23663 8147 23697
rect 8185 23663 8218 23697
rect 8218 23663 8219 23697
rect 8257 23663 8286 23697
rect 8286 23663 8291 23697
rect 8329 23663 8354 23697
rect 8354 23663 8363 23697
rect 8401 23663 8422 23697
rect 8422 23663 8435 23697
rect 8473 23663 8490 23697
rect 8490 23663 8507 23697
rect 8545 23663 8558 23697
rect 8558 23663 8579 23697
rect 8617 23663 8626 23697
rect 8626 23663 8651 23697
rect 8689 23663 8694 23697
rect 8694 23663 8723 23697
rect 8761 23663 8762 23697
rect 8762 23663 8795 23697
rect 8833 23663 8864 23697
rect 8864 23663 8867 23697
rect 8905 23663 8932 23697
rect 8932 23663 8939 23697
rect 8977 23663 9000 23697
rect 9000 23663 9011 23697
rect 9049 23663 9068 23697
rect 9068 23663 9083 23697
rect 9121 23663 9136 23697
rect 9136 23663 9155 23697
rect 9193 23663 9204 23697
rect 9204 23663 9227 23697
rect 9265 23663 9272 23697
rect 9272 23663 9299 23697
rect 9337 23663 9340 23697
rect 9340 23663 9371 23697
rect 9409 23663 9442 23697
rect 9442 23663 9443 23697
rect 9481 23663 9510 23697
rect 9510 23663 9515 23697
rect 9553 23663 9578 23697
rect 9578 23663 9587 23697
rect 9625 23663 9646 23697
rect 9646 23663 9659 23697
rect 9697 23663 9714 23697
rect 9714 23663 9731 23697
rect 9769 23663 9782 23697
rect 9782 23663 9803 23697
rect 9841 23663 9850 23697
rect 9850 23663 9875 23697
rect 9913 23663 9918 23697
rect 9918 23663 9947 23697
rect 9985 23663 9986 23697
rect 9986 23663 10019 23697
rect 10057 23663 10088 23697
rect 10088 23663 10091 23697
rect 10129 23663 10156 23697
rect 10156 23663 10163 23697
rect 10201 23663 10224 23697
rect 10224 23663 10235 23697
rect 10273 23663 10292 23697
rect 10292 23663 10307 23697
rect 10345 23663 10360 23697
rect 10360 23663 10379 23697
rect 10417 23663 10428 23697
rect 10428 23663 10451 23697
rect 10489 23663 10496 23697
rect 10496 23663 10523 23697
rect 10561 23663 10564 23697
rect 10564 23663 10595 23697
rect 10633 23663 10666 23697
rect 10666 23663 10667 23697
rect 10705 23663 10734 23697
rect 10734 23663 10739 23697
rect 10777 23663 10802 23697
rect 10802 23663 10811 23697
rect 10849 23663 10870 23697
rect 10870 23663 10883 23697
rect 10921 23663 10938 23697
rect 10938 23663 10955 23697
rect 10993 23663 11006 23697
rect 11006 23663 11027 23697
rect 11065 23663 11074 23697
rect 11074 23663 11099 23697
rect 11137 23663 11142 23697
rect 11142 23663 11171 23697
rect 11209 23663 11210 23697
rect 11210 23663 11243 23697
rect 11281 23663 11312 23697
rect 11312 23663 11315 23697
rect 11353 23663 11380 23697
rect 11380 23663 11387 23697
rect 11425 23663 11448 23697
rect 11448 23663 11459 23697
rect 11497 23663 11516 23697
rect 11516 23663 11531 23697
rect 11569 23663 11584 23697
rect 11584 23663 11603 23697
rect 11641 23663 11652 23697
rect 11652 23663 11675 23697
rect 11713 23663 11720 23697
rect 11720 23663 11747 23697
rect 11785 23663 11788 23697
rect 11788 23663 11819 23697
rect 11857 23663 11890 23697
rect 11890 23663 11891 23697
rect 11929 23663 11958 23697
rect 11958 23663 11963 23697
rect 12001 23663 12026 23697
rect 12026 23663 12035 23697
rect 12073 23663 12094 23697
rect 12094 23663 12107 23697
rect 12145 23663 12162 23697
rect 12162 23663 12179 23697
rect 12217 23663 12230 23697
rect 12230 23663 12251 23697
rect 12289 23663 12298 23697
rect 12298 23663 12323 23697
rect 12361 23663 12366 23697
rect 12366 23663 12395 23697
rect 12433 23663 12434 23697
rect 12434 23663 12467 23697
rect 12505 23663 12536 23697
rect 12536 23663 12539 23697
rect 12577 23663 12604 23697
rect 12604 23663 12611 23697
rect 12649 23663 12672 23697
rect 12672 23663 12683 23697
rect 12721 23663 12740 23697
rect 12740 23663 12755 23697
rect 12793 23663 12808 23697
rect 12808 23663 12827 23697
rect 12865 23663 12876 23697
rect 12876 23663 12899 23697
rect 12937 23663 12944 23697
rect 12944 23663 12971 23697
rect 13009 23663 13012 23697
rect 13012 23663 13043 23697
rect 13081 23663 13114 23697
rect 13114 23663 13115 23697
rect 13153 23663 13182 23697
rect 13182 23663 13187 23697
rect 13225 23663 13250 23697
rect 13250 23663 13259 23697
rect 13297 23663 13331 23697
rect 5081 23428 5090 23462
rect 5090 23428 5115 23462
rect 5154 23428 5158 23462
rect 5158 23428 5188 23462
rect 5227 23428 5260 23462
rect 5260 23428 5261 23462
rect 5300 23428 5328 23462
rect 5328 23428 5334 23462
rect 5373 23428 5396 23462
rect 5396 23428 5407 23462
rect 5446 23428 5464 23462
rect 5464 23428 5480 23462
rect 5519 23428 5532 23462
rect 5532 23428 5553 23462
rect 5592 23428 5600 23462
rect 5600 23428 5626 23462
rect 5665 23428 5668 23462
rect 5668 23428 5699 23462
rect 5737 23428 5770 23462
rect 5770 23428 5771 23462
rect 5809 23428 5838 23462
rect 5838 23428 5843 23462
rect 5881 23428 5906 23462
rect 5906 23428 5915 23462
rect 5953 23428 5974 23462
rect 5974 23428 5987 23462
rect 6025 23428 6042 23462
rect 6042 23428 6059 23462
rect 6097 23428 6110 23462
rect 6110 23428 6131 23462
rect 6169 23428 6178 23462
rect 6178 23428 6203 23462
rect 6241 23428 6246 23462
rect 6246 23428 6275 23462
rect 6313 23428 6314 23462
rect 6314 23428 6347 23462
rect 6385 23428 6416 23462
rect 6416 23428 6419 23462
rect 6457 23428 6484 23462
rect 6484 23428 6491 23462
rect 6529 23428 6552 23462
rect 6552 23428 6563 23462
rect 6601 23428 6620 23462
rect 6620 23428 6635 23462
rect 6673 23428 6688 23462
rect 6688 23428 6707 23462
rect 6745 23428 6756 23462
rect 6756 23428 6779 23462
rect 6817 23428 6824 23462
rect 6824 23428 6851 23462
rect 6889 23428 6892 23462
rect 6892 23428 6923 23462
rect 6961 23428 6994 23462
rect 6994 23428 6995 23462
rect 7033 23428 7062 23462
rect 7062 23428 7067 23462
rect 7105 23428 7130 23462
rect 7130 23428 7139 23462
rect 7177 23428 7198 23462
rect 7198 23428 7211 23462
rect 7249 23428 7266 23462
rect 7266 23428 7283 23462
rect 7321 23428 7334 23462
rect 7334 23428 7355 23462
rect 7393 23428 7402 23462
rect 7402 23428 7427 23462
rect 7465 23428 7470 23462
rect 7470 23428 7499 23462
rect 7537 23428 7538 23462
rect 7538 23428 7571 23462
rect 7609 23428 7640 23462
rect 7640 23428 7643 23462
rect 7681 23428 7708 23462
rect 7708 23428 7715 23462
rect 7753 23428 7776 23462
rect 7776 23428 7787 23462
rect 7825 23428 7844 23462
rect 7844 23428 7859 23462
rect 7897 23428 7912 23462
rect 7912 23428 7931 23462
rect 7969 23428 7980 23462
rect 7980 23428 8003 23462
rect 8041 23428 8048 23462
rect 8048 23428 8075 23462
rect 8113 23428 8116 23462
rect 8116 23428 8147 23462
rect 8185 23428 8218 23462
rect 8218 23428 8219 23462
rect 8257 23428 8286 23462
rect 8286 23428 8291 23462
rect 8329 23428 8354 23462
rect 8354 23428 8363 23462
rect 8401 23428 8422 23462
rect 8422 23428 8435 23462
rect 8473 23428 8490 23462
rect 8490 23428 8507 23462
rect 8545 23428 8558 23462
rect 8558 23428 8579 23462
rect 8617 23428 8626 23462
rect 8626 23428 8651 23462
rect 8689 23428 8694 23462
rect 8694 23428 8723 23462
rect 8761 23428 8762 23462
rect 8762 23428 8795 23462
rect 8833 23428 8864 23462
rect 8864 23428 8867 23462
rect 8905 23428 8932 23462
rect 8932 23428 8939 23462
rect 8977 23428 9000 23462
rect 9000 23428 9011 23462
rect 9049 23428 9068 23462
rect 9068 23428 9083 23462
rect 9121 23428 9136 23462
rect 9136 23428 9155 23462
rect 9193 23428 9204 23462
rect 9204 23428 9227 23462
rect 9265 23428 9272 23462
rect 9272 23428 9299 23462
rect 9337 23428 9340 23462
rect 9340 23428 9371 23462
rect 9409 23428 9442 23462
rect 9442 23428 9443 23462
rect 9481 23428 9510 23462
rect 9510 23428 9515 23462
rect 9553 23428 9578 23462
rect 9578 23428 9587 23462
rect 9625 23428 9646 23462
rect 9646 23428 9659 23462
rect 9697 23428 9714 23462
rect 9714 23428 9731 23462
rect 9769 23428 9782 23462
rect 9782 23428 9803 23462
rect 9841 23428 9850 23462
rect 9850 23428 9875 23462
rect 9913 23428 9918 23462
rect 9918 23428 9947 23462
rect 9985 23428 9986 23462
rect 9986 23428 10019 23462
rect 10057 23428 10088 23462
rect 10088 23428 10091 23462
rect 10129 23428 10156 23462
rect 10156 23428 10163 23462
rect 10201 23428 10224 23462
rect 10224 23428 10235 23462
rect 10273 23428 10292 23462
rect 10292 23428 10307 23462
rect 10345 23428 10360 23462
rect 10360 23428 10379 23462
rect 10417 23428 10428 23462
rect 10428 23428 10451 23462
rect 10489 23428 10496 23462
rect 10496 23428 10523 23462
rect 10561 23428 10564 23462
rect 10564 23428 10595 23462
rect 10633 23428 10666 23462
rect 10666 23428 10667 23462
rect 10705 23428 10734 23462
rect 10734 23428 10739 23462
rect 10777 23428 10802 23462
rect 10802 23428 10811 23462
rect 10849 23428 10870 23462
rect 10870 23428 10883 23462
rect 10921 23428 10938 23462
rect 10938 23428 10955 23462
rect 10993 23428 11006 23462
rect 11006 23428 11027 23462
rect 11065 23428 11074 23462
rect 11074 23428 11099 23462
rect 11137 23428 11142 23462
rect 11142 23428 11171 23462
rect 11209 23428 11210 23462
rect 11210 23428 11243 23462
rect 11281 23428 11312 23462
rect 11312 23428 11315 23462
rect 11353 23428 11380 23462
rect 11380 23428 11387 23462
rect 11425 23428 11448 23462
rect 11448 23428 11459 23462
rect 11497 23428 11516 23462
rect 11516 23428 11531 23462
rect 11569 23428 11584 23462
rect 11584 23428 11603 23462
rect 11641 23428 11652 23462
rect 11652 23428 11675 23462
rect 11713 23428 11720 23462
rect 11720 23428 11747 23462
rect 11785 23428 11788 23462
rect 11788 23428 11819 23462
rect 11857 23428 11890 23462
rect 11890 23428 11891 23462
rect 11929 23428 11958 23462
rect 11958 23428 11963 23462
rect 12001 23428 12026 23462
rect 12026 23428 12035 23462
rect 12073 23428 12094 23462
rect 12094 23428 12107 23462
rect 12145 23428 12162 23462
rect 12162 23428 12179 23462
rect 12217 23428 12230 23462
rect 12230 23428 12251 23462
rect 12289 23428 12298 23462
rect 12298 23428 12323 23462
rect 12361 23428 12366 23462
rect 12366 23428 12395 23462
rect 12433 23428 12434 23462
rect 12434 23428 12467 23462
rect 12505 23428 12536 23462
rect 12536 23428 12539 23462
rect 12577 23428 12604 23462
rect 12604 23428 12611 23462
rect 12649 23428 12672 23462
rect 12672 23428 12683 23462
rect 12721 23428 12740 23462
rect 12740 23428 12755 23462
rect 12793 23428 12808 23462
rect 12808 23428 12827 23462
rect 12865 23428 12876 23462
rect 12876 23428 12899 23462
rect 12937 23428 12944 23462
rect 12944 23428 12971 23462
rect 13009 23428 13012 23462
rect 13012 23428 13043 23462
rect 13081 23428 13114 23462
rect 13114 23428 13115 23462
rect 13153 23428 13182 23462
rect 13182 23428 13187 23462
rect 13225 23428 13250 23462
rect 13250 23428 13259 23462
rect 13297 23428 13331 23462
rect 4727 23076 4761 23110
rect 4727 23003 4761 23037
rect 4727 22930 4761 22964
rect 4727 22857 4761 22891
rect 4727 22784 4761 22818
rect 4727 22711 4761 22745
rect 4727 22638 4761 22672
rect 4727 22565 4761 22599
rect 4727 22492 4761 22526
rect 4727 22419 4761 22453
rect 4727 22346 4761 22380
rect 4727 22272 4761 22306
rect 4727 22198 4761 22232
rect 4727 22124 4761 22158
rect 5073 23032 5107 23066
rect 5073 22959 5107 22993
rect 5073 22886 5107 22920
rect 5073 22813 5107 22847
rect 5073 22740 5107 22774
rect 5073 22667 5107 22701
rect 5073 22594 5107 22628
rect 5073 22522 5107 22556
rect 5073 22450 5107 22484
rect 5073 22378 5107 22412
rect 5073 22306 5107 22340
rect 5073 22234 5107 22268
rect 5073 22162 5107 22196
rect 5073 22090 5107 22124
rect 6718 23020 6752 23054
rect 6718 22942 6752 22976
rect 6718 22864 6752 22898
rect 6718 22786 6752 22820
rect 6718 22708 6752 22742
rect 6718 22630 6752 22664
rect 6718 22552 6752 22586
rect 6718 22475 6752 22509
rect 6718 22398 6752 22432
rect 6718 22321 6752 22355
rect 6718 22244 6752 22278
rect 6718 22167 6752 22201
rect 6718 22090 6752 22124
rect 8374 23020 8408 23054
rect 8374 22942 8408 22976
rect 8374 22864 8408 22898
rect 8374 22786 8408 22820
rect 8374 22708 8408 22742
rect 8374 22630 8408 22664
rect 8374 22552 8408 22586
rect 8374 22475 8408 22509
rect 8374 22398 8408 22432
rect 8374 22321 8408 22355
rect 8374 22244 8408 22278
rect 8374 22167 8408 22201
rect 8374 22090 8408 22124
rect 10030 23020 10064 23054
rect 10030 22942 10064 22976
rect 10030 22864 10064 22898
rect 10030 22786 10064 22820
rect 10030 22708 10064 22742
rect 10030 22630 10064 22664
rect 10030 22552 10064 22586
rect 10030 22475 10064 22509
rect 10030 22398 10064 22432
rect 10030 22321 10064 22355
rect 10030 22244 10064 22278
rect 10030 22167 10064 22201
rect 10030 22090 10064 22124
rect 11686 23020 11720 23054
rect 11686 22942 11720 22976
rect 11686 22864 11720 22898
rect 11686 22786 11720 22820
rect 11686 22708 11720 22742
rect 11686 22630 11720 22664
rect 11686 22552 11720 22586
rect 11686 22475 11720 22509
rect 11686 22398 11720 22432
rect 11686 22321 11720 22355
rect 11686 22244 11720 22278
rect 11686 22167 11720 22201
rect 11686 22090 11720 22124
rect 13342 23020 13376 23054
rect 13342 22942 13376 22976
rect 13342 22864 13376 22898
rect 13342 22786 13376 22820
rect 13342 22708 13376 22742
rect 13342 22630 13376 22664
rect 13342 22552 13376 22586
rect 13342 22475 13376 22509
rect 13342 22398 13376 22432
rect 13342 22321 13376 22355
rect 13342 22244 13376 22278
rect 13342 22167 13376 22201
rect 13342 22090 13376 22124
rect 13521 22217 13617 39027
rect 13617 22217 13699 39099
rect 13521 22144 13555 22178
rect 13593 22144 13617 22178
rect 13617 22144 13627 22178
rect 13665 22144 13699 22178
rect 4727 22050 4761 22084
rect 4727 21976 4761 22010
rect 13521 22071 13555 22105
rect 13593 22071 13617 22105
rect 13617 22071 13627 22105
rect 13665 22071 13699 22105
rect 13521 21998 13555 22032
rect 13593 21998 13617 22032
rect 13617 21998 13627 22032
rect 13665 21998 13699 22032
rect 13521 21925 13555 21959
rect 13593 21925 13617 21959
rect 13617 21925 13627 21959
rect 13665 21925 13699 21959
rect 13521 21852 13555 21886
rect 13593 21852 13617 21886
rect 13617 21852 13627 21886
rect 13665 21852 13699 21886
rect 13521 21779 13555 21813
rect 13593 21779 13617 21813
rect 13617 21779 13627 21813
rect 13665 21779 13699 21813
rect 5079 21729 5090 21763
rect 5090 21729 5113 21763
rect 5152 21729 5158 21763
rect 5158 21729 5186 21763
rect 5225 21729 5226 21763
rect 5226 21729 5259 21763
rect 5298 21729 5328 21763
rect 5328 21729 5332 21763
rect 5371 21729 5396 21763
rect 5396 21729 5405 21763
rect 5444 21729 5464 21763
rect 5464 21729 5478 21763
rect 5517 21729 5532 21763
rect 5532 21729 5551 21763
rect 5590 21729 5600 21763
rect 5600 21729 5624 21763
rect 5663 21729 5668 21763
rect 5668 21729 5697 21763
rect 5736 21729 5770 21763
rect 5809 21729 5838 21763
rect 5838 21729 5843 21763
rect 5881 21729 5906 21763
rect 5906 21729 5915 21763
rect 5953 21729 5974 21763
rect 5974 21729 5987 21763
rect 6025 21729 6042 21763
rect 6042 21729 6059 21763
rect 6097 21729 6110 21763
rect 6110 21729 6131 21763
rect 6169 21729 6178 21763
rect 6178 21729 6203 21763
rect 6241 21729 6246 21763
rect 6246 21729 6275 21763
rect 6313 21729 6314 21763
rect 6314 21729 6347 21763
rect 6385 21729 6416 21763
rect 6416 21729 6419 21763
rect 6457 21729 6484 21763
rect 6484 21729 6491 21763
rect 6529 21729 6552 21763
rect 6552 21729 6563 21763
rect 6601 21729 6620 21763
rect 6620 21729 6635 21763
rect 6673 21729 6688 21763
rect 6688 21729 6707 21763
rect 6745 21729 6756 21763
rect 6756 21729 6779 21763
rect 6817 21729 6824 21763
rect 6824 21729 6851 21763
rect 6889 21729 6892 21763
rect 6892 21729 6923 21763
rect 6961 21729 6994 21763
rect 6994 21729 6995 21763
rect 7033 21729 7062 21763
rect 7062 21729 7067 21763
rect 7105 21729 7130 21763
rect 7130 21729 7139 21763
rect 7177 21729 7198 21763
rect 7198 21729 7211 21763
rect 7249 21729 7266 21763
rect 7266 21729 7283 21763
rect 7321 21729 7334 21763
rect 7334 21729 7355 21763
rect 7393 21729 7402 21763
rect 7402 21729 7427 21763
rect 7465 21729 7470 21763
rect 7470 21729 7499 21763
rect 7537 21729 7538 21763
rect 7538 21729 7571 21763
rect 7609 21729 7640 21763
rect 7640 21729 7643 21763
rect 7681 21729 7708 21763
rect 7708 21729 7715 21763
rect 7753 21729 7776 21763
rect 7776 21729 7787 21763
rect 7825 21729 7844 21763
rect 7844 21729 7859 21763
rect 7897 21729 7912 21763
rect 7912 21729 7931 21763
rect 7969 21729 7980 21763
rect 7980 21729 8003 21763
rect 8041 21729 8048 21763
rect 8048 21729 8075 21763
rect 8113 21729 8116 21763
rect 8116 21729 8147 21763
rect 8185 21729 8218 21763
rect 8218 21729 8219 21763
rect 8257 21729 8286 21763
rect 8286 21729 8291 21763
rect 8329 21729 8354 21763
rect 8354 21729 8363 21763
rect 8401 21729 8422 21763
rect 8422 21729 8435 21763
rect 8473 21729 8490 21763
rect 8490 21729 8507 21763
rect 8545 21729 8558 21763
rect 8558 21729 8579 21763
rect 8617 21729 8626 21763
rect 8626 21729 8651 21763
rect 8689 21729 8694 21763
rect 8694 21729 8723 21763
rect 8761 21729 8762 21763
rect 8762 21729 8795 21763
rect 8833 21729 8864 21763
rect 8864 21729 8867 21763
rect 8905 21729 8932 21763
rect 8932 21729 8939 21763
rect 8977 21729 9000 21763
rect 9000 21729 9011 21763
rect 9049 21729 9068 21763
rect 9068 21729 9083 21763
rect 9121 21729 9136 21763
rect 9136 21729 9155 21763
rect 9193 21729 9204 21763
rect 9204 21729 9227 21763
rect 9265 21729 9272 21763
rect 9272 21729 9299 21763
rect 9337 21729 9340 21763
rect 9340 21729 9371 21763
rect 9409 21729 9442 21763
rect 9442 21729 9443 21763
rect 9481 21729 9510 21763
rect 9510 21729 9515 21763
rect 9553 21729 9578 21763
rect 9578 21729 9587 21763
rect 9625 21729 9646 21763
rect 9646 21729 9659 21763
rect 9697 21729 9714 21763
rect 9714 21729 9731 21763
rect 9769 21729 9782 21763
rect 9782 21729 9803 21763
rect 9841 21729 9850 21763
rect 9850 21729 9875 21763
rect 9913 21729 9918 21763
rect 9918 21729 9947 21763
rect 9985 21729 9986 21763
rect 9986 21729 10019 21763
rect 10057 21729 10088 21763
rect 10088 21729 10091 21763
rect 10129 21729 10156 21763
rect 10156 21729 10163 21763
rect 10201 21729 10224 21763
rect 10224 21729 10235 21763
rect 10273 21729 10292 21763
rect 10292 21729 10307 21763
rect 10345 21729 10360 21763
rect 10360 21729 10379 21763
rect 10417 21729 10428 21763
rect 10428 21729 10451 21763
rect 10489 21729 10496 21763
rect 10496 21729 10523 21763
rect 10561 21729 10564 21763
rect 10564 21729 10595 21763
rect 10633 21729 10666 21763
rect 10666 21729 10667 21763
rect 10705 21729 10734 21763
rect 10734 21729 10739 21763
rect 10777 21729 10802 21763
rect 10802 21729 10811 21763
rect 10849 21729 10870 21763
rect 10870 21729 10883 21763
rect 10921 21729 10938 21763
rect 10938 21729 10955 21763
rect 10993 21729 11006 21763
rect 11006 21729 11027 21763
rect 11065 21729 11074 21763
rect 11074 21729 11099 21763
rect 11137 21729 11142 21763
rect 11142 21729 11171 21763
rect 11209 21729 11210 21763
rect 11210 21729 11243 21763
rect 11281 21729 11312 21763
rect 11312 21729 11315 21763
rect 11353 21729 11380 21763
rect 11380 21729 11387 21763
rect 11425 21729 11448 21763
rect 11448 21729 11459 21763
rect 11497 21729 11516 21763
rect 11516 21729 11531 21763
rect 11569 21729 11584 21763
rect 11584 21729 11603 21763
rect 11641 21729 11652 21763
rect 11652 21729 11675 21763
rect 11713 21729 11720 21763
rect 11720 21729 11747 21763
rect 11785 21729 11788 21763
rect 11788 21729 11819 21763
rect 11857 21729 11890 21763
rect 11890 21729 11891 21763
rect 11929 21729 11958 21763
rect 11958 21729 11963 21763
rect 12001 21729 12026 21763
rect 12026 21729 12035 21763
rect 12073 21729 12094 21763
rect 12094 21729 12107 21763
rect 12145 21729 12162 21763
rect 12162 21729 12179 21763
rect 12217 21729 12230 21763
rect 12230 21729 12251 21763
rect 12289 21729 12298 21763
rect 12298 21729 12323 21763
rect 12361 21729 12366 21763
rect 12366 21729 12395 21763
rect 12433 21729 12434 21763
rect 12434 21729 12467 21763
rect 12505 21729 12536 21763
rect 12536 21729 12539 21763
rect 12577 21729 12604 21763
rect 12604 21729 12611 21763
rect 12649 21729 12672 21763
rect 12672 21729 12683 21763
rect 12721 21729 12740 21763
rect 12740 21729 12755 21763
rect 12793 21729 12808 21763
rect 12808 21729 12827 21763
rect 12865 21729 12876 21763
rect 12876 21729 12899 21763
rect 12937 21729 12944 21763
rect 12944 21729 12971 21763
rect 13009 21729 13012 21763
rect 13012 21729 13043 21763
rect 13081 21729 13114 21763
rect 13114 21729 13115 21763
rect 13153 21729 13182 21763
rect 13182 21729 13187 21763
rect 13225 21729 13250 21763
rect 13250 21729 13259 21763
rect 13297 21729 13331 21763
rect 13521 21706 13555 21740
rect 13593 21706 13617 21740
rect 13617 21706 13627 21740
rect 13665 21706 13699 21740
rect 4727 21601 4761 21635
rect 4727 21527 4761 21561
rect 4727 21453 4761 21487
rect 4727 21379 4761 21413
rect 4727 21305 4761 21339
rect 4727 21231 4761 21265
rect 13521 21633 13555 21667
rect 13593 21633 13617 21667
rect 13617 21633 13627 21667
rect 13665 21633 13699 21667
rect 13521 21560 13555 21594
rect 13593 21560 13617 21594
rect 13617 21560 13627 21594
rect 13665 21560 13699 21594
rect 13521 21487 13555 21521
rect 13593 21487 13617 21521
rect 13617 21487 13627 21521
rect 13665 21487 13699 21521
rect 13521 21414 13555 21448
rect 13593 21414 13617 21448
rect 13617 21414 13627 21448
rect 13665 21414 13699 21448
rect 13521 21341 13555 21375
rect 13593 21341 13617 21375
rect 13617 21341 13627 21375
rect 13665 21341 13699 21375
rect 13521 21268 13555 21302
rect 13593 21268 13617 21302
rect 13617 21268 13627 21302
rect 13665 21268 13699 21302
rect 4727 21157 4761 21191
rect 4727 21083 4761 21117
rect 4727 21009 4761 21043
rect 4727 20935 4761 20969
rect 4727 20861 4761 20895
rect 4727 20788 4761 20822
rect 4727 20715 4761 20749
rect 4727 20642 4761 20676
rect 4727 20569 4761 20603
rect 4727 20496 4761 20530
rect 4727 20423 4761 20457
rect 4727 20350 4761 20384
rect 4727 20277 4761 20311
rect 5073 21217 5107 21251
rect 5073 21144 5107 21178
rect 5073 21071 5107 21105
rect 5073 20998 5107 21032
rect 5073 20925 5107 20959
rect 5073 20853 5107 20887
rect 5073 20781 5107 20815
rect 5073 20709 5107 20743
rect 5073 20637 5107 20671
rect 5073 20565 5107 20599
rect 5073 20493 5107 20527
rect 5073 20421 5107 20455
rect 5073 20349 5107 20383
rect 5073 20277 5107 20311
rect 6718 21217 6752 21251
rect 6718 21144 6752 21178
rect 6718 21071 6752 21105
rect 6718 20998 6752 21032
rect 6718 20925 6752 20959
rect 6718 20853 6752 20887
rect 6718 20781 6752 20815
rect 6718 20709 6752 20743
rect 6718 20637 6752 20671
rect 6718 20565 6752 20599
rect 6718 20493 6752 20527
rect 6718 20421 6752 20455
rect 6718 20349 6752 20383
rect 6718 20277 6752 20311
rect 8374 21217 8408 21251
rect 8374 21144 8408 21178
rect 8374 21071 8408 21105
rect 8374 20998 8408 21032
rect 8374 20925 8408 20959
rect 8374 20853 8408 20887
rect 8374 20781 8408 20815
rect 8374 20709 8408 20743
rect 8374 20637 8408 20671
rect 8374 20565 8408 20599
rect 8374 20493 8408 20527
rect 8374 20421 8408 20455
rect 8374 20349 8408 20383
rect 8374 20277 8408 20311
rect 10030 21217 10064 21251
rect 10030 21144 10064 21178
rect 10030 21071 10064 21105
rect 10030 20998 10064 21032
rect 10030 20925 10064 20959
rect 10030 20853 10064 20887
rect 10030 20781 10064 20815
rect 10030 20709 10064 20743
rect 10030 20637 10064 20671
rect 10030 20565 10064 20599
rect 10030 20493 10064 20527
rect 10030 20421 10064 20455
rect 10030 20349 10064 20383
rect 10030 20277 10064 20311
rect 11686 21217 11720 21251
rect 11686 21144 11720 21178
rect 11686 21071 11720 21105
rect 11686 20998 11720 21032
rect 11686 20925 11720 20959
rect 11686 20853 11720 20887
rect 11686 20781 11720 20815
rect 11686 20709 11720 20743
rect 11686 20637 11720 20671
rect 11686 20565 11720 20599
rect 11686 20493 11720 20527
rect 11686 20421 11720 20455
rect 11686 20349 11720 20383
rect 11686 20277 11720 20311
rect 13342 21217 13376 21251
rect 13342 21144 13376 21178
rect 13342 21071 13376 21105
rect 13342 20998 13376 21032
rect 13342 20925 13376 20959
rect 13342 20853 13376 20887
rect 13342 20781 13376 20815
rect 13342 20709 13376 20743
rect 13342 20637 13376 20671
rect 13342 20565 13376 20599
rect 13342 20493 13376 20527
rect 13342 20421 13376 20455
rect 13342 20349 13376 20383
rect 13342 20277 13376 20311
rect 13521 21195 13555 21229
rect 13593 21195 13617 21229
rect 13617 21195 13627 21229
rect 13665 21195 13699 21229
rect 13521 21122 13555 21156
rect 13593 21122 13617 21156
rect 13617 21122 13627 21156
rect 13665 21122 13699 21156
rect 13521 21049 13555 21083
rect 13593 21049 13617 21083
rect 13617 21049 13627 21083
rect 13665 21049 13699 21083
rect 13521 20976 13555 21010
rect 13593 20976 13617 21010
rect 13617 20976 13627 21010
rect 13665 20976 13699 21010
rect 13521 20903 13555 20937
rect 13593 20903 13617 20937
rect 13617 20903 13627 20937
rect 13665 20903 13699 20937
rect 13521 20830 13555 20864
rect 13593 20830 13617 20864
rect 13617 20830 13627 20864
rect 13665 20830 13699 20864
rect 13521 20757 13555 20791
rect 13593 20757 13617 20791
rect 13617 20757 13627 20791
rect 13665 20757 13699 20791
rect 13521 20684 13555 20718
rect 13593 20684 13617 20718
rect 13617 20684 13627 20718
rect 13665 20684 13699 20718
rect 13521 20611 13555 20645
rect 13593 20611 13617 20645
rect 13617 20611 13627 20645
rect 13665 20611 13699 20645
rect 13521 20538 13555 20572
rect 13593 20538 13617 20572
rect 13617 20538 13627 20572
rect 13665 20538 13699 20572
rect 13521 20496 13555 20499
rect 13593 20496 13627 20499
rect 13521 20465 13549 20496
rect 13549 20465 13555 20496
rect 13593 20465 13617 20496
rect 13617 20465 13627 20496
rect 13665 20465 13699 20499
rect 13521 20393 13549 20426
rect 13549 20393 13555 20426
rect 13593 20393 13617 20426
rect 13617 20393 13627 20426
rect 13521 20392 13555 20393
rect 13593 20392 13627 20393
rect 13665 20392 13699 20426
rect 13521 20324 13549 20353
rect 13549 20324 13555 20353
rect 13593 20324 13617 20353
rect 13617 20324 13627 20353
rect 13521 20319 13555 20324
rect 13593 20319 13627 20324
rect 13665 20319 13699 20353
rect 13521 20255 13549 20280
rect 13549 20255 13555 20280
rect 13593 20255 13617 20280
rect 13617 20255 13627 20280
rect 13521 20246 13555 20255
rect 13593 20246 13627 20255
rect 13665 20246 13699 20280
rect 13521 20173 13525 20207
rect 13525 20173 13555 20207
rect 13593 20173 13627 20207
rect 13665 20173 13699 20207
rect 13838 26620 13840 39287
rect 13840 26620 13942 39287
rect 13942 26620 13944 39287
rect 13838 26547 13840 26581
rect 13840 26547 13872 26581
rect 13910 26547 13942 26581
rect 13942 26547 13944 26581
rect 13838 26474 13840 26508
rect 13840 26474 13872 26508
rect 13910 26474 13942 26508
rect 13942 26474 13944 26508
rect 13838 26401 13840 26435
rect 13840 26401 13872 26435
rect 13910 26401 13942 26435
rect 13942 26401 13944 26435
rect 13838 26328 13840 26362
rect 13840 26328 13872 26362
rect 13910 26328 13942 26362
rect 13942 26328 13944 26362
rect 13838 26255 13840 26289
rect 13840 26255 13872 26289
rect 13910 26255 13942 26289
rect 13942 26255 13944 26289
rect 13838 26182 13840 26216
rect 13840 26182 13872 26216
rect 13910 26182 13942 26216
rect 13942 26182 13944 26216
rect 13838 26109 13840 26143
rect 13840 26109 13872 26143
rect 13910 26109 13942 26143
rect 13942 26109 13944 26143
rect 13838 26036 13840 26070
rect 13840 26036 13872 26070
rect 13910 26036 13942 26070
rect 13942 26036 13944 26070
rect 13838 25963 13840 25997
rect 13840 25963 13872 25997
rect 13910 25963 13942 25997
rect 13942 25963 13944 25997
rect 13838 25890 13840 25924
rect 13840 25890 13872 25924
rect 13910 25890 13942 25924
rect 13942 25890 13944 25924
rect 13838 25817 13840 25851
rect 13840 25817 13872 25851
rect 13910 25817 13942 25851
rect 13942 25817 13944 25851
rect 13838 25744 13840 25778
rect 13840 25744 13872 25778
rect 13910 25744 13942 25778
rect 13942 25744 13944 25778
rect 13838 25671 13840 25705
rect 13840 25671 13872 25705
rect 13910 25671 13942 25705
rect 13942 25671 13944 25705
rect 13838 25598 13840 25632
rect 13840 25598 13872 25632
rect 13910 25598 13942 25632
rect 13942 25598 13944 25632
rect 13838 25525 13840 25559
rect 13840 25525 13872 25559
rect 13910 25525 13942 25559
rect 13942 25525 13944 25559
rect 13838 25452 13840 25486
rect 13840 25452 13872 25486
rect 13910 25452 13942 25486
rect 13942 25452 13944 25486
rect 13838 25379 13840 25413
rect 13840 25379 13872 25413
rect 13910 25379 13942 25413
rect 13942 25379 13944 25413
rect 13838 25306 13840 25340
rect 13840 25306 13872 25340
rect 13910 25306 13942 25340
rect 13942 25306 13944 25340
rect 13838 25233 13840 25267
rect 13840 25233 13872 25267
rect 13910 25233 13942 25267
rect 13942 25233 13944 25267
rect 13838 25160 13840 25194
rect 13840 25160 13872 25194
rect 13910 25160 13942 25194
rect 13942 25160 13944 25194
rect 13838 25087 13840 25121
rect 13840 25087 13872 25121
rect 13910 25087 13942 25121
rect 13942 25087 13944 25121
rect 13838 25014 13840 25048
rect 13840 25014 13872 25048
rect 13910 25014 13942 25048
rect 13942 25014 13944 25048
rect 13838 24941 13840 24975
rect 13840 24941 13872 24975
rect 13910 24941 13942 24975
rect 13942 24941 13944 24975
rect 13838 24868 13840 24902
rect 13840 24868 13872 24902
rect 13910 24868 13942 24902
rect 13942 24868 13944 24902
rect 13838 24795 13840 24829
rect 13840 24795 13872 24829
rect 13910 24795 13942 24829
rect 13942 24795 13944 24829
rect 13838 24722 13840 24756
rect 13840 24722 13872 24756
rect 13910 24722 13942 24756
rect 13942 24722 13944 24756
rect 13838 24649 13840 24683
rect 13840 24649 13872 24683
rect 13910 24649 13942 24683
rect 13942 24649 13944 24683
rect 13838 24576 13840 24610
rect 13840 24576 13872 24610
rect 13910 24576 13942 24610
rect 13942 24576 13944 24610
rect 13838 24503 13840 24537
rect 13840 24503 13872 24537
rect 13910 24503 13942 24537
rect 13942 24503 13944 24537
rect 13838 24430 13840 24464
rect 13840 24430 13872 24464
rect 13910 24430 13942 24464
rect 13942 24430 13944 24464
rect 13838 24357 13840 24391
rect 13840 24357 13872 24391
rect 13910 24357 13942 24391
rect 13942 24357 13944 24391
rect 13838 24284 13840 24318
rect 13840 24284 13872 24318
rect 13910 24284 13942 24318
rect 13942 24284 13944 24318
rect 13838 24211 13840 24245
rect 13840 24211 13872 24245
rect 13910 24211 13942 24245
rect 13942 24211 13944 24245
rect 13838 24138 13840 24172
rect 13840 24138 13872 24172
rect 13910 24138 13942 24172
rect 13942 24138 13944 24172
rect 13838 24065 13840 24099
rect 13840 24065 13872 24099
rect 13910 24065 13942 24099
rect 13942 24065 13944 24099
rect 13838 23992 13840 24026
rect 13840 23992 13872 24026
rect 13910 23992 13942 24026
rect 13942 23992 13944 24026
rect 13838 23919 13840 23953
rect 13840 23919 13872 23953
rect 13910 23919 13942 23953
rect 13942 23919 13944 23953
rect 13838 23846 13840 23880
rect 13840 23846 13872 23880
rect 13910 23846 13942 23880
rect 13942 23846 13944 23880
rect 13838 23773 13840 23807
rect 13840 23773 13872 23807
rect 13910 23773 13942 23807
rect 13942 23773 13944 23807
rect 13838 23700 13840 23734
rect 13840 23700 13872 23734
rect 13910 23700 13942 23734
rect 13942 23700 13944 23734
rect 13838 23627 13840 23661
rect 13840 23627 13872 23661
rect 13910 23627 13942 23661
rect 13942 23627 13944 23661
rect 13838 23554 13840 23588
rect 13840 23554 13872 23588
rect 13910 23554 13942 23588
rect 13942 23554 13944 23588
rect 13838 23481 13840 23515
rect 13840 23481 13872 23515
rect 13910 23481 13942 23515
rect 13942 23481 13944 23515
rect 13838 23408 13840 23442
rect 13840 23408 13872 23442
rect 13910 23408 13942 23442
rect 13942 23408 13944 23442
rect 13838 23335 13840 23369
rect 13840 23335 13872 23369
rect 13910 23335 13942 23369
rect 13942 23335 13944 23369
rect 13838 23262 13840 23296
rect 13840 23262 13872 23296
rect 13910 23262 13942 23296
rect 13942 23262 13944 23296
rect 13838 23189 13840 23223
rect 13840 23189 13872 23223
rect 13910 23189 13942 23223
rect 13942 23189 13944 23223
rect 13838 23116 13840 23150
rect 13840 23116 13872 23150
rect 13910 23116 13942 23150
rect 13942 23116 13944 23150
rect 13838 23043 13840 23077
rect 13840 23043 13872 23077
rect 13910 23043 13942 23077
rect 13942 23043 13944 23077
rect 13838 22970 13840 23004
rect 13840 22970 13872 23004
rect 13910 22970 13942 23004
rect 13942 22970 13944 23004
rect 13838 22897 13840 22931
rect 13840 22897 13872 22931
rect 13910 22897 13942 22931
rect 13942 22897 13944 22931
rect 13838 22824 13840 22858
rect 13840 22824 13872 22858
rect 13910 22824 13942 22858
rect 13942 22824 13944 22858
rect 13838 22751 13840 22785
rect 13840 22751 13872 22785
rect 13910 22751 13942 22785
rect 13942 22751 13944 22785
rect 13838 22678 13840 22712
rect 13840 22678 13872 22712
rect 13910 22678 13942 22712
rect 13942 22678 13944 22712
rect 13838 22605 13840 22639
rect 13840 22605 13872 22639
rect 13910 22605 13942 22639
rect 13942 22605 13944 22639
rect 13838 22532 13840 22566
rect 13840 22532 13872 22566
rect 13910 22532 13942 22566
rect 13942 22532 13944 22566
rect 13838 22459 13840 22493
rect 13840 22459 13872 22493
rect 13910 22459 13942 22493
rect 13942 22459 13944 22493
rect 13838 22386 13840 22420
rect 13840 22386 13872 22420
rect 13910 22386 13942 22420
rect 13942 22386 13944 22420
rect 13838 22313 13840 22347
rect 13840 22313 13872 22347
rect 13910 22313 13942 22347
rect 13942 22313 13944 22347
rect 13838 22240 13840 22274
rect 13840 22240 13872 22274
rect 13910 22240 13942 22274
rect 13942 22240 13944 22274
rect 13838 22167 13840 22201
rect 13840 22167 13872 22201
rect 13910 22167 13942 22201
rect 13942 22167 13944 22201
rect 13838 22094 13840 22128
rect 13840 22094 13872 22128
rect 13910 22094 13942 22128
rect 13942 22094 13944 22128
rect 13838 22021 13840 22055
rect 13840 22021 13872 22055
rect 13910 22021 13942 22055
rect 13942 22021 13944 22055
rect 13838 21948 13840 21982
rect 13840 21948 13872 21982
rect 13910 21948 13942 21982
rect 13942 21948 13944 21982
rect 13838 21875 13840 21909
rect 13840 21875 13872 21909
rect 13910 21875 13942 21909
rect 13942 21875 13944 21909
rect 13838 21802 13840 21836
rect 13840 21802 13872 21836
rect 13910 21802 13942 21836
rect 13942 21802 13944 21836
rect 13838 21729 13840 21763
rect 13840 21729 13872 21763
rect 13910 21729 13942 21763
rect 13942 21729 13944 21763
rect 13838 21656 13840 21690
rect 13840 21656 13872 21690
rect 13910 21656 13942 21690
rect 13942 21656 13944 21690
rect 13838 21583 13840 21617
rect 13840 21583 13872 21617
rect 13910 21583 13942 21617
rect 13942 21583 13944 21617
rect 13838 21510 13840 21544
rect 13840 21510 13872 21544
rect 13910 21510 13942 21544
rect 13942 21510 13944 21544
rect 13838 21437 13840 21471
rect 13840 21437 13872 21471
rect 13910 21437 13942 21471
rect 13942 21437 13944 21471
rect 1943 19443 1946 19477
rect 1946 19443 1977 19477
rect 2015 19443 2048 19477
rect 2048 19443 2049 19477
rect 1943 19369 1946 19403
rect 1946 19369 1977 19403
rect 2015 19369 2048 19403
rect 2048 19369 2049 19403
rect 1943 19295 1946 19329
rect 1946 19295 1977 19329
rect 2015 19295 2048 19329
rect 2048 19295 2049 19329
rect 1943 19221 1946 19255
rect 1946 19221 1977 19255
rect 2015 19221 2048 19255
rect 2048 19221 2049 19255
rect 1943 19147 1946 19181
rect 1946 19147 1977 19181
rect 2015 19147 2048 19181
rect 2048 19147 2049 19181
rect 1943 19073 1946 19107
rect 1946 19073 1977 19107
rect 2015 19073 2048 19107
rect 2048 19073 2049 19107
rect 1943 18999 1946 19033
rect 1946 18999 1977 19033
rect 2015 18999 2048 19033
rect 2048 18999 2049 19033
rect 1943 18925 1946 18959
rect 1946 18925 1977 18959
rect 2015 18925 2048 18959
rect 2048 18925 2049 18959
rect 1943 18850 1946 18884
rect 1946 18850 1977 18884
rect 2015 18850 2048 18884
rect 2048 18850 2049 18884
rect 1943 18775 1946 18809
rect 1946 18775 1977 18809
rect 2015 18775 2048 18809
rect 2048 18775 2049 18809
rect 1943 18700 1946 18734
rect 1946 18700 1977 18734
rect 2015 18700 2048 18734
rect 2048 18700 2049 18734
rect 1943 18625 1946 18659
rect 1946 18625 1977 18659
rect 2015 18625 2048 18659
rect 2048 18625 2049 18659
rect 1943 18550 1946 18584
rect 1946 18550 1977 18584
rect 2015 18550 2048 18584
rect 2048 18550 2049 18584
rect 1943 18475 1946 18509
rect 1946 18475 1977 18509
rect 2015 18475 2048 18509
rect 2048 18475 2049 18509
rect 1943 18400 1946 18434
rect 1946 18400 1977 18434
rect 2015 18400 2048 18434
rect 2048 18400 2049 18434
rect 1943 18325 1946 18359
rect 1946 18325 1977 18359
rect 2015 18325 2048 18359
rect 2048 18325 2049 18359
rect 1943 18250 1946 18284
rect 1946 18250 1977 18284
rect 2015 18250 2048 18284
rect 2048 18250 2049 18284
rect 1943 18175 1946 18209
rect 1946 18175 1977 18209
rect 2015 18175 2048 18209
rect 2048 18175 2049 18209
rect 1943 18100 1946 18134
rect 1946 18100 1977 18134
rect 2015 18100 2048 18134
rect 2048 18100 2049 18134
rect 1943 18025 1946 18059
rect 1946 18025 1977 18059
rect 2015 18025 2048 18059
rect 2048 18025 2049 18059
rect 1943 17950 1946 17984
rect 1946 17950 1977 17984
rect 2015 17950 2048 17984
rect 2048 17950 2049 17984
rect 1943 17875 1946 17909
rect 1946 17875 1977 17909
rect 2015 17875 2048 17909
rect 2048 17875 2049 17909
rect 4923 19708 4943 19742
rect 4943 19708 4957 19742
rect 4996 19708 5011 19742
rect 5011 19708 5030 19742
rect 5069 19708 5079 19742
rect 5079 19708 5103 19742
rect 5142 19708 5147 19742
rect 5147 19708 5176 19742
rect 5215 19708 5249 19742
rect 5288 19708 5317 19742
rect 5317 19708 5322 19742
rect 5361 19708 5385 19742
rect 5385 19708 5395 19742
rect 5434 19708 5453 19742
rect 5453 19708 5468 19742
rect 5507 19708 5521 19742
rect 5521 19708 5541 19742
rect 5580 19708 5589 19742
rect 5589 19708 5614 19742
rect 5653 19708 5657 19742
rect 5657 19708 5687 19742
rect 5726 19708 5759 19742
rect 5759 19708 5760 19742
rect 5799 19708 5827 19742
rect 5827 19708 5833 19742
rect 5872 19708 5895 19742
rect 5895 19708 5906 19742
rect 5945 19708 5963 19742
rect 5963 19708 5979 19742
rect 6017 19708 6031 19742
rect 6031 19708 6051 19742
rect 6089 19708 6099 19742
rect 6099 19708 6123 19742
rect 6161 19708 6167 19742
rect 6167 19708 6195 19742
rect 6233 19708 6235 19742
rect 6235 19708 6267 19742
rect 6305 19708 6337 19742
rect 6337 19708 6339 19742
rect 6377 19708 6405 19742
rect 6405 19708 6411 19742
rect 6449 19708 6473 19742
rect 6473 19708 6483 19742
rect 6521 19708 6541 19742
rect 6541 19708 6555 19742
rect 6593 19708 6609 19742
rect 6609 19708 6627 19742
rect 6665 19708 6677 19742
rect 6677 19708 6699 19742
rect 6737 19708 6745 19742
rect 6745 19708 6771 19742
rect 6809 19708 6813 19742
rect 6813 19708 6843 19742
rect 6881 19708 6915 19742
rect 6953 19708 6983 19742
rect 6983 19708 6987 19742
rect 7025 19708 7051 19742
rect 7051 19708 7059 19742
rect 7097 19708 7119 19742
rect 7119 19708 7131 19742
rect 7169 19708 7187 19742
rect 7187 19708 7203 19742
rect 7241 19708 7255 19742
rect 7255 19708 7275 19742
rect 7313 19708 7323 19742
rect 7323 19708 7347 19742
rect 7385 19708 7391 19742
rect 7391 19708 7419 19742
rect 7457 19708 7459 19742
rect 7459 19708 7491 19742
rect 7529 19708 7561 19742
rect 7561 19708 7563 19742
rect 7601 19708 7629 19742
rect 7629 19708 7635 19742
rect 7673 19708 7697 19742
rect 7697 19708 7707 19742
rect 7745 19708 7765 19742
rect 7765 19708 7779 19742
rect 7817 19708 7833 19742
rect 7833 19708 7851 19742
rect 7889 19708 7901 19742
rect 7901 19708 7923 19742
rect 7961 19708 7969 19742
rect 7969 19708 7995 19742
rect 8033 19708 8037 19742
rect 8037 19708 8067 19742
rect 8105 19708 8139 19742
rect 8177 19708 8207 19742
rect 8207 19708 8211 19742
rect 8249 19708 8275 19742
rect 8275 19708 8283 19742
rect 8321 19708 8343 19742
rect 8343 19708 8355 19742
rect 8393 19708 8411 19742
rect 8411 19708 8427 19742
rect 8465 19708 8479 19742
rect 8479 19708 8499 19742
rect 8537 19708 8547 19742
rect 8547 19708 8571 19742
rect 8609 19708 8615 19742
rect 8615 19708 8643 19742
rect 8681 19708 8683 19742
rect 8683 19708 8715 19742
rect 8753 19708 8785 19742
rect 8785 19708 8787 19742
rect 8825 19708 8853 19742
rect 8853 19708 8859 19742
rect 8897 19708 8921 19742
rect 8921 19708 8931 19742
rect 8969 19708 8989 19742
rect 8989 19708 9003 19742
rect 9041 19708 9057 19742
rect 9057 19708 9075 19742
rect 9113 19708 9125 19742
rect 9125 19708 9147 19742
rect 9185 19708 9193 19742
rect 9193 19708 9219 19742
rect 9257 19708 9261 19742
rect 9261 19708 9291 19742
rect 9329 19708 9363 19742
rect 9401 19708 9431 19742
rect 9431 19708 9435 19742
rect 9473 19708 9499 19742
rect 9499 19708 9507 19742
rect 9545 19708 9567 19742
rect 9567 19708 9579 19742
rect 9617 19708 9635 19742
rect 9635 19708 9651 19742
rect 9689 19708 9703 19742
rect 9703 19708 9723 19742
rect 9761 19708 9771 19742
rect 9771 19708 9795 19742
rect 9833 19708 9839 19742
rect 9839 19708 9867 19742
rect 9905 19708 9907 19742
rect 9907 19708 9939 19742
rect 9977 19708 10009 19742
rect 10009 19708 10011 19742
rect 10049 19708 10077 19742
rect 10077 19708 10083 19742
rect 10121 19708 10145 19742
rect 10145 19708 10155 19742
rect 10193 19708 10213 19742
rect 10213 19708 10227 19742
rect 10265 19708 10281 19742
rect 10281 19708 10299 19742
rect 10337 19708 10349 19742
rect 10349 19708 10371 19742
rect 10409 19708 10417 19742
rect 10417 19708 10443 19742
rect 10481 19708 10485 19742
rect 10485 19708 10515 19742
rect 10553 19708 10587 19742
rect 10625 19708 10655 19742
rect 10655 19708 10659 19742
rect 10697 19708 10723 19742
rect 10723 19708 10731 19742
rect 10769 19708 10791 19742
rect 10791 19708 10803 19742
rect 10841 19708 10859 19742
rect 10859 19708 10875 19742
rect 10913 19708 10927 19742
rect 10927 19708 10947 19742
rect 10985 19708 10995 19742
rect 10995 19708 11019 19742
rect 11057 19708 11063 19742
rect 11063 19708 11091 19742
rect 11129 19708 11131 19742
rect 11131 19708 11163 19742
rect 11201 19708 11233 19742
rect 11233 19708 11235 19742
rect 11273 19708 11301 19742
rect 11301 19708 11307 19742
rect 11345 19708 11369 19742
rect 11369 19708 11379 19742
rect 11417 19708 11437 19742
rect 11437 19708 11451 19742
rect 11489 19708 11505 19742
rect 11505 19708 11523 19742
rect 11561 19708 11573 19742
rect 11573 19708 11595 19742
rect 11633 19708 11641 19742
rect 11641 19708 11667 19742
rect 11705 19708 11709 19742
rect 11709 19708 11739 19742
rect 11777 19708 11811 19742
rect 11849 19708 11879 19742
rect 11879 19708 11883 19742
rect 11921 19708 11947 19742
rect 11947 19708 11955 19742
rect 11993 19708 12015 19742
rect 12015 19708 12027 19742
rect 12065 19708 12083 19742
rect 12083 19708 12099 19742
rect 12137 19708 12151 19742
rect 12151 19708 12171 19742
rect 12209 19708 12219 19742
rect 12219 19708 12243 19742
rect 12281 19708 12287 19742
rect 12287 19708 12315 19742
rect 12353 19708 12355 19742
rect 12355 19708 12387 19742
rect 12425 19708 12457 19742
rect 12457 19708 12459 19742
rect 12497 19708 12525 19742
rect 12525 19708 12531 19742
rect 12569 19708 12593 19742
rect 12593 19708 12603 19742
rect 12641 19708 12661 19742
rect 12661 19708 12675 19742
rect 12713 19708 12729 19742
rect 12729 19708 12747 19742
rect 12785 19708 12797 19742
rect 12797 19708 12819 19742
rect 12857 19708 12865 19742
rect 12865 19708 12891 19742
rect 12929 19708 12933 19742
rect 12933 19708 12963 19742
rect 13490 19701 13596 19745
rect 2184 16883 2218 16917
rect 2258 16883 2292 16917
rect 2332 16883 2366 16917
rect 2184 16764 2218 16798
rect 2258 16764 2292 16798
rect 2332 16764 2366 16798
rect 3899 16883 3933 16917
rect 3973 16883 4007 16917
rect 4047 16883 4081 16917
rect 3899 16764 3933 16798
rect 3973 16764 4007 16798
rect 4047 16764 4081 16798
rect 4486 19544 4520 19578
rect 4622 19544 4656 19578
rect 4486 19471 4520 19505
rect 4622 19471 4656 19505
rect 4486 19398 4520 19432
rect 4622 19398 4656 19432
rect 4486 19325 4520 19359
rect 4622 19325 4656 19359
rect 4486 19252 4520 19286
rect 4622 19252 4656 19286
rect 4486 19179 4520 19213
rect 4622 19179 4656 19213
rect 4486 19106 4520 19140
rect 4622 19106 4656 19140
rect 4486 19033 4520 19067
rect 4622 19033 4656 19067
rect 4486 18960 4520 18994
rect 4622 18960 4656 18994
rect 4486 18887 4520 18921
rect 4622 18887 4656 18921
rect 4486 18814 4520 18848
rect 4622 18814 4656 18848
rect 4486 18741 4520 18775
rect 4622 18741 4656 18775
rect 4486 18668 4520 18702
rect 4622 18668 4656 18702
rect 4486 18595 4520 18629
rect 4622 18595 4656 18629
rect 4486 18522 4520 18556
rect 4622 18522 4656 18556
rect 4486 18449 4520 18483
rect 4622 18449 4656 18483
rect 4486 18376 4520 18410
rect 4622 18376 4656 18410
rect 4486 18303 4520 18337
rect 4622 18303 4656 18337
rect 4486 18230 4520 18264
rect 4622 18230 4656 18264
rect 4737 19580 4771 19614
rect 4809 19580 4843 19614
rect 4737 19506 4771 19540
rect 4809 19506 4843 19540
rect 4737 19432 4771 19466
rect 4809 19432 4843 19466
rect 4737 19358 4771 19392
rect 4809 19358 4843 19392
rect 13342 19540 13376 19574
rect 13342 19464 13376 19498
rect 13342 19388 13376 19422
rect 4737 19284 4771 19318
rect 4809 19284 4843 19318
rect 4737 19210 4771 19244
rect 4809 19210 4843 19244
rect 4737 19136 4771 19170
rect 4809 19136 4843 19170
rect 4737 19062 4771 19096
rect 4809 19062 4843 19096
rect 4737 18988 4771 19022
rect 4809 18988 4843 19022
rect 4737 18914 4771 18948
rect 4809 18914 4843 18948
rect 4737 18840 4771 18874
rect 4809 18840 4843 18874
rect 4737 18767 4771 18801
rect 4809 18767 4843 18801
rect 4737 18694 4771 18728
rect 4809 18694 4843 18728
rect 4737 18621 4771 18655
rect 4809 18621 4843 18655
rect 4737 18548 4771 18582
rect 4809 18548 4843 18582
rect 4737 18475 4771 18509
rect 4809 18475 4843 18509
rect 4737 18402 4771 18436
rect 4809 18402 4843 18436
rect 5062 19351 5096 19385
rect 5062 19276 5096 19310
rect 5062 19201 5096 19235
rect 5062 19126 5096 19160
rect 5062 19052 5096 19086
rect 5062 18978 5096 19012
rect 5062 18904 5096 18938
rect 5062 18830 5096 18864
rect 5062 18756 5096 18790
rect 5062 18682 5096 18716
rect 5062 18608 5096 18642
rect 5062 18534 5096 18568
rect 5062 18460 5096 18494
rect 5062 18386 5096 18420
rect 6718 19351 6752 19385
rect 6718 19276 6752 19310
rect 6718 19201 6752 19235
rect 6718 19126 6752 19160
rect 6718 19052 6752 19086
rect 6718 18978 6752 19012
rect 6718 18904 6752 18938
rect 6718 18830 6752 18864
rect 6718 18756 6752 18790
rect 6718 18682 6752 18716
rect 6718 18608 6752 18642
rect 6718 18534 6752 18568
rect 6718 18460 6752 18494
rect 6718 18386 6752 18420
rect 8374 19351 8408 19385
rect 8374 19276 8408 19310
rect 8374 19201 8408 19235
rect 8374 19126 8408 19160
rect 8374 19052 8408 19086
rect 8374 18978 8408 19012
rect 8374 18904 8408 18938
rect 8374 18830 8408 18864
rect 8374 18756 8408 18790
rect 8374 18682 8408 18716
rect 8374 18608 8408 18642
rect 8374 18534 8408 18568
rect 8374 18460 8408 18494
rect 8374 18386 8408 18420
rect 10030 19351 10064 19385
rect 10030 19276 10064 19310
rect 10030 19201 10064 19235
rect 10030 19126 10064 19160
rect 10030 19052 10064 19086
rect 10030 18978 10064 19012
rect 10030 18904 10064 18938
rect 10030 18830 10064 18864
rect 10030 18756 10064 18790
rect 10030 18682 10064 18716
rect 10030 18608 10064 18642
rect 10030 18534 10064 18568
rect 10030 18460 10064 18494
rect 10030 18386 10064 18420
rect 11686 19351 11720 19385
rect 11686 19276 11720 19310
rect 11686 19201 11720 19235
rect 11686 19126 11720 19160
rect 11686 19052 11720 19086
rect 11686 18978 11720 19012
rect 11686 18904 11720 18938
rect 11686 18830 11720 18864
rect 11686 18756 11720 18790
rect 11686 18682 11720 18716
rect 11686 18608 11720 18642
rect 11686 18534 11720 18568
rect 11686 18460 11720 18494
rect 11686 18386 11720 18420
rect 13342 19312 13376 19346
rect 13342 19236 13376 19270
rect 13342 19160 13376 19194
rect 13342 19084 13376 19118
rect 13342 19008 13376 19042
rect 13342 18932 13376 18966
rect 13342 18856 13376 18890
rect 13342 18781 13376 18815
rect 13342 18706 13376 18740
rect 13342 18631 13376 18665
rect 13342 18556 13376 18590
rect 13342 18481 13376 18515
rect 13342 18406 13376 18440
rect 4737 18329 4771 18363
rect 4809 18329 4843 18363
rect 4737 18256 4771 18290
rect 4809 18256 4843 18290
rect 13342 18331 13376 18365
rect 13342 18256 13376 18290
rect 4486 18157 4520 18191
rect 4622 18157 4656 18191
rect 4486 18084 4520 18118
rect 4622 18084 4656 18118
rect 4486 18011 4520 18045
rect 4622 18011 4656 18045
rect 4923 18009 4943 18043
rect 4943 18009 4957 18043
rect 4996 18009 5011 18043
rect 5011 18009 5030 18043
rect 5069 18009 5079 18043
rect 5079 18009 5103 18043
rect 5142 18009 5147 18043
rect 5147 18009 5176 18043
rect 5215 18009 5249 18043
rect 5288 18009 5317 18043
rect 5317 18009 5322 18043
rect 5361 18009 5385 18043
rect 5385 18009 5395 18043
rect 5434 18009 5453 18043
rect 5453 18009 5468 18043
rect 5507 18009 5521 18043
rect 5521 18009 5541 18043
rect 5580 18009 5589 18043
rect 5589 18009 5614 18043
rect 5653 18009 5657 18043
rect 5657 18009 5687 18043
rect 5726 18009 5759 18043
rect 5759 18009 5760 18043
rect 5799 18009 5827 18043
rect 5827 18009 5833 18043
rect 5872 18009 5895 18043
rect 5895 18009 5906 18043
rect 5945 18009 5963 18043
rect 5963 18009 5979 18043
rect 6017 18009 6031 18043
rect 6031 18009 6051 18043
rect 6089 18009 6099 18043
rect 6099 18009 6123 18043
rect 6161 18009 6167 18043
rect 6167 18009 6195 18043
rect 6233 18009 6235 18043
rect 6235 18009 6267 18043
rect 6305 18009 6337 18043
rect 6337 18009 6339 18043
rect 6377 18009 6405 18043
rect 6405 18009 6411 18043
rect 6449 18009 6473 18043
rect 6473 18009 6483 18043
rect 6521 18009 6541 18043
rect 6541 18009 6555 18043
rect 6593 18009 6609 18043
rect 6609 18009 6627 18043
rect 6665 18009 6677 18043
rect 6677 18009 6699 18043
rect 6737 18009 6745 18043
rect 6745 18009 6771 18043
rect 6809 18009 6813 18043
rect 6813 18009 6843 18043
rect 6881 18009 6915 18043
rect 6953 18009 6983 18043
rect 6983 18009 6987 18043
rect 7025 18009 7051 18043
rect 7051 18009 7059 18043
rect 7097 18009 7119 18043
rect 7119 18009 7131 18043
rect 7169 18009 7187 18043
rect 7187 18009 7203 18043
rect 7241 18009 7255 18043
rect 7255 18009 7275 18043
rect 7313 18009 7323 18043
rect 7323 18009 7347 18043
rect 7385 18009 7391 18043
rect 7391 18009 7419 18043
rect 7457 18009 7459 18043
rect 7459 18009 7491 18043
rect 7529 18009 7561 18043
rect 7561 18009 7563 18043
rect 7601 18009 7629 18043
rect 7629 18009 7635 18043
rect 7673 18009 7697 18043
rect 7697 18009 7707 18043
rect 7745 18009 7765 18043
rect 7765 18009 7779 18043
rect 7817 18009 7833 18043
rect 7833 18009 7851 18043
rect 7889 18009 7901 18043
rect 7901 18009 7923 18043
rect 7961 18009 7969 18043
rect 7969 18009 7995 18043
rect 8033 18009 8037 18043
rect 8037 18009 8067 18043
rect 8105 18009 8139 18043
rect 8177 18009 8207 18043
rect 8207 18009 8211 18043
rect 8249 18009 8275 18043
rect 8275 18009 8283 18043
rect 8321 18009 8343 18043
rect 8343 18009 8355 18043
rect 8393 18009 8411 18043
rect 8411 18009 8427 18043
rect 8465 18009 8479 18043
rect 8479 18009 8499 18043
rect 8537 18009 8547 18043
rect 8547 18009 8571 18043
rect 8609 18009 8615 18043
rect 8615 18009 8643 18043
rect 8681 18009 8683 18043
rect 8683 18009 8715 18043
rect 8753 18009 8785 18043
rect 8785 18009 8787 18043
rect 8825 18009 8853 18043
rect 8853 18009 8859 18043
rect 8897 18009 8921 18043
rect 8921 18009 8931 18043
rect 8969 18009 8989 18043
rect 8989 18009 9003 18043
rect 9041 18009 9057 18043
rect 9057 18009 9075 18043
rect 9113 18009 9125 18043
rect 9125 18009 9147 18043
rect 9185 18009 9193 18043
rect 9193 18009 9219 18043
rect 9257 18009 9261 18043
rect 9261 18009 9291 18043
rect 9329 18009 9363 18043
rect 9401 18009 9431 18043
rect 9431 18009 9435 18043
rect 9473 18009 9499 18043
rect 9499 18009 9507 18043
rect 9545 18009 9567 18043
rect 9567 18009 9579 18043
rect 9617 18009 9635 18043
rect 9635 18009 9651 18043
rect 9689 18009 9703 18043
rect 9703 18009 9723 18043
rect 9761 18009 9771 18043
rect 9771 18009 9795 18043
rect 9833 18009 9839 18043
rect 9839 18009 9867 18043
rect 9905 18009 9907 18043
rect 9907 18009 9939 18043
rect 9977 18009 10009 18043
rect 10009 18009 10011 18043
rect 10049 18009 10077 18043
rect 10077 18009 10083 18043
rect 10121 18009 10145 18043
rect 10145 18009 10155 18043
rect 10193 18009 10213 18043
rect 10213 18009 10227 18043
rect 10265 18009 10281 18043
rect 10281 18009 10299 18043
rect 10337 18009 10349 18043
rect 10349 18009 10371 18043
rect 10409 18009 10417 18043
rect 10417 18009 10443 18043
rect 10481 18009 10485 18043
rect 10485 18009 10515 18043
rect 10553 18009 10587 18043
rect 10625 18009 10655 18043
rect 10655 18009 10659 18043
rect 10697 18009 10723 18043
rect 10723 18009 10731 18043
rect 10769 18009 10791 18043
rect 10791 18009 10803 18043
rect 10841 18009 10859 18043
rect 10859 18009 10875 18043
rect 10913 18009 10927 18043
rect 10927 18009 10947 18043
rect 10985 18009 10995 18043
rect 10995 18009 11019 18043
rect 11057 18009 11063 18043
rect 11063 18009 11091 18043
rect 11129 18009 11131 18043
rect 11131 18009 11163 18043
rect 11201 18009 11233 18043
rect 11233 18009 11235 18043
rect 11273 18009 11301 18043
rect 11301 18009 11307 18043
rect 11345 18009 11369 18043
rect 11369 18009 11379 18043
rect 11417 18009 11437 18043
rect 11437 18009 11451 18043
rect 11489 18009 11505 18043
rect 11505 18009 11523 18043
rect 11561 18009 11573 18043
rect 11573 18009 11595 18043
rect 11633 18009 11641 18043
rect 11641 18009 11667 18043
rect 11705 18009 11709 18043
rect 11709 18009 11739 18043
rect 11777 18009 11811 18043
rect 11849 18009 11879 18043
rect 11879 18009 11883 18043
rect 11921 18009 11947 18043
rect 11947 18009 11955 18043
rect 11993 18009 12015 18043
rect 12015 18009 12027 18043
rect 12065 18009 12083 18043
rect 12083 18009 12099 18043
rect 12137 18009 12151 18043
rect 12151 18009 12171 18043
rect 12209 18009 12219 18043
rect 12219 18009 12243 18043
rect 12281 18009 12287 18043
rect 12287 18009 12315 18043
rect 12353 18009 12355 18043
rect 12355 18009 12387 18043
rect 12425 18009 12457 18043
rect 12457 18009 12459 18043
rect 12497 18009 12525 18043
rect 12525 18009 12531 18043
rect 12569 18009 12593 18043
rect 12593 18009 12603 18043
rect 12641 18009 12661 18043
rect 12661 18009 12675 18043
rect 12713 18009 12729 18043
rect 12729 18009 12747 18043
rect 12785 18009 12797 18043
rect 12797 18009 12819 18043
rect 12857 18009 12865 18043
rect 12865 18009 12891 18043
rect 12929 18009 12933 18043
rect 12933 18009 12963 18043
rect 4486 17938 4520 17972
rect 4622 17938 4656 17972
rect 4486 17865 4520 17899
rect 4622 17865 4656 17899
rect 4486 17792 4520 17826
rect 4622 17792 4656 17826
rect 4486 17719 4520 17753
rect 4622 17719 4656 17753
rect 4486 17645 4520 17679
rect 4622 17645 4656 17679
rect 4486 17571 4520 17605
rect 4622 17571 4656 17605
rect 4486 17497 4520 17531
rect 4622 17497 4656 17531
rect 4486 17423 4520 17457
rect 4622 17423 4656 17457
rect 4486 17349 4520 17383
rect 4622 17349 4656 17383
rect 4486 17275 4520 17309
rect 4622 17275 4656 17309
rect 4486 17201 4520 17235
rect 4622 17201 4656 17235
rect 4486 17127 4520 17161
rect 4622 17127 4656 17161
rect 4486 17053 4520 17087
rect 4622 17053 4656 17087
rect 4486 16979 4520 17013
rect 4622 16979 4656 17013
rect 4486 16905 4520 16939
rect 4622 16905 4656 16939
rect 4486 16831 4520 16865
rect 4622 16831 4656 16865
rect 4486 16757 4520 16791
rect 4622 16757 4656 16791
rect 4486 16683 4520 16717
rect 4622 16683 4656 16717
rect 4486 16609 4520 16643
rect 4622 16609 4656 16643
rect 4486 16535 4520 16569
rect 4622 16535 4656 16569
rect 4737 17881 4771 17915
rect 4809 17881 4843 17915
rect 4737 17807 4771 17841
rect 4809 17807 4843 17841
rect 13342 17841 13376 17875
rect 4737 17733 4771 17767
rect 4809 17733 4843 17767
rect 4737 17659 4771 17693
rect 4809 17659 4843 17693
rect 4737 17585 4771 17619
rect 4809 17585 4843 17619
rect 4737 17511 4771 17545
rect 4809 17511 4843 17545
rect 4737 17437 4771 17471
rect 4809 17437 4843 17471
rect 4737 17363 4771 17397
rect 4809 17363 4843 17397
rect 4737 17289 4771 17323
rect 4809 17289 4843 17323
rect 4737 17215 4771 17249
rect 4809 17215 4843 17249
rect 4737 17141 4771 17175
rect 4809 17141 4843 17175
rect 4737 17068 4771 17102
rect 4809 17068 4843 17102
rect 4737 16995 4771 17029
rect 4809 16995 4843 17029
rect 4737 16922 4771 16956
rect 4809 16922 4843 16956
rect 4737 16849 4771 16883
rect 4809 16849 4843 16883
rect 4737 16776 4771 16810
rect 4809 16776 4843 16810
rect 4737 16703 4771 16737
rect 4809 16703 4843 16737
rect 4737 16630 4771 16664
rect 4809 16630 4843 16664
rect 4737 16557 4771 16591
rect 4809 16557 4843 16591
rect 5062 17770 5096 17804
rect 5062 17696 5096 17730
rect 5062 17622 5096 17656
rect 5062 17548 5096 17582
rect 5062 17474 5096 17508
rect 5062 17400 5096 17434
rect 5062 17326 5096 17360
rect 5062 17252 5096 17286
rect 5062 17178 5096 17212
rect 5062 17104 5096 17138
rect 5062 17030 5096 17064
rect 5062 16956 5096 16990
rect 5062 16882 5096 16916
rect 5062 16808 5096 16842
rect 5062 16733 5096 16767
rect 5062 16658 5096 16692
rect 5062 16583 5096 16617
rect 6718 17770 6752 17804
rect 6718 17696 6752 17730
rect 6718 17622 6752 17656
rect 6718 17548 6752 17582
rect 6718 17474 6752 17508
rect 6718 17400 6752 17434
rect 6718 17326 6752 17360
rect 6718 17252 6752 17286
rect 6718 17178 6752 17212
rect 6718 17104 6752 17138
rect 6718 17030 6752 17064
rect 6718 16956 6752 16990
rect 6718 16882 6752 16916
rect 6718 16808 6752 16842
rect 6718 16733 6752 16767
rect 6718 16658 6752 16692
rect 6718 16583 6752 16617
rect 8374 17770 8408 17804
rect 8374 17696 8408 17730
rect 8374 17622 8408 17656
rect 8374 17548 8408 17582
rect 8374 17474 8408 17508
rect 8374 17400 8408 17434
rect 8374 17326 8408 17360
rect 8374 17252 8408 17286
rect 8374 17178 8408 17212
rect 8374 17104 8408 17138
rect 8374 17030 8408 17064
rect 8374 16956 8408 16990
rect 8374 16882 8408 16916
rect 8374 16808 8408 16842
rect 8374 16733 8408 16767
rect 8374 16658 8408 16692
rect 8374 16583 8408 16617
rect 10030 17770 10064 17804
rect 10030 17696 10064 17730
rect 10030 17622 10064 17656
rect 10030 17548 10064 17582
rect 10030 17474 10064 17508
rect 10030 17400 10064 17434
rect 10030 17326 10064 17360
rect 10030 17252 10064 17286
rect 10030 17178 10064 17212
rect 10030 17104 10064 17138
rect 10030 17030 10064 17064
rect 10030 16956 10064 16990
rect 10030 16882 10064 16916
rect 10030 16808 10064 16842
rect 10030 16733 10064 16767
rect 10030 16658 10064 16692
rect 10030 16583 10064 16617
rect 11686 17770 11720 17804
rect 11686 17696 11720 17730
rect 11686 17622 11720 17656
rect 11686 17548 11720 17582
rect 11686 17474 11720 17508
rect 11686 17400 11720 17434
rect 11686 17326 11720 17360
rect 11686 17252 11720 17286
rect 11686 17178 11720 17212
rect 11686 17104 11720 17138
rect 11686 17030 11720 17064
rect 11686 16956 11720 16990
rect 11686 16882 11720 16916
rect 11686 16808 11720 16842
rect 11686 16733 11720 16767
rect 11686 16658 11720 16692
rect 11686 16583 11720 16617
rect 13342 17766 13376 17800
rect 13342 17691 13376 17725
rect 13342 17616 13376 17650
rect 13342 17541 13376 17575
rect 13342 17466 13376 17500
rect 13342 17391 13376 17425
rect 13342 17316 13376 17350
rect 13342 17241 13376 17275
rect 13342 17165 13376 17199
rect 13342 17089 13376 17123
rect 13342 17013 13376 17047
rect 13342 16937 13376 16971
rect 13342 16861 13376 16895
rect 13342 16785 13376 16819
rect 13342 16709 13376 16743
rect 13342 16633 13376 16667
rect 13342 16557 13376 16591
rect 4486 16461 4520 16495
rect 4622 16466 4656 16495
rect 4622 16461 4656 16466
rect 4486 16417 4520 16421
rect 1944 15922 1946 16100
rect 1946 15922 2048 16100
rect 2048 15922 2050 16100
rect 1944 15849 1946 15883
rect 1946 15849 1978 15883
rect 2016 15849 2048 15883
rect 2048 15849 2050 15883
rect 1944 15776 1946 15810
rect 1946 15776 1978 15810
rect 2016 15776 2048 15810
rect 2048 15776 2050 15810
rect 1944 15703 1946 15737
rect 1946 15703 1978 15737
rect 2016 15703 2048 15737
rect 2048 15703 2050 15737
rect 1944 15630 1946 15664
rect 1946 15630 1978 15664
rect 2016 15630 2048 15664
rect 2048 15630 2050 15664
rect 1944 15557 1946 15591
rect 1946 15557 1978 15591
rect 2016 15557 2048 15591
rect 2048 15557 2050 15591
rect 1944 15484 1946 15518
rect 1946 15484 1978 15518
rect 2016 15484 2048 15518
rect 2048 15484 2050 15518
rect 1944 15411 1946 15445
rect 1946 15411 1978 15445
rect 2016 15411 2048 15445
rect 2048 15411 2050 15445
rect 1944 15338 1946 15372
rect 1946 15338 1978 15372
rect 2016 15338 2048 15372
rect 2048 15338 2050 15372
rect 1944 14940 1946 14974
rect 1946 14940 1978 14974
rect 2016 14940 2048 14974
rect 2048 14940 2050 14974
rect 1944 14865 1946 14899
rect 1946 14865 1978 14899
rect 2016 14865 2048 14899
rect 2048 14865 2050 14899
rect 1944 14790 1946 14824
rect 1946 14790 1978 14824
rect 2016 14790 2048 14824
rect 2048 14790 2050 14824
rect 1944 14715 1946 14749
rect 1946 14715 1978 14749
rect 2016 14715 2048 14749
rect 2048 14715 2050 14749
rect 1944 14640 1946 14674
rect 1946 14640 1978 14674
rect 2016 14640 2048 14674
rect 2048 14640 2050 14674
rect 1944 14565 1946 14599
rect 1946 14565 1978 14599
rect 2016 14565 2048 14599
rect 2048 14565 2050 14599
rect 1944 14490 1946 14524
rect 1946 14490 1978 14524
rect 2016 14490 2048 14524
rect 2048 14490 2050 14524
rect 1944 14415 1946 14449
rect 1946 14415 1978 14449
rect 2016 14415 2048 14449
rect 2048 14415 2050 14449
rect 1944 14340 1946 14374
rect 1946 14340 1978 14374
rect 2016 14340 2048 14374
rect 2048 14340 2050 14374
rect 1944 14265 1946 14299
rect 1946 14265 1978 14299
rect 2016 14265 2048 14299
rect 2048 14265 2050 14299
rect 1944 14190 1946 14224
rect 1946 14190 1978 14224
rect 2016 14190 2048 14224
rect 2048 14190 2050 14224
rect 1944 14115 1946 14149
rect 1946 14115 1978 14149
rect 2016 14115 2048 14149
rect 2048 14115 2050 14149
rect 1944 14041 1946 14075
rect 1946 14041 1978 14075
rect 2016 14041 2048 14075
rect 2048 14041 2050 14075
rect 1944 13967 1946 14001
rect 1946 13967 1978 14001
rect 2016 13967 2048 14001
rect 2048 13967 2050 14001
rect 1944 13893 1946 13927
rect 1946 13893 1978 13927
rect 2016 13893 2048 13927
rect 2048 13893 2050 13927
rect 1944 13819 1946 13853
rect 1946 13819 1978 13853
rect 2016 13819 2048 13853
rect 2048 13819 2050 13853
rect 1944 13745 1946 13779
rect 1946 13745 1978 13779
rect 2016 13745 2048 13779
rect 2048 13745 2050 13779
rect 1944 13671 1946 13705
rect 1946 13671 1978 13705
rect 2016 13671 2048 13705
rect 2048 13671 2050 13705
rect 1944 13597 1946 13631
rect 1946 13597 1978 13631
rect 2016 13597 2048 13631
rect 2048 13597 2050 13631
rect 1944 13523 1946 13557
rect 1946 13523 1978 13557
rect 2016 13523 2048 13557
rect 2048 13523 2050 13557
rect 1944 13449 1946 13483
rect 1946 13449 1978 13483
rect 2016 13449 2048 13483
rect 2048 13449 2050 13483
rect 1944 13375 1946 13409
rect 1946 13375 1978 13409
rect 2016 13375 2048 13409
rect 2048 13375 2050 13409
rect 1944 13301 1946 13335
rect 1946 13301 1978 13335
rect 2016 13301 2048 13335
rect 2048 13301 2050 13335
rect 1944 12855 1946 12889
rect 1946 12855 1978 12889
rect 2016 12855 2048 12889
rect 2048 12855 2050 12889
rect 1944 12780 1946 12814
rect 1946 12780 1978 12814
rect 2016 12780 2048 12814
rect 2048 12780 2050 12814
rect 1944 12705 1946 12739
rect 1946 12705 1978 12739
rect 2016 12705 2048 12739
rect 2048 12705 2050 12739
rect 1944 12630 1946 12664
rect 1946 12630 1978 12664
rect 2016 12630 2048 12664
rect 2048 12630 2050 12664
rect 1944 12555 1946 12589
rect 1946 12555 1978 12589
rect 2016 12555 2048 12589
rect 2048 12555 2050 12589
rect 1944 12480 1946 12514
rect 1946 12480 1978 12514
rect 2016 12480 2048 12514
rect 2048 12480 2050 12514
rect 1944 12405 1946 12439
rect 1946 12405 1978 12439
rect 2016 12405 2048 12439
rect 2048 12405 2050 12439
rect 1944 12330 1946 12364
rect 1946 12330 1978 12364
rect 2016 12330 2048 12364
rect 2048 12330 2050 12364
rect 1944 12255 1946 12289
rect 1946 12255 1978 12289
rect 2016 12255 2048 12289
rect 2048 12255 2050 12289
rect 1944 12180 1946 12214
rect 1946 12180 1978 12214
rect 2016 12180 2048 12214
rect 2048 12180 2050 12214
rect 1944 12105 1946 12139
rect 1946 12105 1978 12139
rect 2016 12105 2048 12139
rect 2048 12105 2050 12139
rect 1944 12030 1946 12064
rect 1946 12030 1978 12064
rect 2016 12030 2048 12064
rect 2048 12030 2050 12064
rect 1944 11955 1946 11989
rect 1946 11955 1978 11989
rect 2016 11955 2048 11989
rect 2048 11955 2050 11989
rect 1944 11880 1946 11914
rect 1946 11880 1978 11914
rect 2016 11880 2048 11914
rect 2048 11880 2050 11914
rect 1944 11805 1946 11839
rect 1946 11805 1978 11839
rect 2016 11805 2048 11839
rect 2048 11805 2050 11839
rect 1944 11730 1946 11764
rect 1946 11730 1978 11764
rect 2016 11730 2048 11764
rect 2048 11730 2050 11764
rect 1944 11655 1946 11689
rect 1946 11655 1978 11689
rect 2016 11655 2048 11689
rect 2048 11655 2050 11689
rect 1944 11580 1946 11614
rect 1946 11580 1978 11614
rect 2016 11580 2048 11614
rect 2048 11580 2050 11614
rect 1944 11505 1946 11539
rect 1946 11505 1978 11539
rect 2016 11505 2048 11539
rect 2048 11505 2050 11539
rect 1944 11430 1946 11464
rect 1946 11430 1978 11464
rect 2016 11430 2048 11464
rect 2048 11430 2050 11464
rect 1944 11355 1946 11389
rect 1946 11355 1978 11389
rect 2016 11355 2048 11389
rect 2048 11355 2050 11389
rect 1944 11279 1946 11313
rect 1946 11279 1978 11313
rect 2016 11279 2048 11313
rect 2048 11279 2050 11313
rect 1944 10813 1946 10847
rect 1946 10813 1978 10847
rect 2016 10813 2048 10847
rect 2048 10813 2050 10847
rect 1944 10737 1946 10771
rect 1946 10737 1978 10771
rect 2016 10737 2048 10771
rect 2048 10737 2050 10771
rect 1944 10661 1946 10695
rect 1946 10661 1978 10695
rect 2016 10661 2048 10695
rect 2048 10661 2050 10695
rect 1944 10586 1946 10620
rect 1946 10586 1978 10620
rect 2016 10586 2048 10620
rect 2048 10586 2050 10620
rect 1944 10511 1946 10545
rect 1946 10511 1978 10545
rect 2016 10511 2048 10545
rect 2048 10511 2050 10545
rect 1944 10436 1946 10470
rect 1946 10436 1978 10470
rect 2016 10436 2048 10470
rect 2048 10436 2050 10470
rect 1944 10361 1946 10395
rect 1946 10361 1978 10395
rect 2016 10361 2048 10395
rect 2048 10361 2050 10395
rect 1944 10286 1946 10320
rect 1946 10286 1978 10320
rect 2016 10286 2048 10320
rect 2048 10286 2050 10320
rect 1944 10211 1946 10245
rect 1946 10211 1978 10245
rect 2016 10211 2048 10245
rect 2048 10211 2050 10245
rect 1944 10136 1946 10170
rect 1946 10136 1978 10170
rect 2016 10136 2048 10170
rect 2048 10136 2050 10170
rect 1944 10061 1946 10095
rect 1946 10061 1978 10095
rect 2016 10061 2048 10095
rect 2048 10061 2050 10095
rect 1944 9986 1946 10020
rect 1946 9986 1978 10020
rect 2016 9986 2048 10020
rect 2048 9986 2050 10020
rect 1944 9911 1946 9945
rect 1946 9911 1978 9945
rect 2016 9911 2048 9945
rect 2048 9911 2050 9945
rect 1944 9836 1946 9870
rect 1946 9836 1978 9870
rect 2016 9836 2048 9870
rect 2048 9836 2050 9870
rect 1944 9761 1946 9795
rect 1946 9761 1978 9795
rect 2016 9761 2048 9795
rect 2048 9761 2050 9795
rect 1944 9686 1946 9720
rect 1946 9686 1978 9720
rect 2016 9686 2048 9720
rect 2048 9686 2050 9720
rect 1944 9611 1946 9645
rect 1946 9611 1978 9645
rect 2016 9611 2048 9645
rect 2048 9611 2050 9645
rect 1944 9536 1946 9570
rect 1946 9536 1978 9570
rect 2016 9536 2048 9570
rect 2048 9536 2050 9570
rect 1944 9461 1946 9495
rect 1946 9461 1978 9495
rect 2016 9461 2048 9495
rect 2048 9461 2050 9495
rect 1944 9386 1946 9420
rect 1946 9386 1978 9420
rect 2016 9386 2048 9420
rect 2048 9386 2050 9420
rect 4486 16387 4520 16417
rect 4622 16398 4656 16421
rect 4622 16387 4656 16398
rect 4923 16209 4927 16243
rect 4927 16209 4957 16243
rect 4996 16209 5029 16243
rect 5029 16209 5030 16243
rect 5069 16209 5097 16243
rect 5097 16209 5103 16243
rect 5142 16209 5165 16243
rect 5165 16209 5176 16243
rect 5215 16209 5233 16243
rect 5233 16209 5249 16243
rect 5288 16209 5301 16243
rect 5301 16209 5322 16243
rect 5361 16209 5369 16243
rect 5369 16209 5395 16243
rect 5434 16209 5437 16243
rect 5437 16209 5468 16243
rect 5507 16209 5539 16243
rect 5539 16209 5541 16243
rect 5580 16209 5607 16243
rect 5607 16209 5614 16243
rect 5653 16209 5675 16243
rect 5675 16209 5687 16243
rect 5726 16209 5743 16243
rect 5743 16209 5760 16243
rect 5799 16209 5811 16243
rect 5811 16209 5833 16243
rect 5872 16209 5879 16243
rect 5879 16209 5906 16243
rect 5945 16209 5947 16243
rect 5947 16209 5979 16243
rect 6017 16209 6049 16243
rect 6049 16209 6051 16243
rect 6089 16209 6117 16243
rect 6117 16209 6123 16243
rect 6161 16209 6185 16243
rect 6185 16209 6195 16243
rect 6233 16209 6253 16243
rect 6253 16209 6267 16243
rect 6305 16209 6321 16243
rect 6321 16209 6339 16243
rect 6377 16209 6389 16243
rect 6389 16209 6411 16243
rect 6449 16209 6457 16243
rect 6457 16209 6483 16243
rect 6521 16209 6525 16243
rect 6525 16209 6555 16243
rect 6593 16209 6627 16243
rect 6665 16209 6695 16243
rect 6695 16209 6699 16243
rect 6737 16209 6763 16243
rect 6763 16209 6771 16243
rect 6809 16209 6831 16243
rect 6831 16209 6843 16243
rect 6881 16209 6899 16243
rect 6899 16209 6915 16243
rect 6953 16209 6967 16243
rect 6967 16209 6987 16243
rect 7025 16209 7035 16243
rect 7035 16209 7059 16243
rect 7097 16209 7103 16243
rect 7103 16209 7131 16243
rect 7169 16209 7171 16243
rect 7171 16209 7203 16243
rect 7241 16209 7273 16243
rect 7273 16209 7275 16243
rect 7313 16209 7341 16243
rect 7341 16209 7347 16243
rect 7385 16209 7409 16243
rect 7409 16209 7419 16243
rect 7457 16209 7477 16243
rect 7477 16209 7491 16243
rect 7529 16209 7545 16243
rect 7545 16209 7563 16243
rect 7601 16209 7613 16243
rect 7613 16209 7635 16243
rect 7673 16209 7681 16243
rect 7681 16209 7707 16243
rect 7745 16209 7749 16243
rect 7749 16209 7779 16243
rect 7817 16209 7851 16243
rect 7889 16209 7919 16243
rect 7919 16209 7923 16243
rect 7961 16209 7987 16243
rect 7987 16209 7995 16243
rect 8033 16209 8055 16243
rect 8055 16209 8067 16243
rect 8105 16209 8123 16243
rect 8123 16209 8139 16243
rect 8177 16209 8191 16243
rect 8191 16209 8211 16243
rect 8249 16209 8259 16243
rect 8259 16209 8283 16243
rect 8321 16209 8327 16243
rect 8327 16209 8355 16243
rect 8393 16209 8395 16243
rect 8395 16209 8427 16243
rect 8465 16209 8497 16243
rect 8497 16209 8499 16243
rect 8537 16209 8565 16243
rect 8565 16209 8571 16243
rect 8609 16209 8633 16243
rect 8633 16209 8643 16243
rect 8681 16209 8701 16243
rect 8701 16209 8715 16243
rect 8753 16209 8769 16243
rect 8769 16209 8787 16243
rect 8825 16209 8837 16243
rect 8837 16209 8859 16243
rect 8897 16209 8905 16243
rect 8905 16209 8931 16243
rect 8969 16209 8973 16243
rect 8973 16209 9003 16243
rect 9041 16209 9075 16243
rect 9113 16209 9143 16243
rect 9143 16209 9147 16243
rect 9185 16209 9211 16243
rect 9211 16209 9219 16243
rect 9257 16209 9279 16243
rect 9279 16209 9291 16243
rect 9329 16209 9347 16243
rect 9347 16209 9363 16243
rect 9401 16209 9415 16243
rect 9415 16209 9435 16243
rect 9473 16209 9483 16243
rect 9483 16209 9507 16243
rect 9545 16209 9551 16243
rect 9551 16209 9579 16243
rect 9617 16209 9619 16243
rect 9619 16209 9651 16243
rect 9689 16209 9721 16243
rect 9721 16209 9723 16243
rect 9761 16209 9789 16243
rect 9789 16209 9795 16243
rect 9833 16209 9857 16243
rect 9857 16209 9867 16243
rect 9905 16209 9925 16243
rect 9925 16209 9939 16243
rect 9977 16209 9993 16243
rect 9993 16209 10011 16243
rect 10049 16209 10061 16243
rect 10061 16209 10083 16243
rect 10121 16209 10129 16243
rect 10129 16209 10155 16243
rect 10193 16209 10197 16243
rect 10197 16209 10227 16243
rect 10265 16209 10299 16243
rect 10337 16209 10367 16243
rect 10367 16209 10371 16243
rect 10409 16209 10435 16243
rect 10435 16209 10443 16243
rect 10481 16209 10503 16243
rect 10503 16209 10515 16243
rect 10553 16209 10571 16243
rect 10571 16209 10587 16243
rect 10625 16209 10639 16243
rect 10639 16209 10659 16243
rect 10697 16209 10707 16243
rect 10707 16209 10731 16243
rect 10769 16209 10775 16243
rect 10775 16209 10803 16243
rect 10841 16209 10843 16243
rect 10843 16209 10875 16243
rect 10913 16209 10945 16243
rect 10945 16209 10947 16243
rect 10985 16209 11013 16243
rect 11013 16209 11019 16243
rect 11057 16209 11081 16243
rect 11081 16209 11091 16243
rect 11129 16209 11149 16243
rect 11149 16209 11163 16243
rect 11201 16209 11217 16243
rect 11217 16209 11235 16243
rect 11273 16209 11285 16243
rect 11285 16209 11307 16243
rect 11345 16209 11353 16243
rect 11353 16209 11379 16243
rect 11417 16209 11421 16243
rect 11421 16209 11451 16243
rect 11489 16209 11523 16243
rect 11561 16209 11591 16243
rect 11591 16209 11595 16243
rect 11633 16209 11659 16243
rect 11659 16209 11667 16243
rect 11705 16209 11727 16243
rect 11727 16209 11739 16243
rect 11777 16209 11795 16243
rect 11795 16209 11811 16243
rect 11849 16209 11863 16243
rect 11863 16209 11883 16243
rect 11921 16209 11931 16243
rect 11931 16209 11955 16243
rect 11993 16209 11999 16243
rect 11999 16209 12027 16243
rect 12065 16209 12067 16243
rect 12067 16209 12099 16243
rect 12137 16209 12169 16243
rect 12169 16209 12171 16243
rect 12209 16209 12237 16243
rect 12237 16209 12243 16243
rect 12281 16209 12305 16243
rect 12305 16209 12315 16243
rect 12353 16209 12373 16243
rect 12373 16209 12387 16243
rect 12425 16209 12441 16243
rect 12441 16209 12459 16243
rect 12497 16209 12509 16243
rect 12509 16209 12531 16243
rect 12569 16209 12577 16243
rect 12577 16209 12603 16243
rect 12641 16209 12645 16243
rect 12645 16209 12675 16243
rect 12713 16209 12747 16243
rect 12785 16209 12815 16243
rect 12815 16209 12819 16243
rect 12857 16209 12883 16243
rect 12883 16209 12891 16243
rect 12929 16209 12951 16243
rect 12951 16209 12963 16243
rect 13342 16073 13376 16107
rect 2280 16006 2314 16040
rect 2404 16006 2438 16040
rect 2280 15931 2314 15965
rect 2404 15931 2438 15965
rect 2280 15856 2314 15890
rect 2404 15856 2438 15890
rect 2280 15781 2314 15815
rect 2404 15781 2438 15815
rect 2280 15706 2314 15740
rect 2404 15706 2438 15740
rect 2280 15631 2314 15665
rect 2404 15631 2438 15665
rect 2280 15555 2314 15589
rect 2404 15555 2438 15589
rect 2280 15479 2314 15513
rect 2404 15479 2438 15513
rect 2280 15403 2314 15437
rect 2404 15403 2438 15437
rect 2280 15327 2314 15361
rect 2404 15327 2438 15361
rect 2280 15251 2314 15285
rect 2404 15251 2438 15285
rect 2280 15175 2314 15209
rect 2404 15175 2438 15209
rect 2550 16026 2584 16060
rect 2550 15953 2584 15987
rect 2550 15880 2584 15914
rect 2550 15807 2584 15841
rect 2550 15734 2584 15768
rect 2550 15661 2584 15695
rect 2550 15589 2584 15623
rect 2550 15517 2584 15551
rect 2550 15445 2584 15479
rect 2550 15373 2584 15407
rect 2550 15301 2584 15335
rect 2550 15229 2584 15263
rect 2550 15157 2584 15191
rect 3406 16026 3440 16060
rect 3406 15953 3440 15987
rect 3406 15880 3440 15914
rect 3406 15807 3440 15841
rect 3406 15734 3440 15768
rect 3406 15661 3440 15695
rect 3406 15589 3440 15623
rect 3406 15517 3440 15551
rect 3406 15445 3440 15479
rect 3406 15373 3440 15407
rect 3406 15301 3440 15335
rect 3406 15229 3440 15263
rect 3406 15157 3440 15191
rect 5062 16026 5096 16060
rect 5062 15953 5096 15987
rect 5062 15880 5096 15914
rect 5062 15807 5096 15841
rect 5062 15734 5096 15768
rect 5062 15661 5096 15695
rect 5062 15589 5096 15623
rect 5062 15517 5096 15551
rect 5062 15445 5096 15479
rect 5062 15373 5096 15407
rect 5062 15301 5096 15335
rect 5062 15229 5096 15263
rect 5062 15157 5096 15191
rect 6718 16026 6752 16060
rect 6718 15953 6752 15987
rect 6718 15880 6752 15914
rect 6718 15807 6752 15841
rect 6718 15734 6752 15768
rect 6718 15661 6752 15695
rect 6718 15589 6752 15623
rect 6718 15517 6752 15551
rect 6718 15445 6752 15479
rect 6718 15373 6752 15407
rect 6718 15301 6752 15335
rect 6718 15229 6752 15263
rect 6718 15157 6752 15191
rect 8374 16026 8408 16060
rect 8374 15953 8408 15987
rect 8374 15880 8408 15914
rect 8374 15807 8408 15841
rect 8374 15734 8408 15768
rect 8374 15661 8408 15695
rect 8374 15589 8408 15623
rect 8374 15517 8408 15551
rect 8374 15445 8408 15479
rect 8374 15373 8408 15407
rect 8374 15301 8408 15335
rect 8374 15229 8408 15263
rect 8374 15157 8408 15191
rect 10030 16026 10064 16060
rect 10030 15953 10064 15987
rect 10030 15880 10064 15914
rect 10030 15807 10064 15841
rect 10030 15734 10064 15768
rect 10030 15661 10064 15695
rect 10030 15589 10064 15623
rect 10030 15517 10064 15551
rect 10030 15445 10064 15479
rect 10030 15373 10064 15407
rect 10030 15301 10064 15335
rect 10030 15229 10064 15263
rect 10030 15157 10064 15191
rect 11686 16026 11720 16060
rect 11686 15953 11720 15987
rect 11686 15880 11720 15914
rect 11686 15807 11720 15841
rect 11686 15734 11720 15768
rect 11686 15661 11720 15695
rect 11686 15589 11720 15623
rect 11686 15517 11720 15551
rect 11686 15445 11720 15479
rect 11686 15373 11720 15407
rect 11686 15301 11720 15335
rect 11686 15229 11720 15263
rect 11686 15157 11720 15191
rect 13342 15996 13376 16030
rect 13342 15919 13376 15953
rect 13342 15842 13376 15876
rect 13342 15765 13376 15799
rect 13342 15689 13376 15723
rect 13342 15613 13376 15647
rect 13342 15537 13376 15571
rect 13342 15461 13376 15495
rect 13342 15385 13376 15419
rect 13342 15309 13376 15343
rect 13342 15233 13376 15267
rect 13342 15157 13376 15191
rect 2280 14953 2314 14987
rect 2404 14953 2438 14987
rect 2280 14878 2314 14912
rect 2404 14878 2438 14912
rect 2280 14803 2314 14837
rect 2404 14803 2438 14837
rect 2280 14728 2314 14762
rect 2404 14728 2438 14762
rect 2280 14653 2314 14687
rect 2404 14653 2438 14687
rect 2280 14578 2314 14612
rect 2404 14578 2438 14612
rect 2280 14503 2314 14537
rect 2404 14503 2438 14537
rect 2280 14428 2314 14462
rect 2404 14428 2438 14462
rect 2280 14353 2314 14387
rect 2404 14353 2438 14387
rect 2280 14278 2314 14312
rect 2404 14278 2438 14312
rect 2280 14203 2314 14237
rect 2404 14203 2438 14237
rect 2280 14128 2314 14162
rect 2404 14128 2438 14162
rect 2280 14053 2314 14087
rect 2404 14053 2438 14087
rect 2280 13978 2314 14012
rect 2404 13978 2438 14012
rect 2280 13903 2314 13937
rect 2404 13903 2438 13937
rect 2280 13828 2314 13862
rect 2404 13828 2438 13862
rect 2280 13753 2314 13787
rect 2404 13753 2438 13787
rect 2280 13678 2314 13712
rect 2404 13678 2438 13712
rect 2280 13602 2314 13636
rect 2404 13602 2438 13636
rect 2280 13526 2314 13560
rect 2404 13526 2438 13560
rect 2280 13450 2314 13484
rect 2404 13450 2438 13484
rect 2280 13374 2314 13408
rect 2404 13374 2438 13408
rect 2679 14311 2713 14345
rect 2751 14311 2785 14345
rect 2679 14233 2713 14267
rect 2751 14233 2785 14267
rect 2679 14155 2713 14189
rect 2751 14155 2785 14189
rect 2679 14077 2713 14111
rect 2751 14077 2785 14111
rect 2679 13999 2713 14033
rect 2751 13999 2785 14033
rect 2679 13921 2713 13955
rect 2751 13921 2785 13955
rect 2679 13843 2713 13877
rect 2751 13843 2785 13877
rect 2679 13765 2713 13799
rect 2751 13765 2785 13799
rect 2679 13688 2713 13722
rect 2751 13688 2785 13722
rect 2679 13611 2713 13645
rect 2751 13611 2785 13645
rect 2679 13534 2713 13568
rect 2751 13534 2785 13568
rect 2679 13457 2713 13491
rect 2751 13457 2785 13491
rect 2679 13380 2713 13414
rect 2751 13380 2785 13414
rect 2956 14311 2990 14345
rect 3028 14311 3062 14345
rect 2956 14233 2990 14267
rect 3028 14233 3062 14267
rect 2956 14155 2990 14189
rect 3028 14155 3062 14189
rect 2956 14077 2990 14111
rect 3028 14077 3062 14111
rect 2956 13999 2990 14033
rect 3028 13999 3062 14033
rect 2956 13921 2990 13955
rect 3028 13921 3062 13955
rect 2956 13843 2990 13877
rect 3028 13843 3062 13877
rect 2956 13765 2990 13799
rect 3028 13765 3062 13799
rect 2956 13688 2990 13722
rect 3028 13688 3062 13722
rect 2956 13611 2990 13645
rect 3028 13611 3062 13645
rect 2956 13534 2990 13568
rect 3028 13534 3062 13568
rect 2956 13457 2990 13491
rect 3028 13457 3062 13491
rect 2956 13380 2990 13414
rect 3028 13380 3062 13414
rect 3233 14311 3267 14345
rect 3305 14311 3339 14345
rect 3233 14233 3267 14267
rect 3305 14233 3339 14267
rect 3233 14155 3267 14189
rect 3305 14155 3339 14189
rect 3233 14077 3267 14111
rect 3305 14077 3339 14111
rect 3233 13999 3267 14033
rect 3305 13999 3339 14033
rect 3233 13921 3267 13955
rect 3305 13921 3339 13955
rect 3233 13843 3267 13877
rect 3305 13843 3339 13877
rect 3233 13765 3267 13799
rect 3305 13765 3339 13799
rect 3233 13688 3267 13722
rect 3305 13688 3339 13722
rect 3233 13611 3267 13645
rect 3305 13611 3339 13645
rect 3233 13534 3267 13568
rect 3305 13534 3339 13568
rect 3233 13457 3267 13491
rect 3305 13457 3339 13491
rect 3233 13380 3267 13414
rect 3305 13380 3339 13414
rect 3510 14311 3544 14345
rect 3582 14311 3616 14345
rect 3510 14233 3544 14267
rect 3582 14233 3616 14267
rect 3510 14155 3544 14189
rect 3582 14155 3616 14189
rect 3510 14077 3544 14111
rect 3582 14077 3616 14111
rect 3510 13999 3544 14033
rect 3582 13999 3616 14033
rect 3510 13921 3544 13955
rect 3582 13921 3616 13955
rect 3510 13843 3544 13877
rect 3582 13843 3616 13877
rect 3510 13765 3544 13799
rect 3582 13765 3616 13799
rect 3510 13688 3544 13722
rect 3582 13688 3616 13722
rect 3510 13611 3544 13645
rect 3582 13611 3616 13645
rect 3510 13534 3544 13568
rect 3582 13534 3616 13568
rect 3510 13457 3544 13491
rect 3582 13457 3616 13491
rect 3510 13380 3544 13414
rect 3582 13380 3616 13414
rect 3787 14311 3821 14345
rect 3859 14311 3893 14345
rect 3787 14233 3821 14267
rect 3859 14233 3893 14267
rect 3787 14155 3821 14189
rect 3859 14155 3893 14189
rect 3787 14077 3821 14111
rect 3859 14077 3893 14111
rect 3787 13999 3821 14033
rect 3859 13999 3893 14033
rect 3787 13921 3821 13955
rect 3859 13921 3893 13955
rect 3787 13843 3821 13877
rect 3859 13843 3893 13877
rect 3787 13765 3821 13799
rect 3859 13765 3893 13799
rect 3787 13688 3821 13722
rect 3859 13688 3893 13722
rect 3787 13611 3821 13645
rect 3859 13611 3893 13645
rect 3787 13534 3821 13568
rect 3859 13534 3893 13568
rect 3787 13457 3821 13491
rect 3859 13457 3893 13491
rect 3787 13380 3821 13414
rect 3859 13380 3893 13414
rect 4064 14311 4098 14345
rect 4136 14311 4170 14345
rect 4064 14233 4098 14267
rect 4136 14233 4170 14267
rect 4064 14155 4098 14189
rect 4136 14155 4170 14189
rect 4064 14077 4098 14111
rect 4136 14077 4170 14111
rect 4064 13999 4098 14033
rect 4136 13999 4170 14033
rect 4064 13921 4098 13955
rect 4136 13921 4170 13955
rect 4064 13843 4098 13877
rect 4136 13843 4170 13877
rect 4064 13765 4098 13799
rect 4136 13765 4170 13799
rect 4064 13688 4098 13722
rect 4136 13688 4170 13722
rect 4064 13611 4098 13645
rect 4136 13611 4170 13645
rect 4064 13534 4098 13568
rect 4136 13534 4170 13568
rect 4064 13457 4098 13491
rect 4136 13457 4170 13491
rect 4064 13380 4098 13414
rect 4136 13380 4170 13414
rect 4341 14311 4375 14345
rect 4413 14311 4447 14345
rect 4341 14233 4375 14267
rect 4413 14233 4447 14267
rect 4341 14155 4375 14189
rect 4413 14155 4447 14189
rect 4341 14077 4375 14111
rect 4413 14077 4447 14111
rect 4341 13999 4375 14033
rect 4413 13999 4447 14033
rect 4341 13921 4375 13955
rect 4413 13921 4447 13955
rect 4341 13843 4375 13877
rect 4413 13843 4447 13877
rect 4341 13765 4375 13799
rect 4413 13765 4447 13799
rect 4341 13688 4375 13722
rect 4413 13688 4447 13722
rect 4341 13611 4375 13645
rect 4413 13611 4447 13645
rect 4341 13534 4375 13568
rect 4413 13534 4447 13568
rect 4341 13457 4375 13491
rect 4413 13457 4447 13491
rect 4341 13380 4375 13414
rect 4413 13380 4447 13414
rect 4618 14311 4652 14345
rect 4690 14311 4724 14345
rect 4618 14233 4652 14267
rect 4690 14233 4724 14267
rect 4618 14155 4652 14189
rect 4690 14155 4724 14189
rect 4618 14077 4652 14111
rect 4690 14077 4724 14111
rect 4618 13999 4652 14033
rect 4690 13999 4724 14033
rect 4618 13921 4652 13955
rect 4690 13921 4724 13955
rect 4618 13843 4652 13877
rect 4690 13843 4724 13877
rect 4618 13765 4652 13799
rect 4690 13765 4724 13799
rect 4618 13688 4652 13722
rect 4690 13688 4724 13722
rect 4618 13611 4652 13645
rect 4690 13611 4724 13645
rect 4618 13534 4652 13568
rect 4690 13534 4724 13568
rect 4618 13457 4652 13491
rect 4690 13457 4724 13491
rect 4618 13380 4652 13414
rect 4690 13380 4724 13414
rect 4895 14311 4929 14345
rect 4967 14311 5001 14345
rect 4895 14233 4929 14267
rect 4967 14233 5001 14267
rect 4895 14155 4929 14189
rect 4967 14155 5001 14189
rect 4895 14077 4929 14111
rect 4967 14077 5001 14111
rect 4895 13999 4929 14033
rect 4967 13999 5001 14033
rect 4895 13921 4929 13955
rect 4967 13921 5001 13955
rect 4895 13843 4929 13877
rect 4967 13843 5001 13877
rect 4895 13765 4929 13799
rect 4967 13765 5001 13799
rect 4895 13688 4929 13722
rect 4967 13688 5001 13722
rect 4895 13611 4929 13645
rect 4967 13611 5001 13645
rect 4895 13534 4929 13568
rect 4967 13534 5001 13568
rect 4895 13457 4929 13491
rect 4967 13457 5001 13491
rect 4895 13380 4929 13414
rect 4967 13380 5001 13414
rect 5172 14311 5206 14345
rect 5244 14311 5278 14345
rect 5172 14233 5206 14267
rect 5244 14233 5278 14267
rect 5172 14155 5206 14189
rect 5244 14155 5278 14189
rect 5172 14077 5206 14111
rect 5244 14077 5278 14111
rect 5172 13999 5206 14033
rect 5244 13999 5278 14033
rect 5172 13921 5206 13955
rect 5244 13921 5278 13955
rect 5172 13843 5206 13877
rect 5244 13843 5278 13877
rect 5172 13765 5206 13799
rect 5244 13765 5278 13799
rect 5172 13688 5206 13722
rect 5244 13688 5278 13722
rect 5172 13611 5206 13645
rect 5244 13611 5278 13645
rect 5172 13534 5206 13568
rect 5244 13534 5278 13568
rect 5172 13457 5206 13491
rect 5244 13457 5278 13491
rect 5172 13380 5206 13414
rect 5244 13380 5278 13414
rect 5449 14311 5483 14345
rect 5521 14311 5555 14345
rect 5449 14233 5483 14267
rect 5521 14233 5555 14267
rect 5449 14155 5483 14189
rect 5521 14155 5555 14189
rect 5449 14077 5483 14111
rect 5521 14077 5555 14111
rect 5449 13999 5483 14033
rect 5521 13999 5555 14033
rect 5449 13921 5483 13955
rect 5521 13921 5555 13955
rect 5449 13843 5483 13877
rect 5521 13843 5555 13877
rect 5449 13765 5483 13799
rect 5521 13765 5555 13799
rect 5449 13688 5483 13722
rect 5521 13688 5555 13722
rect 5449 13611 5483 13645
rect 5521 13611 5555 13645
rect 5449 13534 5483 13568
rect 5521 13534 5555 13568
rect 5449 13457 5483 13491
rect 5521 13457 5555 13491
rect 5449 13380 5483 13414
rect 5521 13380 5555 13414
rect 5726 14311 5760 14345
rect 5798 14311 5832 14345
rect 5726 14233 5760 14267
rect 5798 14233 5832 14267
rect 5726 14155 5760 14189
rect 5798 14155 5832 14189
rect 5726 14077 5760 14111
rect 5798 14077 5832 14111
rect 5726 13999 5760 14033
rect 5798 13999 5832 14033
rect 5726 13921 5760 13955
rect 5798 13921 5832 13955
rect 5726 13843 5760 13877
rect 5798 13843 5832 13877
rect 5726 13765 5760 13799
rect 5798 13765 5832 13799
rect 5726 13688 5760 13722
rect 5798 13688 5832 13722
rect 5726 13611 5760 13645
rect 5798 13611 5832 13645
rect 5726 13534 5760 13568
rect 5798 13534 5832 13568
rect 5726 13457 5760 13491
rect 5798 13457 5832 13491
rect 5726 13380 5760 13414
rect 5798 13380 5832 13414
rect 6003 14311 6037 14345
rect 6075 14311 6109 14345
rect 6003 14233 6037 14267
rect 6075 14233 6109 14267
rect 6003 14155 6037 14189
rect 6075 14155 6109 14189
rect 6003 14077 6037 14111
rect 6075 14077 6109 14111
rect 6003 13999 6037 14033
rect 6075 13999 6109 14033
rect 6003 13921 6037 13955
rect 6075 13921 6109 13955
rect 6003 13843 6037 13877
rect 6075 13843 6109 13877
rect 6003 13765 6037 13799
rect 6075 13765 6109 13799
rect 6003 13688 6037 13722
rect 6075 13688 6109 13722
rect 6003 13611 6037 13645
rect 6075 13611 6109 13645
rect 6003 13534 6037 13568
rect 6075 13534 6109 13568
rect 6003 13457 6037 13491
rect 6075 13457 6109 13491
rect 6003 13380 6037 13414
rect 6075 13380 6109 13414
rect 6280 14311 6314 14345
rect 6352 14311 6386 14345
rect 6280 14233 6314 14267
rect 6352 14233 6386 14267
rect 6280 14155 6314 14189
rect 6352 14155 6386 14189
rect 6280 14077 6314 14111
rect 6352 14077 6386 14111
rect 6280 13999 6314 14033
rect 6352 13999 6386 14033
rect 6280 13921 6314 13955
rect 6352 13921 6386 13955
rect 6280 13843 6314 13877
rect 6352 13843 6386 13877
rect 6280 13765 6314 13799
rect 6352 13765 6386 13799
rect 6280 13688 6314 13722
rect 6352 13688 6386 13722
rect 6280 13611 6314 13645
rect 6352 13611 6386 13645
rect 6280 13534 6314 13568
rect 6352 13534 6386 13568
rect 6280 13457 6314 13491
rect 6352 13457 6386 13491
rect 6280 13380 6314 13414
rect 6352 13380 6386 13414
rect 6557 14311 6591 14345
rect 6629 14311 6663 14345
rect 6557 14233 6591 14267
rect 6629 14233 6663 14267
rect 6557 14155 6591 14189
rect 6629 14155 6663 14189
rect 6557 14077 6591 14111
rect 6629 14077 6663 14111
rect 6557 13999 6591 14033
rect 6629 13999 6663 14033
rect 6557 13921 6591 13955
rect 6629 13921 6663 13955
rect 6557 13843 6591 13877
rect 6629 13843 6663 13877
rect 6557 13765 6591 13799
rect 6629 13765 6663 13799
rect 6557 13688 6591 13722
rect 6629 13688 6663 13722
rect 6557 13611 6591 13645
rect 6629 13611 6663 13645
rect 6557 13534 6591 13568
rect 6629 13534 6663 13568
rect 6557 13457 6591 13491
rect 6629 13457 6663 13491
rect 6557 13380 6591 13414
rect 6629 13380 6663 13414
rect 6834 14311 6868 14345
rect 6906 14311 6940 14345
rect 6834 14233 6868 14267
rect 6906 14233 6940 14267
rect 6834 14155 6868 14189
rect 6906 14155 6940 14189
rect 6834 14077 6868 14111
rect 6906 14077 6940 14111
rect 6834 13999 6868 14033
rect 6906 13999 6940 14033
rect 6834 13921 6868 13955
rect 6906 13921 6940 13955
rect 6834 13843 6868 13877
rect 6906 13843 6940 13877
rect 6834 13765 6868 13799
rect 6906 13765 6940 13799
rect 6834 13688 6868 13722
rect 6906 13688 6940 13722
rect 6834 13611 6868 13645
rect 6906 13611 6940 13645
rect 6834 13534 6868 13568
rect 6906 13534 6940 13568
rect 6834 13457 6868 13491
rect 6906 13457 6940 13491
rect 6834 13380 6868 13414
rect 6906 13380 6940 13414
rect 7111 14311 7145 14345
rect 7183 14311 7217 14345
rect 7111 14233 7145 14267
rect 7183 14233 7217 14267
rect 7111 14155 7145 14189
rect 7183 14155 7217 14189
rect 7111 14077 7145 14111
rect 7183 14077 7217 14111
rect 7111 13999 7145 14033
rect 7183 13999 7217 14033
rect 7111 13921 7145 13955
rect 7183 13921 7217 13955
rect 7111 13843 7145 13877
rect 7183 13843 7217 13877
rect 7111 13765 7145 13799
rect 7183 13765 7217 13799
rect 7111 13688 7145 13722
rect 7183 13688 7217 13722
rect 7111 13611 7145 13645
rect 7183 13611 7217 13645
rect 7111 13534 7145 13568
rect 7183 13534 7217 13568
rect 7111 13457 7145 13491
rect 7183 13457 7217 13491
rect 7111 13380 7145 13414
rect 7183 13380 7217 13414
rect 7388 14311 7422 14345
rect 7460 14311 7494 14345
rect 7388 14233 7422 14267
rect 7460 14233 7494 14267
rect 7388 14155 7422 14189
rect 7460 14155 7494 14189
rect 7388 14077 7422 14111
rect 7460 14077 7494 14111
rect 7388 13999 7422 14033
rect 7460 13999 7494 14033
rect 7388 13921 7422 13955
rect 7460 13921 7494 13955
rect 7388 13843 7422 13877
rect 7460 13843 7494 13877
rect 7388 13765 7422 13799
rect 7460 13765 7494 13799
rect 7388 13688 7422 13722
rect 7460 13688 7494 13722
rect 7388 13611 7422 13645
rect 7460 13611 7494 13645
rect 7388 13534 7422 13568
rect 7460 13534 7494 13568
rect 7388 13457 7422 13491
rect 7460 13457 7494 13491
rect 7388 13380 7422 13414
rect 7460 13380 7494 13414
rect 7665 14311 7699 14345
rect 7737 14311 7771 14345
rect 7665 14233 7699 14267
rect 7737 14233 7771 14267
rect 7665 14155 7699 14189
rect 7737 14155 7771 14189
rect 7665 14077 7699 14111
rect 7737 14077 7771 14111
rect 7665 13999 7699 14033
rect 7737 13999 7771 14033
rect 7665 13921 7699 13955
rect 7737 13921 7771 13955
rect 7665 13843 7699 13877
rect 7737 13843 7771 13877
rect 7665 13765 7699 13799
rect 7737 13765 7771 13799
rect 7665 13688 7699 13722
rect 7737 13688 7771 13722
rect 7665 13611 7699 13645
rect 7737 13611 7771 13645
rect 7665 13534 7699 13568
rect 7737 13534 7771 13568
rect 7665 13457 7699 13491
rect 7737 13457 7771 13491
rect 7665 13380 7699 13414
rect 7737 13380 7771 13414
rect 7942 14311 7976 14345
rect 8014 14311 8048 14345
rect 7942 14233 7976 14267
rect 8014 14233 8048 14267
rect 7942 14155 7976 14189
rect 8014 14155 8048 14189
rect 7942 14077 7976 14111
rect 8014 14077 8048 14111
rect 7942 13999 7976 14033
rect 8014 13999 8048 14033
rect 7942 13921 7976 13955
rect 8014 13921 8048 13955
rect 7942 13843 7976 13877
rect 8014 13843 8048 13877
rect 7942 13765 7976 13799
rect 8014 13765 8048 13799
rect 7942 13688 7976 13722
rect 8014 13688 8048 13722
rect 7942 13611 7976 13645
rect 8014 13611 8048 13645
rect 7942 13534 7976 13568
rect 8014 13534 8048 13568
rect 7942 13457 7976 13491
rect 8014 13457 8048 13491
rect 7942 13380 7976 13414
rect 8014 13380 8048 13414
rect 8219 14311 8253 14345
rect 8291 14311 8325 14345
rect 8219 14233 8253 14267
rect 8291 14233 8325 14267
rect 8219 14155 8253 14189
rect 8291 14155 8325 14189
rect 8219 14077 8253 14111
rect 8291 14077 8325 14111
rect 8219 13999 8253 14033
rect 8291 13999 8325 14033
rect 8219 13921 8253 13955
rect 8291 13921 8325 13955
rect 8219 13843 8253 13877
rect 8291 13843 8325 13877
rect 8219 13765 8253 13799
rect 8291 13765 8325 13799
rect 8219 13688 8253 13722
rect 8291 13688 8325 13722
rect 8219 13611 8253 13645
rect 8291 13611 8325 13645
rect 8219 13534 8253 13568
rect 8291 13534 8325 13568
rect 8219 13457 8253 13491
rect 8291 13457 8325 13491
rect 8219 13380 8253 13414
rect 8291 13380 8325 13414
rect 8496 14311 8530 14345
rect 8568 14311 8602 14345
rect 8496 14233 8530 14267
rect 8568 14233 8602 14267
rect 8496 14155 8530 14189
rect 8568 14155 8602 14189
rect 8496 14077 8530 14111
rect 8568 14077 8602 14111
rect 8496 13999 8530 14033
rect 8568 13999 8602 14033
rect 8496 13921 8530 13955
rect 8568 13921 8602 13955
rect 8496 13843 8530 13877
rect 8568 13843 8602 13877
rect 8496 13765 8530 13799
rect 8568 13765 8602 13799
rect 8496 13688 8530 13722
rect 8568 13688 8602 13722
rect 8496 13611 8530 13645
rect 8568 13611 8602 13645
rect 8496 13534 8530 13568
rect 8568 13534 8602 13568
rect 8496 13457 8530 13491
rect 8568 13457 8602 13491
rect 8496 13380 8530 13414
rect 8568 13380 8602 13414
rect 8773 14311 8807 14345
rect 8845 14311 8879 14345
rect 8773 14233 8807 14267
rect 8845 14233 8879 14267
rect 8773 14155 8807 14189
rect 8845 14155 8879 14189
rect 8773 14077 8807 14111
rect 8845 14077 8879 14111
rect 8773 13999 8807 14033
rect 8845 13999 8879 14033
rect 8773 13921 8807 13955
rect 8845 13921 8879 13955
rect 8773 13843 8807 13877
rect 8845 13843 8879 13877
rect 8773 13765 8807 13799
rect 8845 13765 8879 13799
rect 8773 13688 8807 13722
rect 8845 13688 8879 13722
rect 8773 13611 8807 13645
rect 8845 13611 8879 13645
rect 8773 13534 8807 13568
rect 8845 13534 8879 13568
rect 8773 13457 8807 13491
rect 8845 13457 8879 13491
rect 8773 13380 8807 13414
rect 8845 13380 8879 13414
rect 9050 14311 9084 14345
rect 9122 14311 9156 14345
rect 9050 14233 9084 14267
rect 9122 14233 9156 14267
rect 9050 14155 9084 14189
rect 9122 14155 9156 14189
rect 9050 14077 9084 14111
rect 9122 14077 9156 14111
rect 9050 13999 9084 14033
rect 9122 13999 9156 14033
rect 9050 13921 9084 13955
rect 9122 13921 9156 13955
rect 9050 13843 9084 13877
rect 9122 13843 9156 13877
rect 9050 13765 9084 13799
rect 9122 13765 9156 13799
rect 9050 13688 9084 13722
rect 9122 13688 9156 13722
rect 9050 13611 9084 13645
rect 9122 13611 9156 13645
rect 9050 13534 9084 13568
rect 9122 13534 9156 13568
rect 9050 13457 9084 13491
rect 9122 13457 9156 13491
rect 9050 13380 9084 13414
rect 9122 13380 9156 13414
rect 9327 14311 9361 14345
rect 9399 14311 9433 14345
rect 9327 14233 9361 14267
rect 9399 14233 9433 14267
rect 9327 14155 9361 14189
rect 9399 14155 9433 14189
rect 9327 14077 9361 14111
rect 9399 14077 9433 14111
rect 9327 13999 9361 14033
rect 9399 13999 9433 14033
rect 9327 13921 9361 13955
rect 9399 13921 9433 13955
rect 9327 13843 9361 13877
rect 9399 13843 9433 13877
rect 9327 13765 9361 13799
rect 9399 13765 9433 13799
rect 9327 13688 9361 13722
rect 9399 13688 9433 13722
rect 9327 13611 9361 13645
rect 9399 13611 9433 13645
rect 9327 13534 9361 13568
rect 9399 13534 9433 13568
rect 9327 13457 9361 13491
rect 9399 13457 9433 13491
rect 9327 13380 9361 13414
rect 9399 13380 9433 13414
rect 9604 14311 9638 14345
rect 9676 14311 9710 14345
rect 9604 14233 9638 14267
rect 9676 14233 9710 14267
rect 9604 14155 9638 14189
rect 9676 14155 9710 14189
rect 9604 14077 9638 14111
rect 9676 14077 9710 14111
rect 9604 13999 9638 14033
rect 9676 13999 9710 14033
rect 9604 13921 9638 13955
rect 9676 13921 9710 13955
rect 9604 13843 9638 13877
rect 9676 13843 9710 13877
rect 9604 13765 9638 13799
rect 9676 13765 9710 13799
rect 9604 13688 9638 13722
rect 9676 13688 9710 13722
rect 9604 13611 9638 13645
rect 9676 13611 9710 13645
rect 9604 13534 9638 13568
rect 9676 13534 9710 13568
rect 9604 13457 9638 13491
rect 9676 13457 9710 13491
rect 9604 13380 9638 13414
rect 9676 13380 9710 13414
rect 9881 14311 9915 14345
rect 9953 14311 9987 14345
rect 9881 14233 9915 14267
rect 9953 14233 9987 14267
rect 9881 14155 9915 14189
rect 9953 14155 9987 14189
rect 9881 14077 9915 14111
rect 9953 14077 9987 14111
rect 9881 13999 9915 14033
rect 9953 13999 9987 14033
rect 9881 13921 9915 13955
rect 9953 13921 9987 13955
rect 9881 13843 9915 13877
rect 9953 13843 9987 13877
rect 9881 13765 9915 13799
rect 9953 13765 9987 13799
rect 9881 13688 9915 13722
rect 9953 13688 9987 13722
rect 9881 13611 9915 13645
rect 9953 13611 9987 13645
rect 9881 13534 9915 13568
rect 9953 13534 9987 13568
rect 9881 13457 9915 13491
rect 9953 13457 9987 13491
rect 9881 13380 9915 13414
rect 9953 13380 9987 13414
rect 10158 14311 10192 14345
rect 10230 14311 10264 14345
rect 10158 14233 10192 14267
rect 10230 14233 10264 14267
rect 10158 14155 10192 14189
rect 10230 14155 10264 14189
rect 10158 14077 10192 14111
rect 10230 14077 10264 14111
rect 10158 13999 10192 14033
rect 10230 13999 10264 14033
rect 10158 13921 10192 13955
rect 10230 13921 10264 13955
rect 10158 13843 10192 13877
rect 10230 13843 10264 13877
rect 10158 13765 10192 13799
rect 10230 13765 10264 13799
rect 10158 13688 10192 13722
rect 10230 13688 10264 13722
rect 10158 13611 10192 13645
rect 10230 13611 10264 13645
rect 10158 13534 10192 13568
rect 10230 13534 10264 13568
rect 10158 13457 10192 13491
rect 10230 13457 10264 13491
rect 10158 13380 10192 13414
rect 10230 13380 10264 13414
rect 10435 14311 10469 14345
rect 10507 14311 10541 14345
rect 10435 14233 10469 14267
rect 10507 14233 10541 14267
rect 10435 14155 10469 14189
rect 10507 14155 10541 14189
rect 10435 14077 10469 14111
rect 10507 14077 10541 14111
rect 10435 13999 10469 14033
rect 10507 13999 10541 14033
rect 10435 13921 10469 13955
rect 10507 13921 10541 13955
rect 10435 13843 10469 13877
rect 10507 13843 10541 13877
rect 10435 13765 10469 13799
rect 10507 13765 10541 13799
rect 10435 13688 10469 13722
rect 10507 13688 10541 13722
rect 10435 13611 10469 13645
rect 10507 13611 10541 13645
rect 10435 13534 10469 13568
rect 10507 13534 10541 13568
rect 10435 13457 10469 13491
rect 10507 13457 10541 13491
rect 10435 13380 10469 13414
rect 10507 13380 10541 13414
rect 10712 14311 10746 14345
rect 10784 14311 10818 14345
rect 10712 14233 10746 14267
rect 10784 14233 10818 14267
rect 10712 14155 10746 14189
rect 10784 14155 10818 14189
rect 10712 14077 10746 14111
rect 10784 14077 10818 14111
rect 10712 13999 10746 14033
rect 10784 13999 10818 14033
rect 10712 13921 10746 13955
rect 10784 13921 10818 13955
rect 10712 13843 10746 13877
rect 10784 13843 10818 13877
rect 10712 13765 10746 13799
rect 10784 13765 10818 13799
rect 10712 13688 10746 13722
rect 10784 13688 10818 13722
rect 10712 13611 10746 13645
rect 10784 13611 10818 13645
rect 10712 13534 10746 13568
rect 10784 13534 10818 13568
rect 10712 13457 10746 13491
rect 10784 13457 10818 13491
rect 10712 13380 10746 13414
rect 10784 13380 10818 13414
rect 10989 14311 11023 14345
rect 11061 14311 11095 14345
rect 10989 14233 11023 14267
rect 11061 14233 11095 14267
rect 10989 14155 11023 14189
rect 11061 14155 11095 14189
rect 10989 14077 11023 14111
rect 11061 14077 11095 14111
rect 10989 13999 11023 14033
rect 11061 13999 11095 14033
rect 10989 13921 11023 13955
rect 11061 13921 11095 13955
rect 10989 13843 11023 13877
rect 11061 13843 11095 13877
rect 10989 13765 11023 13799
rect 11061 13765 11095 13799
rect 10989 13688 11023 13722
rect 11061 13688 11095 13722
rect 10989 13611 11023 13645
rect 11061 13611 11095 13645
rect 10989 13534 11023 13568
rect 11061 13534 11095 13568
rect 10989 13457 11023 13491
rect 11061 13457 11095 13491
rect 10989 13380 11023 13414
rect 11061 13380 11095 13414
rect 11266 14311 11300 14345
rect 11338 14311 11372 14345
rect 11266 14233 11300 14267
rect 11338 14233 11372 14267
rect 11266 14155 11300 14189
rect 11338 14155 11372 14189
rect 11266 14077 11300 14111
rect 11338 14077 11372 14111
rect 11266 13999 11300 14033
rect 11338 13999 11372 14033
rect 11266 13921 11300 13955
rect 11338 13921 11372 13955
rect 11266 13843 11300 13877
rect 11338 13843 11372 13877
rect 11266 13765 11300 13799
rect 11338 13765 11372 13799
rect 11266 13688 11300 13722
rect 11338 13688 11372 13722
rect 11266 13611 11300 13645
rect 11338 13611 11372 13645
rect 11266 13534 11300 13568
rect 11338 13534 11372 13568
rect 11266 13457 11300 13491
rect 11338 13457 11372 13491
rect 11266 13380 11300 13414
rect 11338 13380 11372 13414
rect 11543 14311 11577 14345
rect 11615 14311 11649 14345
rect 11543 14233 11577 14267
rect 11615 14233 11649 14267
rect 11543 14155 11577 14189
rect 11615 14155 11649 14189
rect 11543 14077 11577 14111
rect 11615 14077 11649 14111
rect 11543 13999 11577 14033
rect 11615 13999 11649 14033
rect 11543 13921 11577 13955
rect 11615 13921 11649 13955
rect 11543 13843 11577 13877
rect 11615 13843 11649 13877
rect 11543 13765 11577 13799
rect 11615 13765 11649 13799
rect 11543 13688 11577 13722
rect 11615 13688 11649 13722
rect 11543 13611 11577 13645
rect 11615 13611 11649 13645
rect 11543 13534 11577 13568
rect 11615 13534 11649 13568
rect 11543 13457 11577 13491
rect 11615 13457 11649 13491
rect 11543 13380 11577 13414
rect 11615 13380 11649 13414
rect 11820 14311 11854 14345
rect 11892 14311 11926 14345
rect 11820 14233 11854 14267
rect 11892 14233 11926 14267
rect 11820 14155 11854 14189
rect 11892 14155 11926 14189
rect 11820 14077 11854 14111
rect 11892 14077 11926 14111
rect 11820 13999 11854 14033
rect 11892 13999 11926 14033
rect 11820 13921 11854 13955
rect 11892 13921 11926 13955
rect 11820 13843 11854 13877
rect 11892 13843 11926 13877
rect 11820 13765 11854 13799
rect 11892 13765 11926 13799
rect 11820 13688 11854 13722
rect 11892 13688 11926 13722
rect 11820 13611 11854 13645
rect 11892 13611 11926 13645
rect 11820 13534 11854 13568
rect 11892 13534 11926 13568
rect 11820 13457 11854 13491
rect 11892 13457 11926 13491
rect 11820 13380 11854 13414
rect 11892 13380 11926 13414
rect 12097 14311 12131 14345
rect 12169 14311 12203 14345
rect 12097 14233 12131 14267
rect 12169 14233 12203 14267
rect 12097 14155 12131 14189
rect 12169 14155 12203 14189
rect 12097 14077 12131 14111
rect 12169 14077 12203 14111
rect 12097 13999 12131 14033
rect 12169 13999 12203 14033
rect 12097 13921 12131 13955
rect 12169 13921 12203 13955
rect 12097 13843 12131 13877
rect 12169 13843 12203 13877
rect 12097 13765 12131 13799
rect 12169 13765 12203 13799
rect 12097 13688 12131 13722
rect 12169 13688 12203 13722
rect 12097 13611 12131 13645
rect 12169 13611 12203 13645
rect 12097 13534 12131 13568
rect 12169 13534 12203 13568
rect 12097 13457 12131 13491
rect 12169 13457 12203 13491
rect 12097 13380 12131 13414
rect 12169 13380 12203 13414
rect 12374 14311 12408 14345
rect 12446 14311 12480 14345
rect 12374 14233 12408 14267
rect 12446 14233 12480 14267
rect 12374 14155 12408 14189
rect 12446 14155 12480 14189
rect 12374 14077 12408 14111
rect 12446 14077 12480 14111
rect 12374 13999 12408 14033
rect 12446 13999 12480 14033
rect 12374 13921 12408 13955
rect 12446 13921 12480 13955
rect 12374 13843 12408 13877
rect 12446 13843 12480 13877
rect 12374 13765 12408 13799
rect 12446 13765 12480 13799
rect 12374 13688 12408 13722
rect 12446 13688 12480 13722
rect 12374 13611 12408 13645
rect 12446 13611 12480 13645
rect 12374 13534 12408 13568
rect 12446 13534 12480 13568
rect 12374 13457 12408 13491
rect 12446 13457 12480 13491
rect 12374 13380 12408 13414
rect 12446 13380 12480 13414
rect 12651 14311 12685 14345
rect 12723 14311 12757 14345
rect 12651 14233 12685 14267
rect 12723 14233 12757 14267
rect 12651 14155 12685 14189
rect 12723 14155 12757 14189
rect 12651 14077 12685 14111
rect 12723 14077 12757 14111
rect 12651 13999 12685 14033
rect 12723 13999 12757 14033
rect 12651 13921 12685 13955
rect 12723 13921 12757 13955
rect 12651 13843 12685 13877
rect 12723 13843 12757 13877
rect 12651 13765 12685 13799
rect 12723 13765 12757 13799
rect 12651 13688 12685 13722
rect 12723 13688 12757 13722
rect 12651 13611 12685 13645
rect 12723 13611 12757 13645
rect 12651 13534 12685 13568
rect 12723 13534 12757 13568
rect 12651 13457 12685 13491
rect 12723 13457 12757 13491
rect 12651 13380 12685 13414
rect 12723 13380 12757 13414
rect 12928 14311 12962 14345
rect 13000 14311 13034 14345
rect 12928 14233 12962 14267
rect 13000 14233 13034 14267
rect 12928 14155 12962 14189
rect 13000 14155 13034 14189
rect 12928 14077 12962 14111
rect 13000 14077 13034 14111
rect 12928 13999 12962 14033
rect 13000 13999 13034 14033
rect 12928 13921 12962 13955
rect 13000 13921 13034 13955
rect 12928 13843 12962 13877
rect 13000 13843 13034 13877
rect 12928 13765 12962 13799
rect 13000 13765 13034 13799
rect 12928 13688 12962 13722
rect 13000 13688 13034 13722
rect 12928 13611 12962 13645
rect 13000 13611 13034 13645
rect 12928 13534 12962 13568
rect 13000 13534 13034 13568
rect 12928 13457 12962 13491
rect 13000 13457 13034 13491
rect 12928 13380 12962 13414
rect 13000 13380 13034 13414
rect 13205 14311 13239 14345
rect 13277 14311 13311 14345
rect 13205 14233 13239 14267
rect 13277 14233 13311 14267
rect 13205 14155 13239 14189
rect 13277 14155 13311 14189
rect 13205 14077 13239 14111
rect 13277 14077 13311 14111
rect 13205 13999 13239 14033
rect 13277 13999 13311 14033
rect 13205 13921 13239 13955
rect 13277 13921 13311 13955
rect 13205 13843 13239 13877
rect 13277 13843 13311 13877
rect 13205 13765 13239 13799
rect 13277 13765 13311 13799
rect 13205 13688 13239 13722
rect 13277 13688 13311 13722
rect 13205 13611 13239 13645
rect 13277 13611 13311 13645
rect 13205 13534 13239 13568
rect 13277 13534 13311 13568
rect 13205 13457 13239 13491
rect 13277 13457 13311 13491
rect 13205 13380 13239 13414
rect 13277 13380 13311 13414
rect 2280 13298 2314 13332
rect 2404 13298 2438 13332
rect 2669 13184 2703 13218
rect 2741 13184 2775 13218
rect 2669 13077 2703 13111
rect 2741 13077 2775 13111
rect 2669 12970 2703 13004
rect 2741 12970 2775 13004
rect 2255 11891 2274 12789
rect 2274 11891 2361 12789
rect 2255 11818 2274 11852
rect 2274 11818 2289 11852
rect 2327 11818 2361 11852
rect 2255 11745 2274 11779
rect 2274 11745 2289 11779
rect 2327 11745 2361 11779
rect 2255 11672 2274 11706
rect 2274 11672 2289 11706
rect 2327 11672 2361 11706
rect 2255 11599 2274 11633
rect 2274 11599 2289 11633
rect 2327 11599 2361 11633
rect 2255 11526 2274 11560
rect 2274 11526 2289 11560
rect 2327 11526 2361 11560
rect 2255 11453 2274 11487
rect 2274 11453 2289 11487
rect 2327 11453 2361 11487
rect 2255 11380 2274 11414
rect 2274 11380 2289 11414
rect 2327 11380 2361 11414
rect 2679 12680 2713 12714
rect 2751 12680 2785 12714
rect 2679 12607 2713 12641
rect 2751 12607 2785 12641
rect 2679 12534 2713 12568
rect 2751 12534 2785 12568
rect 2679 12461 2713 12495
rect 2751 12461 2785 12495
rect 2679 11380 2785 12422
rect 2956 12680 2990 12714
rect 3028 12680 3062 12714
rect 2956 12607 2990 12641
rect 3028 12607 3062 12641
rect 2956 12534 2990 12568
rect 3028 12534 3062 12568
rect 2956 12461 2990 12495
rect 3028 12461 3062 12495
rect 2956 11380 3062 12422
rect 3233 12680 3267 12714
rect 3305 12680 3339 12714
rect 3233 12607 3267 12641
rect 3305 12607 3339 12641
rect 3233 12534 3267 12568
rect 3305 12534 3339 12568
rect 3233 12461 3267 12495
rect 3305 12461 3339 12495
rect 3233 11380 3339 12422
rect 3510 12680 3544 12714
rect 3582 12680 3616 12714
rect 3510 12607 3544 12641
rect 3582 12607 3616 12641
rect 3510 12534 3544 12568
rect 3582 12534 3616 12568
rect 3510 12461 3544 12495
rect 3582 12461 3616 12495
rect 3510 11380 3616 12422
rect 3787 12680 3821 12714
rect 3859 12680 3893 12714
rect 3787 12607 3821 12641
rect 3859 12607 3893 12641
rect 3787 12534 3821 12568
rect 3859 12534 3893 12568
rect 3787 12461 3821 12495
rect 3859 12461 3893 12495
rect 3787 11380 3893 12422
rect 4064 12680 4098 12714
rect 4136 12680 4170 12714
rect 4064 12607 4098 12641
rect 4136 12607 4170 12641
rect 4064 12534 4098 12568
rect 4136 12534 4170 12568
rect 4064 12461 4098 12495
rect 4136 12461 4170 12495
rect 4064 11380 4170 12422
rect 4341 12680 4375 12714
rect 4413 12680 4447 12714
rect 4341 12607 4375 12641
rect 4413 12607 4447 12641
rect 4341 12534 4375 12568
rect 4413 12534 4447 12568
rect 4341 12461 4375 12495
rect 4413 12461 4447 12495
rect 4341 11380 4447 12422
rect 4618 12680 4652 12714
rect 4690 12680 4724 12714
rect 4618 12607 4652 12641
rect 4690 12607 4724 12641
rect 4618 12534 4652 12568
rect 4690 12534 4724 12568
rect 4618 12461 4652 12495
rect 4690 12461 4724 12495
rect 4618 11380 4724 12422
rect 4895 12680 4929 12714
rect 4967 12680 5001 12714
rect 4895 12607 4929 12641
rect 4967 12607 5001 12641
rect 4895 12534 4929 12568
rect 4967 12534 5001 12568
rect 4895 12461 4929 12495
rect 4967 12461 5001 12495
rect 4895 11380 5001 12422
rect 5172 12680 5206 12714
rect 5244 12680 5278 12714
rect 5172 12607 5206 12641
rect 5244 12607 5278 12641
rect 5172 12534 5206 12568
rect 5244 12534 5278 12568
rect 5172 12461 5206 12495
rect 5244 12461 5278 12495
rect 5172 11380 5278 12422
rect 5449 12680 5483 12714
rect 5521 12680 5555 12714
rect 5449 12607 5483 12641
rect 5521 12607 5555 12641
rect 5449 12534 5483 12568
rect 5521 12534 5555 12568
rect 5449 12461 5483 12495
rect 5521 12461 5555 12495
rect 5449 11380 5555 12422
rect 5726 12680 5760 12714
rect 5798 12680 5832 12714
rect 5726 12607 5760 12641
rect 5798 12607 5832 12641
rect 5726 12534 5760 12568
rect 5798 12534 5832 12568
rect 5726 12461 5760 12495
rect 5798 12461 5832 12495
rect 5726 11380 5832 12422
rect 6003 12680 6037 12714
rect 6075 12680 6109 12714
rect 6003 12607 6037 12641
rect 6075 12607 6109 12641
rect 6003 12534 6037 12568
rect 6075 12534 6109 12568
rect 6003 12461 6037 12495
rect 6075 12461 6109 12495
rect 6003 11380 6109 12422
rect 6280 12680 6314 12714
rect 6352 12680 6386 12714
rect 6280 12607 6314 12641
rect 6352 12607 6386 12641
rect 6280 12534 6314 12568
rect 6352 12534 6386 12568
rect 6280 12461 6314 12495
rect 6352 12461 6386 12495
rect 6280 11380 6386 12422
rect 6557 12680 6591 12714
rect 6629 12680 6663 12714
rect 6557 12607 6591 12641
rect 6629 12607 6663 12641
rect 6557 12534 6591 12568
rect 6629 12534 6663 12568
rect 6557 12461 6591 12495
rect 6629 12461 6663 12495
rect 6557 11380 6663 12422
rect 6834 12680 6868 12714
rect 6906 12680 6940 12714
rect 6834 12607 6868 12641
rect 6906 12607 6940 12641
rect 6834 12534 6868 12568
rect 6906 12534 6940 12568
rect 6834 12461 6868 12495
rect 6906 12461 6940 12495
rect 6834 11380 6940 12422
rect 7111 12680 7145 12714
rect 7183 12680 7217 12714
rect 7111 12607 7145 12641
rect 7183 12607 7217 12641
rect 7111 12534 7145 12568
rect 7183 12534 7217 12568
rect 7111 12461 7145 12495
rect 7183 12461 7217 12495
rect 7111 11380 7217 12422
rect 7388 12680 7422 12714
rect 7460 12680 7494 12714
rect 7388 12607 7422 12641
rect 7460 12607 7494 12641
rect 7388 12534 7422 12568
rect 7460 12534 7494 12568
rect 7388 12461 7422 12495
rect 7460 12461 7494 12495
rect 7388 11380 7494 12422
rect 7665 12680 7699 12714
rect 7737 12680 7771 12714
rect 7665 12607 7699 12641
rect 7737 12607 7771 12641
rect 7665 12534 7699 12568
rect 7737 12534 7771 12568
rect 7665 12461 7699 12495
rect 7737 12461 7771 12495
rect 7665 11380 7771 12422
rect 7942 12680 7976 12714
rect 8014 12680 8048 12714
rect 7942 12607 7976 12641
rect 8014 12607 8048 12641
rect 7942 12534 7976 12568
rect 8014 12534 8048 12568
rect 7942 12461 7976 12495
rect 8014 12461 8048 12495
rect 7942 11380 8048 12422
rect 8219 12680 8253 12714
rect 8291 12680 8325 12714
rect 8219 12607 8253 12641
rect 8291 12607 8325 12641
rect 8219 12534 8253 12568
rect 8291 12534 8325 12568
rect 8219 12461 8253 12495
rect 8291 12461 8325 12495
rect 8219 11380 8325 12422
rect 8496 12680 8530 12714
rect 8568 12680 8602 12714
rect 8496 12607 8530 12641
rect 8568 12607 8602 12641
rect 8496 12534 8530 12568
rect 8568 12534 8602 12568
rect 8496 12461 8530 12495
rect 8568 12461 8602 12495
rect 8496 11380 8602 12422
rect 8773 12680 8807 12714
rect 8845 12680 8879 12714
rect 8773 12607 8807 12641
rect 8845 12607 8879 12641
rect 8773 12534 8807 12568
rect 8845 12534 8879 12568
rect 8773 12461 8807 12495
rect 8845 12461 8879 12495
rect 8773 11380 8879 12422
rect 9050 12680 9084 12714
rect 9122 12680 9156 12714
rect 9050 12607 9084 12641
rect 9122 12607 9156 12641
rect 9050 12534 9084 12568
rect 9122 12534 9156 12568
rect 9050 12461 9084 12495
rect 9122 12461 9156 12495
rect 9050 11380 9156 12422
rect 9327 12680 9361 12714
rect 9399 12680 9433 12714
rect 9327 12607 9361 12641
rect 9399 12607 9433 12641
rect 9327 12534 9361 12568
rect 9399 12534 9433 12568
rect 9327 12461 9361 12495
rect 9399 12461 9433 12495
rect 9327 11380 9433 12422
rect 9604 12680 9638 12714
rect 9676 12680 9710 12714
rect 9604 12607 9638 12641
rect 9676 12607 9710 12641
rect 9604 12534 9638 12568
rect 9676 12534 9710 12568
rect 9604 12461 9638 12495
rect 9676 12461 9710 12495
rect 9604 11380 9710 12422
rect 9881 12680 9915 12714
rect 9953 12680 9987 12714
rect 9881 12607 9915 12641
rect 9953 12607 9987 12641
rect 9881 12534 9915 12568
rect 9953 12534 9987 12568
rect 9881 12461 9915 12495
rect 9953 12461 9987 12495
rect 9881 11380 9987 12422
rect 10158 12680 10192 12714
rect 10230 12680 10264 12714
rect 10158 12607 10192 12641
rect 10230 12607 10264 12641
rect 10158 12534 10192 12568
rect 10230 12534 10264 12568
rect 10158 12461 10192 12495
rect 10230 12461 10264 12495
rect 10158 11380 10264 12422
rect 10435 12680 10469 12714
rect 10507 12680 10541 12714
rect 10435 12607 10469 12641
rect 10507 12607 10541 12641
rect 10435 12534 10469 12568
rect 10507 12534 10541 12568
rect 10435 12461 10469 12495
rect 10507 12461 10541 12495
rect 10435 11380 10541 12422
rect 10712 12680 10746 12714
rect 10784 12680 10818 12714
rect 10712 12607 10746 12641
rect 10784 12607 10818 12641
rect 10712 12534 10746 12568
rect 10784 12534 10818 12568
rect 10712 12461 10746 12495
rect 10784 12461 10818 12495
rect 10712 11380 10818 12422
rect 10989 12680 11023 12714
rect 11061 12680 11095 12714
rect 10989 12607 11023 12641
rect 11061 12607 11095 12641
rect 10989 12534 11023 12568
rect 11061 12534 11095 12568
rect 10989 12461 11023 12495
rect 11061 12461 11095 12495
rect 10989 11380 11095 12422
rect 11266 12680 11300 12714
rect 11338 12680 11372 12714
rect 11266 12607 11300 12641
rect 11338 12607 11372 12641
rect 11266 12534 11300 12568
rect 11338 12534 11372 12568
rect 11266 12461 11300 12495
rect 11338 12461 11372 12495
rect 11266 11380 11372 12422
rect 11543 12680 11577 12714
rect 11615 12680 11649 12714
rect 11543 12607 11577 12641
rect 11615 12607 11649 12641
rect 11543 12534 11577 12568
rect 11615 12534 11649 12568
rect 11543 12461 11577 12495
rect 11615 12461 11649 12495
rect 11543 11380 11649 12422
rect 11820 12680 11854 12714
rect 11892 12680 11926 12714
rect 11820 12607 11854 12641
rect 11892 12607 11926 12641
rect 11820 12534 11854 12568
rect 11892 12534 11926 12568
rect 11820 12461 11854 12495
rect 11892 12461 11926 12495
rect 11820 11380 11926 12422
rect 12097 12680 12131 12714
rect 12169 12680 12203 12714
rect 12097 12607 12131 12641
rect 12169 12607 12203 12641
rect 12097 12534 12131 12568
rect 12169 12534 12203 12568
rect 12097 12461 12131 12495
rect 12169 12461 12203 12495
rect 12097 11380 12203 12422
rect 12374 12680 12408 12714
rect 12446 12680 12480 12714
rect 12374 12607 12408 12641
rect 12446 12607 12480 12641
rect 12374 12534 12408 12568
rect 12446 12534 12480 12568
rect 12374 12461 12408 12495
rect 12446 12461 12480 12495
rect 12374 11380 12480 12422
rect 12651 12680 12685 12714
rect 12723 12680 12757 12714
rect 12651 12607 12685 12641
rect 12723 12607 12757 12641
rect 12651 12534 12685 12568
rect 12723 12534 12757 12568
rect 12651 12461 12685 12495
rect 12723 12461 12757 12495
rect 12651 11380 12757 12422
rect 12928 12680 12962 12714
rect 13000 12680 13034 12714
rect 12928 12607 12962 12641
rect 13000 12607 13034 12641
rect 12928 12534 12962 12568
rect 13000 12534 13034 12568
rect 12928 12461 12962 12495
rect 13000 12461 13034 12495
rect 12928 11380 13034 12422
rect 13205 12680 13239 12714
rect 13277 12680 13311 12714
rect 13205 12607 13239 12641
rect 13277 12607 13311 12641
rect 13205 12534 13239 12568
rect 13277 12534 13311 12568
rect 13205 12461 13239 12495
rect 13277 12461 13311 12495
rect 13205 11380 13311 12422
rect 2638 11160 2672 11194
rect 2710 11160 2744 11194
rect 2638 11053 2672 11087
rect 2710 11053 2744 11087
rect 2638 10946 2672 10980
rect 2710 10946 2744 10980
rect 2255 9600 2274 10714
rect 2274 9600 2361 10714
rect 2255 9527 2274 9561
rect 2274 9527 2289 9561
rect 2327 9527 2361 9561
rect 2255 9454 2274 9488
rect 2274 9454 2289 9488
rect 2327 9454 2361 9488
rect 2255 9381 2274 9415
rect 2274 9381 2289 9415
rect 2327 9381 2361 9415
rect 1944 7618 1946 8732
rect 1946 7618 2048 8732
rect 2048 7618 2050 8732
rect 2679 10680 2713 10714
rect 2751 10680 2785 10714
rect 2679 10607 2713 10641
rect 2751 10607 2785 10641
rect 2679 10534 2713 10568
rect 2751 10534 2785 10568
rect 2679 10461 2713 10495
rect 2751 10461 2785 10495
rect 2679 9380 2785 10422
rect 2956 10680 2990 10714
rect 3028 10680 3062 10714
rect 2956 10607 2990 10641
rect 3028 10607 3062 10641
rect 2956 10534 2990 10568
rect 3028 10534 3062 10568
rect 2956 10461 2990 10495
rect 3028 10461 3062 10495
rect 2956 9380 3062 10422
rect 3233 10680 3267 10714
rect 3305 10680 3339 10714
rect 3233 10607 3267 10641
rect 3305 10607 3339 10641
rect 3233 10534 3267 10568
rect 3305 10534 3339 10568
rect 3233 10461 3267 10495
rect 3305 10461 3339 10495
rect 3233 9380 3339 10422
rect 3510 10680 3544 10714
rect 3582 10680 3616 10714
rect 3510 10607 3544 10641
rect 3582 10607 3616 10641
rect 3510 10534 3544 10568
rect 3582 10534 3616 10568
rect 3510 10461 3544 10495
rect 3582 10461 3616 10495
rect 3510 9380 3616 10422
rect 3787 10680 3821 10714
rect 3859 10680 3893 10714
rect 3787 10607 3821 10641
rect 3859 10607 3893 10641
rect 3787 10534 3821 10568
rect 3859 10534 3893 10568
rect 3787 10461 3821 10495
rect 3859 10461 3893 10495
rect 3787 9380 3893 10422
rect 4064 10680 4098 10714
rect 4136 10680 4170 10714
rect 4064 10607 4098 10641
rect 4136 10607 4170 10641
rect 4064 10534 4098 10568
rect 4136 10534 4170 10568
rect 4064 10461 4098 10495
rect 4136 10461 4170 10495
rect 4064 9380 4170 10422
rect 4341 10680 4375 10714
rect 4413 10680 4447 10714
rect 4341 10607 4375 10641
rect 4413 10607 4447 10641
rect 4341 10534 4375 10568
rect 4413 10534 4447 10568
rect 4341 10461 4375 10495
rect 4413 10461 4447 10495
rect 4341 9380 4447 10422
rect 4618 10680 4652 10714
rect 4690 10680 4724 10714
rect 4618 10607 4652 10641
rect 4690 10607 4724 10641
rect 4618 10534 4652 10568
rect 4690 10534 4724 10568
rect 4618 10461 4652 10495
rect 4690 10461 4724 10495
rect 4618 9380 4724 10422
rect 4895 10680 4929 10714
rect 4967 10680 5001 10714
rect 4895 10607 4929 10641
rect 4967 10607 5001 10641
rect 4895 10534 4929 10568
rect 4967 10534 5001 10568
rect 4895 10461 4929 10495
rect 4967 10461 5001 10495
rect 4895 9380 5001 10422
rect 5172 10680 5206 10714
rect 5244 10680 5278 10714
rect 5172 10607 5206 10641
rect 5244 10607 5278 10641
rect 5172 10534 5206 10568
rect 5244 10534 5278 10568
rect 5172 10461 5206 10495
rect 5244 10461 5278 10495
rect 5172 9380 5278 10422
rect 5449 10680 5483 10714
rect 5521 10680 5555 10714
rect 5449 10607 5483 10641
rect 5521 10607 5555 10641
rect 5449 10534 5483 10568
rect 5521 10534 5555 10568
rect 5449 10461 5483 10495
rect 5521 10461 5555 10495
rect 5449 9380 5555 10422
rect 5726 10680 5760 10714
rect 5798 10680 5832 10714
rect 5726 10607 5760 10641
rect 5798 10607 5832 10641
rect 5726 10534 5760 10568
rect 5798 10534 5832 10568
rect 5726 10461 5760 10495
rect 5798 10461 5832 10495
rect 5726 9380 5832 10422
rect 6003 10680 6037 10714
rect 6075 10680 6109 10714
rect 6003 10607 6037 10641
rect 6075 10607 6109 10641
rect 6003 10534 6037 10568
rect 6075 10534 6109 10568
rect 6003 10461 6037 10495
rect 6075 10461 6109 10495
rect 6003 9380 6109 10422
rect 6280 10680 6314 10714
rect 6352 10680 6386 10714
rect 6280 10607 6314 10641
rect 6352 10607 6386 10641
rect 6280 10534 6314 10568
rect 6352 10534 6386 10568
rect 6280 10461 6314 10495
rect 6352 10461 6386 10495
rect 6280 9380 6386 10422
rect 6557 10680 6591 10714
rect 6629 10680 6663 10714
rect 6557 10607 6591 10641
rect 6629 10607 6663 10641
rect 6557 10534 6591 10568
rect 6629 10534 6663 10568
rect 6557 10461 6591 10495
rect 6629 10461 6663 10495
rect 6557 9380 6663 10422
rect 6834 10680 6868 10714
rect 6906 10680 6940 10714
rect 6834 10607 6868 10641
rect 6906 10607 6940 10641
rect 6834 10534 6868 10568
rect 6906 10534 6940 10568
rect 6834 10461 6868 10495
rect 6906 10461 6940 10495
rect 6834 9380 6940 10422
rect 7111 10680 7145 10714
rect 7183 10680 7217 10714
rect 7111 10607 7145 10641
rect 7183 10607 7217 10641
rect 7111 10534 7145 10568
rect 7183 10534 7217 10568
rect 7111 10461 7145 10495
rect 7183 10461 7217 10495
rect 7111 9380 7217 10422
rect 7388 10680 7422 10714
rect 7460 10680 7494 10714
rect 7388 10607 7422 10641
rect 7460 10607 7494 10641
rect 7388 10534 7422 10568
rect 7460 10534 7494 10568
rect 7388 10461 7422 10495
rect 7460 10461 7494 10495
rect 7388 9380 7494 10422
rect 7665 10680 7699 10714
rect 7737 10680 7771 10714
rect 7665 10607 7699 10641
rect 7737 10607 7771 10641
rect 7665 10534 7699 10568
rect 7737 10534 7771 10568
rect 7665 10461 7699 10495
rect 7737 10461 7771 10495
rect 7665 9380 7771 10422
rect 7942 10680 7976 10714
rect 8014 10680 8048 10714
rect 7942 10607 7976 10641
rect 8014 10607 8048 10641
rect 7942 10534 7976 10568
rect 8014 10534 8048 10568
rect 7942 10461 7976 10495
rect 8014 10461 8048 10495
rect 7942 9380 8048 10422
rect 8219 10680 8253 10714
rect 8291 10680 8325 10714
rect 8219 10607 8253 10641
rect 8291 10607 8325 10641
rect 8219 10534 8253 10568
rect 8291 10534 8325 10568
rect 8219 10461 8253 10495
rect 8291 10461 8325 10495
rect 8219 9380 8325 10422
rect 8496 10680 8530 10714
rect 8568 10680 8602 10714
rect 8496 10607 8530 10641
rect 8568 10607 8602 10641
rect 8496 10534 8530 10568
rect 8568 10534 8602 10568
rect 8496 10461 8530 10495
rect 8568 10461 8602 10495
rect 8496 9380 8602 10422
rect 8773 10680 8807 10714
rect 8845 10680 8879 10714
rect 8773 10607 8807 10641
rect 8845 10607 8879 10641
rect 8773 10534 8807 10568
rect 8845 10534 8879 10568
rect 8773 10461 8807 10495
rect 8845 10461 8879 10495
rect 8773 9380 8879 10422
rect 9050 10680 9084 10714
rect 9122 10680 9156 10714
rect 9050 10607 9084 10641
rect 9122 10607 9156 10641
rect 9050 10534 9084 10568
rect 9122 10534 9156 10568
rect 9050 10461 9084 10495
rect 9122 10461 9156 10495
rect 9050 9380 9156 10422
rect 9327 10680 9361 10714
rect 9399 10680 9433 10714
rect 9327 10607 9361 10641
rect 9399 10607 9433 10641
rect 9327 10534 9361 10568
rect 9399 10534 9433 10568
rect 9327 10461 9361 10495
rect 9399 10461 9433 10495
rect 9327 9380 9433 10422
rect 9604 10680 9638 10714
rect 9676 10680 9710 10714
rect 9604 10607 9638 10641
rect 9676 10607 9710 10641
rect 9604 10534 9638 10568
rect 9676 10534 9710 10568
rect 9604 10461 9638 10495
rect 9676 10461 9710 10495
rect 9604 9380 9710 10422
rect 9881 10680 9915 10714
rect 9953 10680 9987 10714
rect 9881 10607 9915 10641
rect 9953 10607 9987 10641
rect 9881 10534 9915 10568
rect 9953 10534 9987 10568
rect 9881 10461 9915 10495
rect 9953 10461 9987 10495
rect 9881 9380 9987 10422
rect 10158 10680 10192 10714
rect 10230 10680 10264 10714
rect 10158 10607 10192 10641
rect 10230 10607 10264 10641
rect 10158 10534 10192 10568
rect 10230 10534 10264 10568
rect 10158 10461 10192 10495
rect 10230 10461 10264 10495
rect 10158 9380 10264 10422
rect 10435 10680 10469 10714
rect 10507 10680 10541 10714
rect 10435 10607 10469 10641
rect 10507 10607 10541 10641
rect 10435 10534 10469 10568
rect 10507 10534 10541 10568
rect 10435 10461 10469 10495
rect 10507 10461 10541 10495
rect 10435 9380 10541 10422
rect 10712 10680 10746 10714
rect 10784 10680 10818 10714
rect 10712 10607 10746 10641
rect 10784 10607 10818 10641
rect 10712 10534 10746 10568
rect 10784 10534 10818 10568
rect 10712 10461 10746 10495
rect 10784 10461 10818 10495
rect 10712 9380 10818 10422
rect 10989 10680 11023 10714
rect 11061 10680 11095 10714
rect 10989 10607 11023 10641
rect 11061 10607 11095 10641
rect 10989 10534 11023 10568
rect 11061 10534 11095 10568
rect 10989 10461 11023 10495
rect 11061 10461 11095 10495
rect 10989 9380 11095 10422
rect 11266 10680 11300 10714
rect 11338 10680 11372 10714
rect 11266 10607 11300 10641
rect 11338 10607 11372 10641
rect 11266 10534 11300 10568
rect 11338 10534 11372 10568
rect 11266 10461 11300 10495
rect 11338 10461 11372 10495
rect 11266 9380 11372 10422
rect 11543 10680 11577 10714
rect 11615 10680 11649 10714
rect 11543 10607 11577 10641
rect 11615 10607 11649 10641
rect 11543 10534 11577 10568
rect 11615 10534 11649 10568
rect 11543 10461 11577 10495
rect 11615 10461 11649 10495
rect 11543 9380 11649 10422
rect 11820 10680 11854 10714
rect 11892 10680 11926 10714
rect 11820 10607 11854 10641
rect 11892 10607 11926 10641
rect 11820 10534 11854 10568
rect 11892 10534 11926 10568
rect 11820 10461 11854 10495
rect 11892 10461 11926 10495
rect 11820 9380 11926 10422
rect 12097 10680 12131 10714
rect 12169 10680 12203 10714
rect 12097 10607 12131 10641
rect 12169 10607 12203 10641
rect 12097 10534 12131 10568
rect 12169 10534 12203 10568
rect 12097 10461 12131 10495
rect 12169 10461 12203 10495
rect 12097 9380 12203 10422
rect 12374 10680 12408 10714
rect 12446 10680 12480 10714
rect 12374 10607 12408 10641
rect 12446 10607 12480 10641
rect 12374 10534 12408 10568
rect 12446 10534 12480 10568
rect 12374 10461 12408 10495
rect 12446 10461 12480 10495
rect 12374 9380 12480 10422
rect 12651 10680 12685 10714
rect 12723 10680 12757 10714
rect 12651 10607 12685 10641
rect 12723 10607 12757 10641
rect 12651 10534 12685 10568
rect 12723 10534 12757 10568
rect 12651 10461 12685 10495
rect 12723 10461 12757 10495
rect 12651 9380 12757 10422
rect 12928 10680 12962 10714
rect 13000 10680 13034 10714
rect 12928 10607 12962 10641
rect 13000 10607 13034 10641
rect 12928 10534 12962 10568
rect 13000 10534 13034 10568
rect 12928 10461 12962 10495
rect 13000 10461 13034 10495
rect 12928 9380 13034 10422
rect 13205 10680 13239 10714
rect 13277 10680 13311 10714
rect 13205 10607 13239 10641
rect 13277 10607 13311 10641
rect 13205 10534 13239 10568
rect 13277 10534 13311 10568
rect 13205 10461 13239 10495
rect 13277 10461 13311 10495
rect 13205 9380 13311 10422
rect 2612 9199 2646 9233
rect 2684 9199 2718 9233
rect 2612 9126 2646 9160
rect 2684 9126 2718 9160
rect 2612 9052 2646 9086
rect 2684 9052 2718 9086
rect 2612 8978 2646 9012
rect 2684 8978 2718 9012
rect 2612 8904 2646 8938
rect 2684 8904 2718 8938
rect 1944 7545 1946 7579
rect 1946 7545 1978 7579
rect 2016 7545 2048 7579
rect 2048 7545 2050 7579
rect 2255 8690 2274 8724
rect 2274 8690 2289 8724
rect 2327 8690 2361 8724
rect 2255 8617 2274 8651
rect 2274 8617 2289 8651
rect 2327 8617 2361 8651
rect 2255 8543 2274 8577
rect 2274 8543 2289 8577
rect 2327 8543 2361 8577
rect 2255 8469 2274 8503
rect 2274 8469 2289 8503
rect 2327 8469 2361 8503
rect 2255 8395 2274 8429
rect 2274 8395 2289 8429
rect 2327 8395 2361 8429
rect 2255 8321 2274 8355
rect 2274 8321 2289 8355
rect 2327 8321 2361 8355
rect 2255 8247 2274 8281
rect 2274 8247 2289 8281
rect 2327 8247 2361 8281
rect 2255 8173 2274 8207
rect 2274 8173 2289 8207
rect 2327 8173 2361 8207
rect 2255 8099 2274 8133
rect 2274 8099 2289 8133
rect 2327 8099 2361 8133
rect 2255 8025 2274 8059
rect 2274 8025 2289 8059
rect 2327 8025 2361 8059
rect 2255 7951 2274 7985
rect 2274 7951 2289 7985
rect 2327 7951 2361 7985
rect 2255 7877 2274 7911
rect 2274 7877 2289 7911
rect 2327 7877 2361 7911
rect 2255 7803 2274 7837
rect 2274 7803 2289 7837
rect 2327 7803 2361 7837
rect 2255 7729 2274 7763
rect 2274 7729 2289 7763
rect 2327 7729 2361 7763
rect 2255 7655 2274 7689
rect 2274 7655 2289 7689
rect 2327 7655 2361 7689
rect 2255 7581 2274 7615
rect 2274 7581 2289 7615
rect 2327 7581 2361 7615
rect 2255 7507 2274 7541
rect 2274 7507 2289 7541
rect 2327 7507 2361 7541
rect 2255 7433 2274 7467
rect 2274 7433 2289 7467
rect 2327 7433 2361 7467
rect 2255 7359 2274 7393
rect 2274 7359 2289 7393
rect 2327 7359 2361 7393
rect 2679 8680 2713 8714
rect 2751 8680 2785 8714
rect 2679 8607 2713 8641
rect 2751 8607 2785 8641
rect 2679 8534 2713 8568
rect 2751 8534 2785 8568
rect 2679 8461 2713 8495
rect 2751 8461 2785 8495
rect 2679 7380 2785 8422
rect 2956 8680 2990 8714
rect 3028 8680 3062 8714
rect 2956 8607 2990 8641
rect 3028 8607 3062 8641
rect 2956 8534 2990 8568
rect 3028 8534 3062 8568
rect 2956 8461 2990 8495
rect 3028 8461 3062 8495
rect 2956 7380 3062 8422
rect 3233 8680 3267 8714
rect 3305 8680 3339 8714
rect 3233 8607 3267 8641
rect 3305 8607 3339 8641
rect 3233 8534 3267 8568
rect 3305 8534 3339 8568
rect 3233 8461 3267 8495
rect 3305 8461 3339 8495
rect 3233 7380 3339 8422
rect 3510 8680 3544 8714
rect 3582 8680 3616 8714
rect 3510 8607 3544 8641
rect 3582 8607 3616 8641
rect 3510 8534 3544 8568
rect 3582 8534 3616 8568
rect 3510 8461 3544 8495
rect 3582 8461 3616 8495
rect 3510 7380 3616 8422
rect 3787 8680 3821 8714
rect 3859 8680 3893 8714
rect 3787 8607 3821 8641
rect 3859 8607 3893 8641
rect 3787 8534 3821 8568
rect 3859 8534 3893 8568
rect 3787 8461 3821 8495
rect 3859 8461 3893 8495
rect 3787 7380 3893 8422
rect 4064 8680 4098 8714
rect 4136 8680 4170 8714
rect 4064 8607 4098 8641
rect 4136 8607 4170 8641
rect 4064 8534 4098 8568
rect 4136 8534 4170 8568
rect 4064 8461 4098 8495
rect 4136 8461 4170 8495
rect 4064 7380 4170 8422
rect 4341 8680 4375 8714
rect 4413 8680 4447 8714
rect 4341 8607 4375 8641
rect 4413 8607 4447 8641
rect 4341 8534 4375 8568
rect 4413 8534 4447 8568
rect 4341 8461 4375 8495
rect 4413 8461 4447 8495
rect 4341 7380 4447 8422
rect 4618 8680 4652 8714
rect 4690 8680 4724 8714
rect 4618 8607 4652 8641
rect 4690 8607 4724 8641
rect 4618 8534 4652 8568
rect 4690 8534 4724 8568
rect 4618 8461 4652 8495
rect 4690 8461 4724 8495
rect 4618 7380 4724 8422
rect 4895 8680 4929 8714
rect 4967 8680 5001 8714
rect 4895 8607 4929 8641
rect 4967 8607 5001 8641
rect 4895 8534 4929 8568
rect 4967 8534 5001 8568
rect 4895 8461 4929 8495
rect 4967 8461 5001 8495
rect 4895 7380 5001 8422
rect 5172 8680 5206 8714
rect 5244 8680 5278 8714
rect 5172 8607 5206 8641
rect 5244 8607 5278 8641
rect 5172 8534 5206 8568
rect 5244 8534 5278 8568
rect 5172 8461 5206 8495
rect 5244 8461 5278 8495
rect 5172 7380 5278 8422
rect 5449 8680 5483 8714
rect 5521 8680 5555 8714
rect 5449 8607 5483 8641
rect 5521 8607 5555 8641
rect 5449 8534 5483 8568
rect 5521 8534 5555 8568
rect 5449 8461 5483 8495
rect 5521 8461 5555 8495
rect 5449 7380 5555 8422
rect 5726 8680 5760 8714
rect 5798 8680 5832 8714
rect 5726 8607 5760 8641
rect 5798 8607 5832 8641
rect 5726 8534 5760 8568
rect 5798 8534 5832 8568
rect 5726 8461 5760 8495
rect 5798 8461 5832 8495
rect 5726 7380 5832 8422
rect 6003 8680 6037 8714
rect 6075 8680 6109 8714
rect 6003 8607 6037 8641
rect 6075 8607 6109 8641
rect 6003 8534 6037 8568
rect 6075 8534 6109 8568
rect 6003 8461 6037 8495
rect 6075 8461 6109 8495
rect 6003 7380 6109 8422
rect 6280 8680 6314 8714
rect 6352 8680 6386 8714
rect 6280 8607 6314 8641
rect 6352 8607 6386 8641
rect 6280 8534 6314 8568
rect 6352 8534 6386 8568
rect 6280 8461 6314 8495
rect 6352 8461 6386 8495
rect 6280 7380 6386 8422
rect 6557 8680 6591 8714
rect 6629 8680 6663 8714
rect 6557 8607 6591 8641
rect 6629 8607 6663 8641
rect 6557 8534 6591 8568
rect 6629 8534 6663 8568
rect 6557 8461 6591 8495
rect 6629 8461 6663 8495
rect 6557 7380 6663 8422
rect 6834 8680 6868 8714
rect 6906 8680 6940 8714
rect 6834 8607 6868 8641
rect 6906 8607 6940 8641
rect 6834 8534 6868 8568
rect 6906 8534 6940 8568
rect 6834 8461 6868 8495
rect 6906 8461 6940 8495
rect 6834 7380 6940 8422
rect 7111 8680 7145 8714
rect 7183 8680 7217 8714
rect 7111 8607 7145 8641
rect 7183 8607 7217 8641
rect 7111 8534 7145 8568
rect 7183 8534 7217 8568
rect 7111 8461 7145 8495
rect 7183 8461 7217 8495
rect 7111 7380 7217 8422
rect 7388 8680 7422 8714
rect 7460 8680 7494 8714
rect 7388 8607 7422 8641
rect 7460 8607 7494 8641
rect 7388 8534 7422 8568
rect 7460 8534 7494 8568
rect 7388 8461 7422 8495
rect 7460 8461 7494 8495
rect 7388 7380 7494 8422
rect 7665 8680 7699 8714
rect 7737 8680 7771 8714
rect 7665 8607 7699 8641
rect 7737 8607 7771 8641
rect 7665 8534 7699 8568
rect 7737 8534 7771 8568
rect 7665 8461 7699 8495
rect 7737 8461 7771 8495
rect 7665 7380 7771 8422
rect 7942 8680 7976 8714
rect 8014 8680 8048 8714
rect 7942 8607 7976 8641
rect 8014 8607 8048 8641
rect 7942 8534 7976 8568
rect 8014 8534 8048 8568
rect 7942 8461 7976 8495
rect 8014 8461 8048 8495
rect 7942 7380 8048 8422
rect 8219 8680 8253 8714
rect 8291 8680 8325 8714
rect 8219 8607 8253 8641
rect 8291 8607 8325 8641
rect 8219 8534 8253 8568
rect 8291 8534 8325 8568
rect 8219 8461 8253 8495
rect 8291 8461 8325 8495
rect 8219 7380 8325 8422
rect 8496 8680 8530 8714
rect 8568 8680 8602 8714
rect 8496 8607 8530 8641
rect 8568 8607 8602 8641
rect 8496 8534 8530 8568
rect 8568 8534 8602 8568
rect 8496 8461 8530 8495
rect 8568 8461 8602 8495
rect 8496 7380 8602 8422
rect 8773 8680 8807 8714
rect 8845 8680 8879 8714
rect 8773 8607 8807 8641
rect 8845 8607 8879 8641
rect 8773 8534 8807 8568
rect 8845 8534 8879 8568
rect 8773 8461 8807 8495
rect 8845 8461 8879 8495
rect 8773 7380 8879 8422
rect 9050 8680 9084 8714
rect 9122 8680 9156 8714
rect 9050 8607 9084 8641
rect 9122 8607 9156 8641
rect 9050 8534 9084 8568
rect 9122 8534 9156 8568
rect 9050 8461 9084 8495
rect 9122 8461 9156 8495
rect 9050 7380 9156 8422
rect 9327 8680 9361 8714
rect 9399 8680 9433 8714
rect 9327 8607 9361 8641
rect 9399 8607 9433 8641
rect 9327 8534 9361 8568
rect 9399 8534 9433 8568
rect 9327 8461 9361 8495
rect 9399 8461 9433 8495
rect 9327 7380 9433 8422
rect 9604 8680 9638 8714
rect 9676 8680 9710 8714
rect 9604 8607 9638 8641
rect 9676 8607 9710 8641
rect 9604 8534 9638 8568
rect 9676 8534 9710 8568
rect 9604 8461 9638 8495
rect 9676 8461 9710 8495
rect 9604 7380 9710 8422
rect 9881 8680 9915 8714
rect 9953 8680 9987 8714
rect 9881 8607 9915 8641
rect 9953 8607 9987 8641
rect 9881 8534 9915 8568
rect 9953 8534 9987 8568
rect 9881 8461 9915 8495
rect 9953 8461 9987 8495
rect 9881 7380 9987 8422
rect 10158 8680 10192 8714
rect 10230 8680 10264 8714
rect 10158 8607 10192 8641
rect 10230 8607 10264 8641
rect 10158 8534 10192 8568
rect 10230 8534 10264 8568
rect 10158 8461 10192 8495
rect 10230 8461 10264 8495
rect 10158 7380 10264 8422
rect 10435 8680 10469 8714
rect 10507 8680 10541 8714
rect 10435 8607 10469 8641
rect 10507 8607 10541 8641
rect 10435 8534 10469 8568
rect 10507 8534 10541 8568
rect 10435 8461 10469 8495
rect 10507 8461 10541 8495
rect 10435 7380 10541 8422
rect 10712 8680 10746 8714
rect 10784 8680 10818 8714
rect 10712 8607 10746 8641
rect 10784 8607 10818 8641
rect 10712 8534 10746 8568
rect 10784 8534 10818 8568
rect 10712 8461 10746 8495
rect 10784 8461 10818 8495
rect 10712 7380 10818 8422
rect 10989 8680 11023 8714
rect 11061 8680 11095 8714
rect 10989 8607 11023 8641
rect 11061 8607 11095 8641
rect 10989 8534 11023 8568
rect 11061 8534 11095 8568
rect 10989 8461 11023 8495
rect 11061 8461 11095 8495
rect 10989 7380 11095 8422
rect 11266 8680 11300 8714
rect 11338 8680 11372 8714
rect 11266 8607 11300 8641
rect 11338 8607 11372 8641
rect 11266 8534 11300 8568
rect 11338 8534 11372 8568
rect 11266 8461 11300 8495
rect 11338 8461 11372 8495
rect 11266 7380 11372 8422
rect 11543 8680 11577 8714
rect 11615 8680 11649 8714
rect 11543 8607 11577 8641
rect 11615 8607 11649 8641
rect 11543 8534 11577 8568
rect 11615 8534 11649 8568
rect 11543 8461 11577 8495
rect 11615 8461 11649 8495
rect 11543 7380 11649 8422
rect 11820 8680 11854 8714
rect 11892 8680 11926 8714
rect 11820 8607 11854 8641
rect 11892 8607 11926 8641
rect 11820 8534 11854 8568
rect 11892 8534 11926 8568
rect 11820 8461 11854 8495
rect 11892 8461 11926 8495
rect 11820 7380 11926 8422
rect 12097 8680 12131 8714
rect 12169 8680 12203 8714
rect 12097 8607 12131 8641
rect 12169 8607 12203 8641
rect 12097 8534 12131 8568
rect 12169 8534 12203 8568
rect 12097 8461 12131 8495
rect 12169 8461 12203 8495
rect 12097 7380 12203 8422
rect 12374 8680 12408 8714
rect 12446 8680 12480 8714
rect 12374 8607 12408 8641
rect 12446 8607 12480 8641
rect 12374 8534 12408 8568
rect 12446 8534 12480 8568
rect 12374 8461 12408 8495
rect 12446 8461 12480 8495
rect 12374 7380 12480 8422
rect 12651 8680 12685 8714
rect 12723 8680 12757 8714
rect 12651 8607 12685 8641
rect 12723 8607 12757 8641
rect 12651 8534 12685 8568
rect 12723 8534 12757 8568
rect 12651 8461 12685 8495
rect 12723 8461 12757 8495
rect 12651 7380 12757 8422
rect 12928 8680 12962 8714
rect 13000 8680 13034 8714
rect 12928 8607 12962 8641
rect 13000 8607 13034 8641
rect 12928 8534 12962 8568
rect 13000 8534 13034 8568
rect 12928 8461 12962 8495
rect 13000 8461 13034 8495
rect 12928 7380 13034 8422
rect 13205 8680 13239 8714
rect 13277 8680 13311 8714
rect 13205 8607 13239 8641
rect 13277 8607 13311 8641
rect 13205 8534 13239 8568
rect 13277 8534 13311 8568
rect 13205 8461 13239 8495
rect 13277 8461 13311 8495
rect 13205 7380 13311 8422
rect 2638 7209 2672 7243
rect 2710 7209 2744 7243
rect 2638 7119 2672 7153
rect 2710 7119 2744 7153
rect 2638 7029 2672 7063
rect 2710 7029 2744 7063
rect 2638 6938 2672 6972
rect 2710 6938 2744 6972
rect 1944 6526 1946 6560
rect 1946 6526 1978 6560
rect 2016 6526 2048 6560
rect 2048 6526 2050 6560
rect 1944 6453 1946 6487
rect 1946 6453 1978 6487
rect 2016 6453 2048 6487
rect 2048 6453 2050 6487
rect 1944 6380 1946 6414
rect 1946 6380 1978 6414
rect 2016 6380 2048 6414
rect 2048 6380 2050 6414
rect 1944 6307 1946 6341
rect 1946 6307 1978 6341
rect 2016 6307 2048 6341
rect 2048 6307 2050 6341
rect 1944 6234 1946 6268
rect 1946 6234 1978 6268
rect 2016 6234 2048 6268
rect 2048 6234 2050 6268
rect 1944 6161 1946 6195
rect 1946 6161 1978 6195
rect 2016 6161 2048 6195
rect 2048 6161 2050 6195
rect 1944 6088 1946 6122
rect 1946 6088 1978 6122
rect 2016 6088 2048 6122
rect 2048 6088 2050 6122
rect 1944 6015 1946 6049
rect 1946 6015 1978 6049
rect 2016 6015 2048 6049
rect 2048 6015 2050 6049
rect 1944 5942 1946 5976
rect 1946 5942 1978 5976
rect 2016 5942 2048 5976
rect 2048 5942 2050 5976
rect 1944 5869 1946 5903
rect 1946 5869 1978 5903
rect 2016 5869 2048 5903
rect 2048 5869 2050 5903
rect 1944 5796 1946 5830
rect 1946 5796 1978 5830
rect 2016 5796 2048 5830
rect 2048 5796 2050 5830
rect 1944 5723 1946 5757
rect 1946 5723 1978 5757
rect 2016 5723 2048 5757
rect 2048 5723 2050 5757
rect 1944 5649 1946 5683
rect 1946 5649 1978 5683
rect 2016 5649 2048 5683
rect 2048 5649 2050 5683
rect 1944 5575 1946 5609
rect 1946 5575 1978 5609
rect 2016 5575 2048 5609
rect 2048 5575 2050 5609
rect 1944 5508 1946 5535
rect 1946 5508 1978 5535
rect 2016 5508 2048 5535
rect 2048 5508 2050 5535
rect 1944 5501 1978 5508
rect 2016 5501 2050 5508
rect 1944 5427 1978 5461
rect 2016 5427 2050 5461
rect 1944 5353 1978 5387
rect 2016 5353 2050 5387
rect 1944 5279 1946 5313
rect 1946 5279 1978 5313
rect 2016 5279 2048 5313
rect 2048 5279 2050 5313
rect 1944 5205 1946 5239
rect 1946 5205 1978 5239
rect 2016 5205 2048 5239
rect 2048 5205 2050 5239
rect 1944 5131 1946 5165
rect 1946 5131 1978 5165
rect 2016 5131 2048 5165
rect 2048 5131 2050 5165
rect 1944 5057 1946 5091
rect 1946 5057 1978 5091
rect 2016 5057 2048 5091
rect 2048 5057 2050 5091
rect 1944 4983 1946 5017
rect 1946 4983 1978 5017
rect 2016 4983 2048 5017
rect 2048 4983 2050 5017
rect 2255 6774 2274 6808
rect 2274 6774 2289 6808
rect 2327 6774 2361 6808
rect 2255 6701 2274 6735
rect 2274 6701 2289 6735
rect 2327 6701 2361 6735
rect 2255 6628 2274 6662
rect 2274 6628 2289 6662
rect 2327 6628 2361 6662
rect 2255 6555 2274 6589
rect 2274 6555 2289 6589
rect 2327 6555 2361 6589
rect 2255 6482 2274 6516
rect 2274 6482 2289 6516
rect 2327 6482 2361 6516
rect 2255 6409 2274 6443
rect 2274 6409 2289 6443
rect 2327 6409 2361 6443
rect 2255 6336 2274 6370
rect 2274 6336 2289 6370
rect 2327 6336 2361 6370
rect 2255 6263 2274 6297
rect 2274 6263 2289 6297
rect 2327 6263 2361 6297
rect 2255 6190 2274 6224
rect 2274 6190 2289 6224
rect 2327 6190 2361 6224
rect 2255 6117 2274 6151
rect 2274 6117 2289 6151
rect 2327 6117 2361 6151
rect 2255 6044 2274 6078
rect 2274 6044 2289 6078
rect 2327 6044 2361 6078
rect 2255 5971 2274 6005
rect 2274 5971 2289 6005
rect 2327 5971 2361 6005
rect 2255 5898 2274 5932
rect 2274 5898 2289 5932
rect 2327 5898 2361 5932
rect 2255 5825 2274 5859
rect 2274 5825 2289 5859
rect 2327 5825 2361 5859
rect 2255 5752 2274 5786
rect 2274 5752 2289 5786
rect 2327 5752 2361 5786
rect 2255 5679 2274 5713
rect 2274 5679 2289 5713
rect 2327 5679 2361 5713
rect 2255 5606 2274 5640
rect 2274 5606 2289 5640
rect 2327 5606 2361 5640
rect 2255 5533 2274 5567
rect 2274 5533 2289 5567
rect 2327 5533 2361 5567
rect 2255 5460 2274 5494
rect 2274 5460 2289 5494
rect 2327 5460 2361 5494
rect 2255 5387 2274 5421
rect 2274 5387 2289 5421
rect 2327 5387 2361 5421
rect 2679 6680 2713 6714
rect 2751 6680 2785 6714
rect 2679 6607 2713 6641
rect 2751 6607 2785 6641
rect 2679 6534 2713 6568
rect 2751 6534 2785 6568
rect 2679 6461 2713 6495
rect 2751 6461 2785 6495
rect 2679 5380 2785 6422
rect 2956 6680 2990 6714
rect 3028 6680 3062 6714
rect 2956 6607 2990 6641
rect 3028 6607 3062 6641
rect 2956 6534 2990 6568
rect 3028 6534 3062 6568
rect 2956 6461 2990 6495
rect 3028 6461 3062 6495
rect 2956 5380 3062 6422
rect 3233 6680 3267 6714
rect 3305 6680 3339 6714
rect 3233 6607 3267 6641
rect 3305 6607 3339 6641
rect 3233 6534 3267 6568
rect 3305 6534 3339 6568
rect 3233 6461 3267 6495
rect 3305 6461 3339 6495
rect 3233 5380 3339 6422
rect 3510 6680 3544 6714
rect 3582 6680 3616 6714
rect 3510 6607 3544 6641
rect 3582 6607 3616 6641
rect 3510 6534 3544 6568
rect 3582 6534 3616 6568
rect 3510 6461 3544 6495
rect 3582 6461 3616 6495
rect 3510 5380 3616 6422
rect 3787 6680 3821 6714
rect 3859 6680 3893 6714
rect 3787 6607 3821 6641
rect 3859 6607 3893 6641
rect 3787 6534 3821 6568
rect 3859 6534 3893 6568
rect 3787 6461 3821 6495
rect 3859 6461 3893 6495
rect 3787 5380 3893 6422
rect 4064 6680 4098 6714
rect 4136 6680 4170 6714
rect 4064 6607 4098 6641
rect 4136 6607 4170 6641
rect 4064 6534 4098 6568
rect 4136 6534 4170 6568
rect 4064 6461 4098 6495
rect 4136 6461 4170 6495
rect 4064 5380 4170 6422
rect 4341 6680 4375 6714
rect 4413 6680 4447 6714
rect 4341 6607 4375 6641
rect 4413 6607 4447 6641
rect 4341 6534 4375 6568
rect 4413 6534 4447 6568
rect 4341 6461 4375 6495
rect 4413 6461 4447 6495
rect 4341 5380 4447 6422
rect 4618 6680 4652 6714
rect 4690 6680 4724 6714
rect 4618 6607 4652 6641
rect 4690 6607 4724 6641
rect 4618 6534 4652 6568
rect 4690 6534 4724 6568
rect 4618 6461 4652 6495
rect 4690 6461 4724 6495
rect 4618 5380 4724 6422
rect 4895 6680 4929 6714
rect 4967 6680 5001 6714
rect 4895 6607 4929 6641
rect 4967 6607 5001 6641
rect 4895 6534 4929 6568
rect 4967 6534 5001 6568
rect 4895 6461 4929 6495
rect 4967 6461 5001 6495
rect 4895 5380 5001 6422
rect 5172 6680 5206 6714
rect 5244 6680 5278 6714
rect 5172 6607 5206 6641
rect 5244 6607 5278 6641
rect 5172 6534 5206 6568
rect 5244 6534 5278 6568
rect 5172 6461 5206 6495
rect 5244 6461 5278 6495
rect 5172 5380 5278 6422
rect 5449 6680 5483 6714
rect 5521 6680 5555 6714
rect 5449 6607 5483 6641
rect 5521 6607 5555 6641
rect 5449 6534 5483 6568
rect 5521 6534 5555 6568
rect 5449 6461 5483 6495
rect 5521 6461 5555 6495
rect 5449 5380 5555 6422
rect 5726 6680 5760 6714
rect 5798 6680 5832 6714
rect 5726 6607 5760 6641
rect 5798 6607 5832 6641
rect 5726 6534 5760 6568
rect 5798 6534 5832 6568
rect 5726 6461 5760 6495
rect 5798 6461 5832 6495
rect 5726 5380 5832 6422
rect 6003 6680 6037 6714
rect 6075 6680 6109 6714
rect 6003 6607 6037 6641
rect 6075 6607 6109 6641
rect 6003 6534 6037 6568
rect 6075 6534 6109 6568
rect 6003 6461 6037 6495
rect 6075 6461 6109 6495
rect 6003 5380 6109 6422
rect 6280 6680 6314 6714
rect 6352 6680 6386 6714
rect 6280 6607 6314 6641
rect 6352 6607 6386 6641
rect 6280 6534 6314 6568
rect 6352 6534 6386 6568
rect 6280 6461 6314 6495
rect 6352 6461 6386 6495
rect 6280 5380 6386 6422
rect 6557 6680 6591 6714
rect 6629 6680 6663 6714
rect 6557 6607 6591 6641
rect 6629 6607 6663 6641
rect 6557 6534 6591 6568
rect 6629 6534 6663 6568
rect 6557 6461 6591 6495
rect 6629 6461 6663 6495
rect 6557 5380 6663 6422
rect 6834 6680 6868 6714
rect 6906 6680 6940 6714
rect 6834 6607 6868 6641
rect 6906 6607 6940 6641
rect 6834 6534 6868 6568
rect 6906 6534 6940 6568
rect 6834 6461 6868 6495
rect 6906 6461 6940 6495
rect 6834 5380 6940 6422
rect 7111 6680 7145 6714
rect 7183 6680 7217 6714
rect 7111 6607 7145 6641
rect 7183 6607 7217 6641
rect 7111 6534 7145 6568
rect 7183 6534 7217 6568
rect 7111 6461 7145 6495
rect 7183 6461 7217 6495
rect 7111 5380 7217 6422
rect 7388 6680 7422 6714
rect 7460 6680 7494 6714
rect 7388 6607 7422 6641
rect 7460 6607 7494 6641
rect 7388 6534 7422 6568
rect 7460 6534 7494 6568
rect 7388 6461 7422 6495
rect 7460 6461 7494 6495
rect 7388 5380 7494 6422
rect 7665 6680 7699 6714
rect 7737 6680 7771 6714
rect 7665 6607 7699 6641
rect 7737 6607 7771 6641
rect 7665 6534 7699 6568
rect 7737 6534 7771 6568
rect 7665 6461 7699 6495
rect 7737 6461 7771 6495
rect 7665 5380 7771 6422
rect 7942 6680 7976 6714
rect 8014 6680 8048 6714
rect 7942 6607 7976 6641
rect 8014 6607 8048 6641
rect 7942 6534 7976 6568
rect 8014 6534 8048 6568
rect 7942 6461 7976 6495
rect 8014 6461 8048 6495
rect 7942 5380 8048 6422
rect 8219 6680 8253 6714
rect 8291 6680 8325 6714
rect 8219 6607 8253 6641
rect 8291 6607 8325 6641
rect 8219 6534 8253 6568
rect 8291 6534 8325 6568
rect 8219 6461 8253 6495
rect 8291 6461 8325 6495
rect 8219 5380 8325 6422
rect 8496 6680 8530 6714
rect 8568 6680 8602 6714
rect 8496 6607 8530 6641
rect 8568 6607 8602 6641
rect 8496 6534 8530 6568
rect 8568 6534 8602 6568
rect 8496 6461 8530 6495
rect 8568 6461 8602 6495
rect 8496 5380 8602 6422
rect 8773 6680 8807 6714
rect 8845 6680 8879 6714
rect 8773 6607 8807 6641
rect 8845 6607 8879 6641
rect 8773 6534 8807 6568
rect 8845 6534 8879 6568
rect 8773 6461 8807 6495
rect 8845 6461 8879 6495
rect 8773 5380 8879 6422
rect 9050 6680 9084 6714
rect 9122 6680 9156 6714
rect 9050 6607 9084 6641
rect 9122 6607 9156 6641
rect 9050 6534 9084 6568
rect 9122 6534 9156 6568
rect 9050 6461 9084 6495
rect 9122 6461 9156 6495
rect 9050 5380 9156 6422
rect 9327 6680 9361 6714
rect 9399 6680 9433 6714
rect 9327 6607 9361 6641
rect 9399 6607 9433 6641
rect 9327 6534 9361 6568
rect 9399 6534 9433 6568
rect 9327 6461 9361 6495
rect 9399 6461 9433 6495
rect 9327 5380 9433 6422
rect 9604 6680 9638 6714
rect 9676 6680 9710 6714
rect 9604 6607 9638 6641
rect 9676 6607 9710 6641
rect 9604 6534 9638 6568
rect 9676 6534 9710 6568
rect 9604 6461 9638 6495
rect 9676 6461 9710 6495
rect 9604 5380 9710 6422
rect 9881 6680 9915 6714
rect 9953 6680 9987 6714
rect 9881 6607 9915 6641
rect 9953 6607 9987 6641
rect 9881 6534 9915 6568
rect 9953 6534 9987 6568
rect 9881 6461 9915 6495
rect 9953 6461 9987 6495
rect 9881 5380 9987 6422
rect 10158 6680 10192 6714
rect 10230 6680 10264 6714
rect 10158 6607 10192 6641
rect 10230 6607 10264 6641
rect 10158 6534 10192 6568
rect 10230 6534 10264 6568
rect 10158 6461 10192 6495
rect 10230 6461 10264 6495
rect 10158 5380 10264 6422
rect 10435 6680 10469 6714
rect 10507 6680 10541 6714
rect 10435 6607 10469 6641
rect 10507 6607 10541 6641
rect 10435 6534 10469 6568
rect 10507 6534 10541 6568
rect 10435 6461 10469 6495
rect 10507 6461 10541 6495
rect 10435 5380 10541 6422
rect 10712 6680 10746 6714
rect 10784 6680 10818 6714
rect 10712 6607 10746 6641
rect 10784 6607 10818 6641
rect 10712 6534 10746 6568
rect 10784 6534 10818 6568
rect 10712 6461 10746 6495
rect 10784 6461 10818 6495
rect 10712 5380 10818 6422
rect 10989 6680 11023 6714
rect 11061 6680 11095 6714
rect 10989 6607 11023 6641
rect 11061 6607 11095 6641
rect 10989 6534 11023 6568
rect 11061 6534 11095 6568
rect 10989 6461 11023 6495
rect 11061 6461 11095 6495
rect 10989 5380 11095 6422
rect 11266 6680 11300 6714
rect 11338 6680 11372 6714
rect 11266 6607 11300 6641
rect 11338 6607 11372 6641
rect 11266 6534 11300 6568
rect 11338 6534 11372 6568
rect 11266 6461 11300 6495
rect 11338 6461 11372 6495
rect 11266 5380 11372 6422
rect 11543 6680 11577 6714
rect 11615 6680 11649 6714
rect 11543 6607 11577 6641
rect 11615 6607 11649 6641
rect 11543 6534 11577 6568
rect 11615 6534 11649 6568
rect 11543 6461 11577 6495
rect 11615 6461 11649 6495
rect 11543 5380 11649 6422
rect 11820 6680 11854 6714
rect 11892 6680 11926 6714
rect 11820 6607 11854 6641
rect 11892 6607 11926 6641
rect 11820 6534 11854 6568
rect 11892 6534 11926 6568
rect 11820 6461 11854 6495
rect 11892 6461 11926 6495
rect 11820 5380 11926 6422
rect 12097 6680 12131 6714
rect 12169 6680 12203 6714
rect 12097 6607 12131 6641
rect 12169 6607 12203 6641
rect 12097 6534 12131 6568
rect 12169 6534 12203 6568
rect 12097 6461 12131 6495
rect 12169 6461 12203 6495
rect 12097 5380 12203 6422
rect 12374 6680 12408 6714
rect 12446 6680 12480 6714
rect 12374 6607 12408 6641
rect 12446 6607 12480 6641
rect 12374 6534 12408 6568
rect 12446 6534 12480 6568
rect 12374 6461 12408 6495
rect 12446 6461 12480 6495
rect 12374 5380 12480 6422
rect 12651 6680 12685 6714
rect 12723 6680 12757 6714
rect 12651 6607 12685 6641
rect 12723 6607 12757 6641
rect 12651 6534 12685 6568
rect 12723 6534 12757 6568
rect 12651 6461 12685 6495
rect 12723 6461 12757 6495
rect 12651 5380 12757 6422
rect 12928 6680 12962 6714
rect 13000 6680 13034 6714
rect 12928 6607 12962 6641
rect 13000 6607 13034 6641
rect 12928 6534 12962 6568
rect 13000 6534 13034 6568
rect 12928 6461 12962 6495
rect 13000 6461 13034 6495
rect 12928 5380 13034 6422
rect 13205 6680 13239 6714
rect 13277 6680 13311 6714
rect 13205 6607 13239 6641
rect 13277 6607 13311 6641
rect 13205 6534 13239 6568
rect 13277 6534 13311 6568
rect 13205 6461 13239 6495
rect 13277 6461 13311 6495
rect 13205 5380 13311 6422
rect 13490 5815 13596 19701
rect 13490 5742 13524 5776
rect 13562 5742 13596 5776
rect 13490 5669 13524 5703
rect 13562 5669 13596 5703
rect 13490 5596 13524 5630
rect 13562 5596 13596 5630
rect 13490 5523 13524 5557
rect 13562 5523 13596 5557
rect 13490 5450 13524 5484
rect 13562 5450 13596 5484
rect 13490 5377 13524 5411
rect 13562 5377 13596 5411
rect 2255 5314 2274 5348
rect 2274 5314 2289 5348
rect 2327 5314 2361 5348
rect 2255 5240 2274 5274
rect 2274 5240 2289 5274
rect 2327 5240 2361 5274
rect 13490 5304 13524 5338
rect 13562 5304 13596 5338
rect 13490 5231 13524 5265
rect 13562 5231 13596 5265
rect 2287 5163 2321 5197
rect 2360 5163 2394 5197
rect 2433 5183 2444 5197
rect 2444 5183 2467 5197
rect 2506 5183 2540 5197
rect 2579 5183 2613 5197
rect 2652 5183 2686 5197
rect 2725 5183 2759 5197
rect 2798 5183 2832 5197
rect 2871 5183 2905 5197
rect 2944 5183 2978 5197
rect 3017 5183 3051 5197
rect 3090 5183 3124 5197
rect 3163 5183 3197 5197
rect 3236 5183 3270 5197
rect 3309 5183 3343 5197
rect 3382 5183 3416 5197
rect 3455 5183 3489 5197
rect 3528 5183 3562 5197
rect 3601 5183 3635 5197
rect 3674 5183 3708 5197
rect 3747 5183 3781 5197
rect 3820 5183 3854 5197
rect 3893 5183 3927 5197
rect 3966 5183 4000 5197
rect 4039 5183 4073 5197
rect 4112 5183 4146 5197
rect 4185 5183 4219 5197
rect 4258 5183 4292 5197
rect 4331 5183 4365 5197
rect 4404 5183 4438 5197
rect 4477 5183 4511 5197
rect 4550 5183 4584 5197
rect 4623 5183 4657 5197
rect 4696 5183 4730 5197
rect 4769 5183 4803 5197
rect 4842 5183 4876 5197
rect 4915 5183 4949 5197
rect 4988 5183 5022 5197
rect 5061 5183 5095 5197
rect 5134 5183 5168 5197
rect 5207 5183 5241 5197
rect 5280 5183 5314 5197
rect 5353 5183 5387 5197
rect 5426 5183 13452 5197
rect 2433 5163 2467 5183
rect 2506 5163 2540 5183
rect 2579 5163 2613 5183
rect 2652 5163 2686 5183
rect 2725 5163 2759 5183
rect 2798 5163 2832 5183
rect 2871 5163 2905 5183
rect 2944 5163 2978 5183
rect 3017 5163 3051 5183
rect 3090 5163 3124 5183
rect 3163 5163 3197 5183
rect 3236 5163 3270 5183
rect 3309 5163 3343 5183
rect 3382 5163 3416 5183
rect 3455 5163 3489 5183
rect 3528 5163 3562 5183
rect 3601 5163 3635 5183
rect 3674 5163 3708 5183
rect 3747 5163 3781 5183
rect 3820 5163 3854 5183
rect 3893 5163 3927 5183
rect 3966 5163 4000 5183
rect 4039 5163 4073 5183
rect 4112 5163 4146 5183
rect 4185 5163 4219 5183
rect 4258 5163 4292 5183
rect 4331 5163 4365 5183
rect 4404 5163 4438 5183
rect 4477 5163 4511 5183
rect 4550 5163 4584 5183
rect 4623 5163 4657 5183
rect 4696 5163 4730 5183
rect 4769 5163 4803 5183
rect 4842 5163 4876 5183
rect 4915 5163 4949 5183
rect 4988 5163 5022 5183
rect 5061 5163 5095 5183
rect 5134 5163 5168 5183
rect 5207 5163 5241 5183
rect 5280 5163 5314 5183
rect 5353 5163 5387 5183
rect 2287 5091 2321 5125
rect 2360 5091 2394 5125
rect 2433 5091 2467 5125
rect 2506 5091 2540 5125
rect 2579 5091 2613 5125
rect 2652 5091 2686 5125
rect 2725 5091 2759 5125
rect 2798 5091 2832 5125
rect 2871 5091 2905 5125
rect 2944 5091 2978 5125
rect 3017 5091 3051 5125
rect 3090 5091 3124 5125
rect 3163 5091 3197 5125
rect 3236 5091 3270 5125
rect 3309 5091 3343 5125
rect 3382 5091 3416 5125
rect 3455 5091 3489 5125
rect 3528 5091 3562 5125
rect 3601 5091 3635 5125
rect 3674 5091 3708 5125
rect 3747 5091 3781 5125
rect 3820 5091 3854 5125
rect 3893 5091 3927 5125
rect 3966 5091 4000 5125
rect 4039 5091 4073 5125
rect 4112 5091 4146 5125
rect 4185 5091 4219 5125
rect 4258 5091 4292 5125
rect 4331 5091 4365 5125
rect 4404 5091 4438 5125
rect 4477 5091 4511 5125
rect 4550 5091 4584 5125
rect 4623 5091 4657 5125
rect 4696 5091 4730 5125
rect 4769 5091 4803 5125
rect 4842 5091 4876 5125
rect 4915 5091 4949 5125
rect 4988 5091 5022 5125
rect 5061 5091 5095 5125
rect 5134 5091 5168 5125
rect 5207 5091 5241 5125
rect 5280 5091 5314 5125
rect 5353 5091 5387 5125
rect 5426 5081 13392 5183
rect 13392 5081 13452 5183
rect 13490 5158 13524 5192
rect 13562 5158 13596 5192
rect 13490 5115 13524 5119
rect 13562 5115 13596 5119
rect 13490 5085 13524 5115
rect 13562 5085 13596 5115
rect 2287 5019 2321 5053
rect 2360 5019 2394 5053
rect 2433 5019 2467 5053
rect 2506 5019 2540 5053
rect 2579 5019 2613 5053
rect 2652 5019 2686 5053
rect 2725 5019 2759 5053
rect 2798 5019 2832 5053
rect 2871 5019 2905 5053
rect 2944 5019 2978 5053
rect 3017 5019 3051 5053
rect 3090 5019 3124 5053
rect 3163 5019 3197 5053
rect 3236 5019 3270 5053
rect 3309 5019 3343 5053
rect 3382 5019 3416 5053
rect 3455 5019 3489 5053
rect 3528 5019 3562 5053
rect 3601 5019 3635 5053
rect 3674 5019 3708 5053
rect 3747 5019 3781 5053
rect 3820 5019 3854 5053
rect 3893 5019 3927 5053
rect 3966 5019 4000 5053
rect 4039 5019 4073 5053
rect 4112 5019 4146 5053
rect 4185 5019 4219 5053
rect 4258 5019 4292 5053
rect 4331 5019 4365 5053
rect 4404 5019 4438 5053
rect 4477 5019 4511 5053
rect 4550 5019 4584 5053
rect 4623 5019 4657 5053
rect 4696 5019 4730 5053
rect 4769 5019 4803 5053
rect 4842 5019 4876 5053
rect 4915 5019 4949 5053
rect 4988 5019 5022 5053
rect 5061 5019 5095 5053
rect 5134 5019 5168 5053
rect 5207 5019 5241 5053
rect 5280 5019 5314 5053
rect 5353 5019 5387 5053
rect 5426 5019 13452 5081
rect 13838 6895 13840 21329
rect 13840 6895 13942 21329
rect 13942 6895 13944 21329
rect 13838 6822 13840 6856
rect 13840 6822 13872 6856
rect 13910 6822 13942 6856
rect 13942 6822 13944 6856
rect 13838 6749 13840 6783
rect 13840 6749 13872 6783
rect 13910 6749 13942 6783
rect 13942 6749 13944 6783
rect 13838 6676 13840 6710
rect 13840 6676 13872 6710
rect 13910 6676 13942 6710
rect 13942 6676 13944 6710
rect 13838 6603 13840 6637
rect 13840 6603 13872 6637
rect 13910 6603 13942 6637
rect 13942 6603 13944 6637
rect 13838 6530 13840 6564
rect 13840 6530 13872 6564
rect 13910 6530 13942 6564
rect 13942 6530 13944 6564
rect 13838 6457 13840 6491
rect 13840 6457 13872 6491
rect 13910 6457 13942 6491
rect 13942 6457 13944 6491
rect 13838 6384 13840 6418
rect 13840 6384 13872 6418
rect 13910 6384 13942 6418
rect 13942 6384 13944 6418
rect 13838 6311 13840 6345
rect 13840 6311 13872 6345
rect 13910 6311 13942 6345
rect 13942 6311 13944 6345
rect 13838 6238 13840 6272
rect 13840 6238 13872 6272
rect 13910 6238 13942 6272
rect 13942 6238 13944 6272
rect 13838 6165 13840 6199
rect 13840 6165 13872 6199
rect 13910 6165 13942 6199
rect 13942 6165 13944 6199
rect 13838 6092 13840 6126
rect 13840 6092 13872 6126
rect 13910 6092 13942 6126
rect 13942 6092 13944 6126
rect 13838 6019 13840 6053
rect 13840 6019 13872 6053
rect 13910 6019 13942 6053
rect 13942 6019 13944 6053
rect 13838 5946 13840 5980
rect 13840 5946 13872 5980
rect 13910 5946 13942 5980
rect 13942 5946 13944 5980
rect 13838 5873 13840 5907
rect 13840 5873 13872 5907
rect 13910 5873 13942 5907
rect 13942 5873 13944 5907
rect 13838 5800 13840 5834
rect 13840 5800 13872 5834
rect 13910 5800 13942 5834
rect 13942 5800 13944 5834
rect 13838 5727 13840 5761
rect 13840 5727 13872 5761
rect 13910 5727 13942 5761
rect 13942 5727 13944 5761
rect 13838 5654 13840 5688
rect 13840 5654 13872 5688
rect 13910 5654 13942 5688
rect 13942 5654 13944 5688
rect 13838 5593 13840 5615
rect 13840 5593 13872 5615
rect 13910 5593 13942 5615
rect 13942 5593 13944 5615
rect 13838 5581 13872 5593
rect 13910 5581 13944 5593
rect 13838 5508 13872 5542
rect 13910 5508 13944 5542
rect 13838 5435 13840 5469
rect 13840 5435 13872 5469
rect 13910 5435 13942 5469
rect 13942 5435 13944 5469
rect 13838 5362 13840 5396
rect 13840 5362 13872 5396
rect 13910 5362 13942 5396
rect 13942 5362 13944 5396
rect 13838 5289 13840 5323
rect 13840 5289 13872 5323
rect 13910 5289 13942 5323
rect 13942 5289 13944 5323
rect 13838 5216 13840 5250
rect 13840 5216 13872 5250
rect 13910 5216 13942 5250
rect 13942 5216 13944 5250
rect 13838 5143 13840 5177
rect 13840 5143 13872 5177
rect 13910 5143 13942 5177
rect 13942 5143 13944 5177
rect 13838 5070 13840 5104
rect 13840 5070 13872 5104
rect 13910 5070 13942 5104
rect 13942 5070 13944 5104
rect 1944 4909 1946 4943
rect 1946 4909 1978 4943
rect 2016 4909 2048 4943
rect 2048 4909 2050 4943
rect 13838 4997 13840 5031
rect 13840 4997 13872 5031
rect 13910 4997 13942 5031
rect 13942 4997 13944 5031
rect 13838 4924 13840 4958
rect 13840 4924 13872 4958
rect 13910 4924 13942 4958
rect 13942 4924 13944 4958
rect 1950 4837 1984 4871
rect 2023 4837 2048 4871
rect 2048 4837 2057 4871
rect 2096 4869 2130 4871
rect 2169 4869 2203 4871
rect 2242 4869 2276 4871
rect 2315 4869 2349 4871
rect 2388 4869 2422 4871
rect 2461 4869 2495 4871
rect 2534 4869 2568 4871
rect 2096 4837 2130 4869
rect 2169 4837 2203 4869
rect 2242 4837 2276 4869
rect 2315 4837 2349 4869
rect 2388 4837 2422 4869
rect 2461 4837 2495 4869
rect 2534 4837 2568 4869
rect 2607 4837 2641 4871
rect 2680 4869 2714 4871
rect 2753 4869 2787 4871
rect 2826 4869 2860 4871
rect 2899 4869 2933 4871
rect 2972 4869 3006 4871
rect 3045 4869 3079 4871
rect 3118 4869 3152 4871
rect 3191 4869 3225 4871
rect 3264 4869 3298 4871
rect 3337 4869 3371 4871
rect 3410 4869 3444 4871
rect 3483 4869 3517 4871
rect 3556 4869 3590 4871
rect 3629 4869 3663 4871
rect 3702 4869 3736 4871
rect 3775 4869 3809 4871
rect 3848 4869 3882 4871
rect 3921 4869 3955 4871
rect 3994 4869 4028 4871
rect 4067 4869 4101 4871
rect 4140 4869 4174 4871
rect 4213 4869 4247 4871
rect 4286 4869 4320 4871
rect 4359 4869 4393 4871
rect 4432 4869 4466 4871
rect 4505 4869 4539 4871
rect 4578 4869 4612 4871
rect 4651 4869 4685 4871
rect 4724 4869 4758 4871
rect 4797 4869 4831 4871
rect 4870 4869 4904 4871
rect 4943 4869 4977 4871
rect 5016 4869 5050 4871
rect 5089 4869 5123 4871
rect 5162 4869 5196 4871
rect 5235 4869 13765 4871
rect 2680 4837 2714 4869
rect 2753 4837 2787 4869
rect 2826 4837 2860 4869
rect 2899 4837 2933 4869
rect 2972 4837 3006 4869
rect 3045 4837 3079 4869
rect 3118 4837 3152 4869
rect 3191 4837 3225 4869
rect 3264 4837 3298 4869
rect 3337 4837 3371 4869
rect 3410 4837 3444 4869
rect 3483 4837 3517 4869
rect 3556 4837 3590 4869
rect 3629 4837 3663 4869
rect 3702 4837 3736 4869
rect 3775 4837 3809 4869
rect 3848 4837 3882 4869
rect 3921 4837 3955 4869
rect 3994 4837 4028 4869
rect 4067 4837 4101 4869
rect 4140 4837 4174 4869
rect 4213 4837 4247 4869
rect 4286 4837 4320 4869
rect 4359 4837 4393 4869
rect 4432 4837 4466 4869
rect 4505 4837 4539 4869
rect 4578 4837 4612 4869
rect 4651 4837 4685 4869
rect 4724 4837 4758 4869
rect 4797 4837 4831 4869
rect 4870 4837 4904 4869
rect 4943 4837 4977 4869
rect 5016 4837 5050 4869
rect 5089 4837 5123 4869
rect 5162 4837 5196 4869
rect 1950 4765 1984 4799
rect 2023 4767 2054 4799
rect 2054 4767 2057 4799
rect 2096 4767 2130 4799
rect 2169 4767 2203 4799
rect 2242 4767 2276 4799
rect 2315 4767 2349 4799
rect 2388 4767 2422 4799
rect 2461 4767 2495 4799
rect 2534 4767 2568 4799
rect 2023 4765 2057 4767
rect 2096 4765 2130 4767
rect 2169 4765 2203 4767
rect 2242 4765 2276 4767
rect 2315 4765 2349 4767
rect 2388 4765 2422 4767
rect 2461 4765 2495 4767
rect 2534 4765 2568 4767
rect 2607 4765 2641 4799
rect 2680 4767 2714 4799
rect 2753 4767 2787 4799
rect 2826 4767 2860 4799
rect 2899 4767 2933 4799
rect 2972 4767 3006 4799
rect 3045 4767 3079 4799
rect 3118 4767 3152 4799
rect 3191 4767 3225 4799
rect 3264 4767 3298 4799
rect 3337 4767 3371 4799
rect 3410 4767 3444 4799
rect 3483 4767 3517 4799
rect 3556 4767 3590 4799
rect 3629 4767 3663 4799
rect 3702 4767 3736 4799
rect 3775 4767 3809 4799
rect 3848 4767 3882 4799
rect 3921 4767 3955 4799
rect 3994 4767 4028 4799
rect 4067 4767 4101 4799
rect 4140 4767 4174 4799
rect 4213 4767 4247 4799
rect 4286 4767 4320 4799
rect 4359 4767 4393 4799
rect 4432 4767 4466 4799
rect 4505 4767 4539 4799
rect 4578 4767 4612 4799
rect 4651 4767 4685 4799
rect 4724 4767 4758 4799
rect 4797 4767 4831 4799
rect 4870 4767 4904 4799
rect 4943 4767 4977 4799
rect 5016 4767 5050 4799
rect 5089 4767 5123 4799
rect 5162 4767 5196 4799
rect 5235 4767 13240 4869
rect 13240 4767 13340 4869
rect 13340 4767 13765 4869
rect 13838 4851 13840 4885
rect 13840 4851 13872 4885
rect 13910 4851 13942 4885
rect 13942 4851 13944 4885
rect 13838 4801 13872 4812
rect 13838 4778 13850 4801
rect 13850 4778 13872 4801
rect 13910 4778 13944 4812
rect 2680 4765 2714 4767
rect 2753 4765 2787 4767
rect 2826 4765 2860 4767
rect 2899 4765 2933 4767
rect 2972 4765 3006 4767
rect 3045 4765 3079 4767
rect 3118 4765 3152 4767
rect 3191 4765 3225 4767
rect 3264 4765 3298 4767
rect 3337 4765 3371 4767
rect 3410 4765 3444 4767
rect 3483 4765 3517 4767
rect 3556 4765 3590 4767
rect 3629 4765 3663 4767
rect 3702 4765 3736 4767
rect 3775 4765 3809 4767
rect 3848 4765 3882 4767
rect 3921 4765 3955 4767
rect 3994 4765 4028 4767
rect 4067 4765 4101 4767
rect 4140 4765 4174 4767
rect 4213 4765 4247 4767
rect 4286 4765 4320 4767
rect 4359 4765 4393 4767
rect 4432 4765 4466 4767
rect 4505 4765 4539 4767
rect 4578 4765 4612 4767
rect 4651 4765 4685 4767
rect 4724 4765 4758 4767
rect 4797 4765 4831 4767
rect 4870 4765 4904 4767
rect 4943 4765 4977 4767
rect 5016 4765 5050 4767
rect 5089 4765 5123 4767
rect 5162 4765 5196 4767
rect 5235 4765 13765 4767
rect 423 4572 457 4606
rect 423 4495 457 4529
rect 995 4568 1029 4602
rect 1099 4568 1133 4602
rect 1202 4568 1236 4602
rect 995 4458 1029 4492
rect 1099 4458 1133 4492
rect 1202 4458 1236 4492
rect 423 4418 457 4452
rect 423 4341 457 4375
rect 423 4264 457 4298
rect 423 4186 457 4220
rect 423 4108 457 4142
rect 1668 3950 1702 3984
rect 1753 3950 1787 3984
rect 1838 3950 1872 3984
rect 13906 3888 13940 3922
rect 14019 3888 14053 3922
rect 13906 3802 13940 3836
rect 14019 3802 14053 3836
rect 14099 3705 14133 3739
rect 14185 3705 14219 3739
rect 368 3555 402 3589
rect 467 3555 501 3589
rect 565 3555 599 3589
rect 368 3483 402 3517
rect 467 3483 501 3517
rect 565 3483 599 3517
rect 1749 3646 1783 3664
rect 1822 3646 1856 3664
rect 1895 3646 1929 3664
rect 1968 3646 2002 3664
rect 2041 3646 2075 3664
rect 2113 3646 2147 3664
rect 2185 3646 2219 3664
rect 2257 3646 2291 3664
rect 2329 3646 2363 3664
rect 2401 3646 2435 3664
rect 2473 3646 2507 3664
rect 2545 3646 2579 3664
rect 2617 3646 2651 3664
rect 2689 3646 2723 3664
rect 1749 3630 1781 3646
rect 1781 3630 1783 3646
rect 1822 3630 1851 3646
rect 1851 3630 1856 3646
rect 1895 3630 1921 3646
rect 1921 3630 1929 3646
rect 1968 3630 1991 3646
rect 1991 3630 2002 3646
rect 2041 3630 2061 3646
rect 2061 3630 2075 3646
rect 2113 3630 2131 3646
rect 2131 3630 2147 3646
rect 2185 3630 2201 3646
rect 2201 3630 2219 3646
rect 2257 3630 2271 3646
rect 2271 3630 2291 3646
rect 2329 3630 2341 3646
rect 2341 3630 2363 3646
rect 2401 3630 2411 3646
rect 2411 3630 2435 3646
rect 2473 3630 2481 3646
rect 2481 3630 2507 3646
rect 2545 3630 2551 3646
rect 2551 3630 2579 3646
rect 2617 3630 2621 3646
rect 2621 3630 2651 3646
rect 2689 3630 2691 3646
rect 2691 3630 2723 3646
rect 2761 3630 2795 3664
rect 2833 3630 2867 3664
rect 2905 3646 2939 3664
rect 2977 3646 3011 3664
rect 3049 3646 3083 3664
rect 3121 3646 3155 3664
rect 3193 3646 3227 3664
rect 3265 3646 3299 3664
rect 2905 3630 2937 3646
rect 2937 3630 2939 3646
rect 2977 3630 3007 3646
rect 3007 3630 3011 3646
rect 3049 3630 3077 3646
rect 3077 3630 3083 3646
rect 3121 3630 3147 3646
rect 3147 3630 3155 3646
rect 3193 3630 3217 3646
rect 3217 3630 3227 3646
rect 3265 3630 3287 3646
rect 3287 3630 3299 3646
rect 1677 3578 1711 3592
rect 1677 3558 1711 3578
rect 1785 3544 1817 3556
rect 1817 3544 1819 3556
rect 1859 3544 1887 3556
rect 1887 3544 1893 3556
rect 1933 3544 1957 3556
rect 1957 3544 1967 3556
rect 2007 3544 2027 3556
rect 2027 3544 2041 3556
rect 2081 3544 2097 3556
rect 2097 3544 2115 3556
rect 2155 3544 2167 3556
rect 2167 3544 2189 3556
rect 2229 3544 2237 3556
rect 2237 3544 2263 3556
rect 2303 3544 2307 3556
rect 2307 3544 2337 3556
rect 2377 3544 2411 3556
rect 2451 3544 2481 3556
rect 2481 3544 2485 3556
rect 2525 3544 2551 3556
rect 2551 3544 2559 3556
rect 2599 3544 2621 3556
rect 2621 3544 2633 3556
rect 2673 3544 2691 3556
rect 2691 3544 2707 3556
rect 2747 3544 2761 3556
rect 2761 3544 2781 3556
rect 2821 3544 2831 3556
rect 2831 3544 2855 3556
rect 2895 3544 2901 3556
rect 2901 3544 2929 3556
rect 2969 3544 2971 3556
rect 2971 3544 3003 3556
rect 1785 3522 1819 3544
rect 1859 3522 1893 3544
rect 1933 3522 1967 3544
rect 2007 3522 2041 3544
rect 2081 3522 2115 3544
rect 2155 3522 2189 3544
rect 2229 3522 2263 3544
rect 2303 3522 2337 3544
rect 2377 3522 2411 3544
rect 2451 3522 2485 3544
rect 2525 3522 2559 3544
rect 2599 3522 2633 3544
rect 2673 3522 2707 3544
rect 2747 3522 2781 3544
rect 2821 3522 2855 3544
rect 2895 3522 2929 3544
rect 2969 3522 3003 3544
rect 3043 3522 3077 3556
rect 3117 3544 3147 3556
rect 3147 3544 3151 3556
rect 3191 3544 3217 3556
rect 3217 3544 3225 3556
rect 3265 3544 3287 3556
rect 3287 3544 3299 3556
rect 3117 3522 3151 3544
rect 3191 3522 3225 3544
rect 3265 3522 3299 3544
rect 1677 3510 1711 3520
rect 3432 3630 3466 3664
rect 3505 3630 3539 3664
rect 3578 3630 3612 3664
rect 3651 3630 3685 3664
rect 3724 3630 3758 3664
rect 3797 3630 3831 3664
rect 3870 3630 3904 3664
rect 3942 3630 3976 3664
rect 4014 3630 4048 3664
rect 4086 3630 4120 3664
rect 4158 3630 4192 3664
rect 4230 3630 4264 3664
rect 4302 3630 4336 3664
rect 4374 3630 4408 3664
rect 4446 3630 4480 3664
rect 4518 3630 4552 3664
rect 4590 3630 4624 3664
rect 4662 3630 4696 3664
rect 4734 3630 4768 3664
rect 4806 3630 4840 3664
rect 4878 3630 4912 3664
rect 4950 3630 4984 3664
rect 5022 3630 5056 3664
rect 5094 3630 5128 3664
rect 5166 3630 5200 3664
rect 5238 3630 5272 3664
rect 5310 3630 5344 3664
rect 5382 3630 5416 3664
rect 5454 3630 5488 3664
rect 5526 3630 5560 3664
rect 5598 3630 5632 3664
rect 5670 3630 5704 3664
rect 5742 3630 5776 3664
rect 5814 3630 5848 3664
rect 5886 3630 5920 3664
rect 5958 3630 5992 3664
rect 6030 3630 6064 3664
rect 6102 3630 6136 3664
rect 6174 3630 6208 3664
rect 6246 3630 6280 3664
rect 6318 3630 6352 3664
rect 6390 3630 6424 3664
rect 6462 3630 6496 3664
rect 6534 3630 6568 3664
rect 6606 3630 6640 3664
rect 6678 3630 6712 3664
rect 6750 3630 6784 3664
rect 6822 3630 6856 3664
rect 6894 3630 6928 3664
rect 6966 3630 7000 3664
rect 7038 3630 7072 3664
rect 7110 3630 7144 3664
rect 7182 3630 7216 3664
rect 7428 3630 7462 3664
rect 7501 3630 7535 3664
rect 7574 3630 7608 3664
rect 7646 3630 7680 3664
rect 7718 3630 7752 3664
rect 7790 3630 7824 3664
rect 7862 3630 7896 3664
rect 7934 3630 7968 3664
rect 8006 3630 8040 3664
rect 8078 3630 8112 3664
rect 8150 3630 8184 3664
rect 8222 3630 8256 3664
rect 8294 3630 8328 3664
rect 8366 3630 8400 3664
rect 8438 3630 8472 3664
rect 8510 3630 8544 3664
rect 8582 3630 8616 3664
rect 8654 3630 8688 3664
rect 8726 3630 8760 3664
rect 8798 3630 8832 3664
rect 8870 3630 8904 3664
rect 8942 3630 8976 3664
rect 9014 3630 9048 3664
rect 9086 3630 9120 3664
rect 9158 3630 9192 3664
rect 9230 3630 9264 3664
rect 9302 3630 9336 3664
rect 9374 3630 9408 3664
rect 9446 3630 9480 3664
rect 9518 3630 9552 3664
rect 9590 3630 9624 3664
rect 9662 3630 9696 3664
rect 9734 3630 9768 3664
rect 9806 3630 9840 3664
rect 9878 3630 9912 3664
rect 9950 3630 9984 3664
rect 10022 3630 10056 3664
rect 10094 3630 10128 3664
rect 10166 3630 10200 3664
rect 10238 3630 10272 3664
rect 10310 3630 10344 3664
rect 10382 3630 10416 3664
rect 10454 3630 10488 3664
rect 10526 3630 10560 3664
rect 10598 3630 10632 3664
rect 10670 3630 10704 3664
rect 10742 3630 10776 3664
rect 10814 3630 10848 3664
rect 10886 3630 10920 3664
rect 10958 3630 10992 3664
rect 11030 3630 11064 3664
rect 11102 3630 11136 3664
rect 11174 3630 11208 3664
rect 14099 3592 14133 3626
rect 14185 3592 14219 3626
rect 3432 3522 3466 3556
rect 3505 3522 3539 3556
rect 3578 3522 3612 3556
rect 3651 3522 3685 3556
rect 3724 3522 3758 3556
rect 3797 3522 3831 3556
rect 3870 3522 3904 3556
rect 3942 3522 3976 3556
rect 4014 3522 4048 3556
rect 4086 3522 4120 3556
rect 4158 3522 4192 3556
rect 4230 3522 4264 3556
rect 4302 3522 4336 3556
rect 4374 3522 4408 3556
rect 4446 3522 4480 3556
rect 4518 3522 4552 3556
rect 4590 3522 4624 3556
rect 4662 3522 4696 3556
rect 4734 3522 4768 3556
rect 4806 3522 4840 3556
rect 4878 3522 4912 3556
rect 4950 3522 4984 3556
rect 5022 3522 5056 3556
rect 5094 3522 5128 3556
rect 5166 3522 5200 3556
rect 5238 3522 5272 3556
rect 5310 3522 5344 3556
rect 5382 3522 5416 3556
rect 5454 3522 5488 3556
rect 5526 3522 5560 3556
rect 5598 3522 5632 3556
rect 5670 3522 5704 3556
rect 5742 3522 5776 3556
rect 5814 3522 5848 3556
rect 5886 3522 5920 3556
rect 5958 3522 5992 3556
rect 6030 3522 6064 3556
rect 6102 3522 6136 3556
rect 6174 3522 6208 3556
rect 6246 3522 6280 3556
rect 6318 3522 6352 3556
rect 6390 3522 6424 3556
rect 6462 3522 6496 3556
rect 6534 3522 6568 3556
rect 6606 3522 6640 3556
rect 6678 3522 6712 3556
rect 6750 3522 6784 3556
rect 6822 3522 6856 3556
rect 6894 3522 6928 3556
rect 6966 3522 7000 3556
rect 7038 3522 7072 3556
rect 7110 3522 7144 3556
rect 7182 3522 7216 3556
rect 7428 3522 7462 3556
rect 7501 3522 7535 3556
rect 7574 3522 7608 3556
rect 7646 3522 7680 3556
rect 7718 3522 7752 3556
rect 7790 3522 7824 3556
rect 7862 3522 7896 3556
rect 7934 3522 7968 3556
rect 8006 3522 8040 3556
rect 8078 3522 8112 3556
rect 8150 3522 8184 3556
rect 8222 3522 8256 3556
rect 8294 3522 8328 3556
rect 8366 3522 8400 3556
rect 8438 3522 8472 3556
rect 8510 3522 8544 3556
rect 8582 3522 8616 3556
rect 8654 3522 8688 3556
rect 8726 3522 8760 3556
rect 8798 3522 8832 3556
rect 8870 3522 8904 3556
rect 8942 3522 8976 3556
rect 9014 3522 9048 3556
rect 9086 3522 9120 3556
rect 9158 3522 9192 3556
rect 9230 3522 9264 3556
rect 9302 3522 9336 3556
rect 9374 3522 9408 3556
rect 9446 3522 9480 3556
rect 9518 3522 9552 3556
rect 9590 3522 9624 3556
rect 9662 3522 9696 3556
rect 9734 3522 9768 3556
rect 9806 3522 9840 3556
rect 9878 3522 9912 3556
rect 9950 3522 9984 3556
rect 10022 3522 10056 3556
rect 10094 3522 10128 3556
rect 10166 3522 10200 3556
rect 10238 3522 10272 3556
rect 10310 3522 10344 3556
rect 10382 3522 10416 3556
rect 10454 3522 10488 3556
rect 10526 3522 10560 3556
rect 10598 3522 10632 3556
rect 10670 3522 10704 3556
rect 10742 3522 10776 3556
rect 10814 3522 10848 3556
rect 10886 3522 10920 3556
rect 10958 3522 10992 3556
rect 11030 3522 11064 3556
rect 11102 3522 11136 3556
rect 11174 3522 11208 3556
rect 1677 3486 1711 3510
rect 1785 3476 1817 3484
rect 1817 3476 1819 3484
rect 1785 3450 1819 3476
rect 345 3408 368 3442
rect 368 3408 379 3442
rect 420 3408 436 3442
rect 436 3408 454 3442
rect 494 3408 504 3442
rect 504 3408 528 3442
rect 568 3408 572 3442
rect 572 3408 602 3442
rect 642 3408 674 3442
rect 674 3408 676 3442
rect 716 3408 742 3442
rect 742 3408 750 3442
rect 791 3408 810 3442
rect 810 3408 825 3442
rect 866 3408 878 3442
rect 878 3408 900 3442
rect 941 3408 946 3442
rect 946 3408 975 3442
rect 1016 3408 1048 3442
rect 1048 3408 1050 3442
rect 1091 3408 1116 3442
rect 1116 3408 1125 3442
rect 1166 3408 1184 3442
rect 1184 3408 1200 3442
rect 1241 3408 1252 3442
rect 1252 3408 1275 3442
rect 1316 3408 1320 3442
rect 1320 3408 1350 3442
rect 270 3340 304 3370
rect 270 3336 304 3340
rect 1388 3366 1422 3370
rect 1388 3336 1422 3366
rect 270 3272 304 3297
rect 270 3263 304 3272
rect 270 3204 304 3224
rect 270 3190 304 3204
rect 270 3136 304 3151
rect 270 3117 304 3136
rect 270 3068 304 3078
rect 270 3044 304 3068
rect 270 3000 304 3005
rect 270 2971 304 3000
rect 270 2898 304 2932
rect 270 2830 304 2859
rect 270 2825 304 2830
rect 270 2762 304 2786
rect 270 2752 304 2762
rect 270 2694 304 2713
rect 270 2679 304 2694
rect 270 2626 304 2640
rect 270 2606 304 2626
rect 270 2558 304 2567
rect 270 2533 304 2558
rect 270 2490 304 2494
rect 270 2460 304 2490
rect 270 2388 304 2421
rect 270 2387 304 2388
rect 270 2320 304 2348
rect 270 2314 304 2320
rect 270 2252 304 2276
rect 270 2242 304 2252
rect 270 2184 304 2204
rect 270 2170 304 2184
rect 270 2116 304 2132
rect 270 2098 304 2116
rect 270 2048 304 2060
rect 270 2026 304 2048
rect 270 1980 304 1988
rect 270 1954 304 1980
rect 369 3288 403 3322
rect 369 3214 403 3248
rect 369 3140 403 3174
rect 369 3066 403 3100
rect 553 3288 587 3322
rect 553 3214 587 3248
rect 553 3140 587 3174
rect 369 2992 403 3026
rect 369 2917 403 2951
rect 369 2842 403 2876
rect 369 2767 403 2801
rect 369 2692 403 2726
rect 369 2617 403 2651
rect 369 2542 403 2576
rect 369 2467 403 2501
rect 369 2392 403 2426
rect 369 2317 403 2351
rect 369 2242 403 2276
rect 369 2167 403 2201
rect 369 2092 403 2126
rect 369 2017 403 2051
rect 461 3054 495 3088
rect 461 2981 495 3015
rect 461 2908 495 2942
rect 461 2835 495 2869
rect 461 2762 495 2796
rect 461 2689 495 2723
rect 461 2616 495 2650
rect 461 2543 495 2577
rect 461 2470 495 2504
rect 461 2397 495 2431
rect 461 2324 495 2358
rect 461 2250 495 2284
rect 461 2176 495 2210
rect 461 2102 495 2136
rect 461 2028 495 2062
rect 553 3066 587 3100
rect 737 3288 771 3322
rect 737 3214 771 3248
rect 737 3140 771 3174
rect 553 2992 587 3026
rect 553 2917 587 2951
rect 553 2842 587 2876
rect 553 2767 587 2801
rect 553 2692 587 2726
rect 553 2617 587 2651
rect 553 2542 587 2576
rect 553 2467 587 2501
rect 553 2392 587 2426
rect 553 2317 587 2351
rect 553 2242 587 2276
rect 553 2167 587 2201
rect 553 2092 587 2126
rect 369 1942 403 1976
rect 553 2017 587 2051
rect 645 3054 679 3088
rect 645 2981 679 3015
rect 645 2908 679 2942
rect 645 2835 679 2869
rect 645 2762 679 2796
rect 645 2689 679 2723
rect 645 2616 679 2650
rect 645 2543 679 2577
rect 645 2470 679 2504
rect 645 2397 679 2431
rect 645 2324 679 2358
rect 645 2250 679 2284
rect 645 2176 679 2210
rect 645 2102 679 2136
rect 645 2028 679 2062
rect 737 3066 771 3100
rect 921 3288 955 3322
rect 921 3214 955 3248
rect 921 3140 955 3174
rect 737 2992 771 3026
rect 737 2917 771 2951
rect 737 2842 771 2876
rect 737 2767 771 2801
rect 737 2692 771 2726
rect 737 2617 771 2651
rect 737 2542 771 2576
rect 737 2467 771 2501
rect 737 2392 771 2426
rect 737 2317 771 2351
rect 737 2242 771 2276
rect 737 2167 771 2201
rect 737 2092 771 2126
rect 553 1942 587 1976
rect 737 2017 771 2051
rect 829 3054 863 3088
rect 829 2981 863 3015
rect 829 2908 863 2942
rect 829 2835 863 2869
rect 829 2762 863 2796
rect 829 2689 863 2723
rect 829 2616 863 2650
rect 829 2543 863 2577
rect 829 2470 863 2504
rect 829 2397 863 2431
rect 829 2324 863 2358
rect 829 2250 863 2284
rect 829 2176 863 2210
rect 829 2102 863 2136
rect 829 2028 863 2062
rect 921 3066 955 3100
rect 1105 3288 1139 3322
rect 1105 3214 1139 3248
rect 1105 3140 1139 3174
rect 921 2992 955 3026
rect 921 2917 955 2951
rect 921 2842 955 2876
rect 921 2767 955 2801
rect 921 2692 955 2726
rect 921 2617 955 2651
rect 921 2542 955 2576
rect 921 2467 955 2501
rect 921 2392 955 2426
rect 921 2317 955 2351
rect 921 2242 955 2276
rect 921 2167 955 2201
rect 921 2092 955 2126
rect 737 1942 771 1976
rect 921 2017 955 2051
rect 1013 3054 1047 3088
rect 1013 2981 1047 3015
rect 1013 2908 1047 2942
rect 1013 2835 1047 2869
rect 1013 2762 1047 2796
rect 1013 2689 1047 2723
rect 1013 2616 1047 2650
rect 1013 2543 1047 2577
rect 1013 2470 1047 2504
rect 1013 2397 1047 2431
rect 1013 2324 1047 2358
rect 1013 2250 1047 2284
rect 1013 2176 1047 2210
rect 1013 2102 1047 2136
rect 1013 2028 1047 2062
rect 1105 3066 1139 3100
rect 1289 3288 1323 3322
rect 1289 3214 1323 3248
rect 1289 3140 1323 3174
rect 1105 2992 1139 3026
rect 1105 2917 1139 2951
rect 1105 2842 1139 2876
rect 1105 2767 1139 2801
rect 1105 2692 1139 2726
rect 1105 2617 1139 2651
rect 1105 2542 1139 2576
rect 1105 2467 1139 2501
rect 1105 2392 1139 2426
rect 1105 2317 1139 2351
rect 1105 2242 1139 2276
rect 1105 2167 1139 2201
rect 1105 2092 1139 2126
rect 921 1942 955 1976
rect 1105 2017 1139 2051
rect 1197 3054 1231 3088
rect 1197 2981 1231 3015
rect 1197 2908 1231 2942
rect 1197 2835 1231 2869
rect 1197 2762 1231 2796
rect 1197 2689 1231 2723
rect 1197 2616 1231 2650
rect 1197 2543 1231 2577
rect 1197 2470 1231 2504
rect 1197 2397 1231 2431
rect 1197 2324 1231 2358
rect 1197 2250 1231 2284
rect 1197 2176 1231 2210
rect 1197 2102 1231 2136
rect 1197 2028 1231 2062
rect 1289 3066 1323 3100
rect 1289 2992 1323 3026
rect 1289 2917 1323 2951
rect 1289 2842 1323 2876
rect 1289 2767 1323 2801
rect 1289 2692 1323 2726
rect 1289 2617 1323 2651
rect 1289 2542 1323 2576
rect 1289 2467 1323 2501
rect 1289 2392 1323 2426
rect 1289 2317 1323 2351
rect 1289 2242 1323 2276
rect 1289 2167 1323 2201
rect 1289 2092 1323 2126
rect 1105 1942 1139 1976
rect 1289 2017 1323 2051
rect 1289 1942 1323 1976
rect 1388 3264 1422 3298
rect 1388 3196 1422 3226
rect 1388 3192 1422 3196
rect 1388 3128 1422 3154
rect 1388 3120 1422 3128
rect 1388 3060 1422 3082
rect 1388 3048 1422 3060
rect 1388 2992 1422 3010
rect 1388 2976 1422 2992
rect 1388 2924 1422 2938
rect 1388 2904 1422 2924
rect 1388 2856 1422 2866
rect 1388 2832 1422 2856
rect 1388 2788 1422 2794
rect 1388 2760 1422 2788
rect 1388 2720 1422 2722
rect 1388 2688 1422 2720
rect 1388 2618 1422 2650
rect 1388 2616 1422 2618
rect 1388 2550 1422 2578
rect 1388 2544 1422 2550
rect 1388 2482 1422 2506
rect 1388 2472 1422 2482
rect 1388 2414 1422 2434
rect 1388 2400 1422 2414
rect 1388 2346 1422 2362
rect 1388 2328 1422 2346
rect 1388 2278 1422 2290
rect 1388 2256 1422 2278
rect 1388 2210 1422 2218
rect 1388 2184 1422 2210
rect 1388 2142 1422 2146
rect 1388 2112 1422 2142
rect 1388 2040 1422 2074
rect 1388 1972 1422 2002
rect 1388 1968 1422 1972
rect 270 1912 304 1916
rect 270 1882 304 1912
rect 1388 1904 1422 1930
rect 1388 1896 1422 1904
rect 270 1810 304 1844
rect 1388 1836 1422 1858
rect 1388 1824 1422 1836
rect 270 1742 304 1772
rect 270 1738 304 1742
rect 270 1674 304 1700
rect 270 1666 304 1674
rect 270 1606 304 1628
rect 270 1594 304 1606
rect 270 1538 304 1556
rect 270 1522 304 1538
rect 270 1470 304 1484
rect 270 1450 304 1470
rect 270 1402 304 1412
rect 270 1378 304 1402
rect 270 1334 304 1340
rect 270 1306 304 1334
rect 270 1266 304 1268
rect 270 1234 304 1266
rect 270 1164 304 1196
rect 270 1162 304 1164
rect 270 1096 304 1124
rect 270 1090 304 1096
rect 270 1028 304 1052
rect 270 1018 304 1028
rect 270 960 304 980
rect 270 946 304 960
rect 270 892 304 908
rect 270 874 304 892
rect 369 1758 403 1792
rect 369 1684 403 1718
rect 369 1610 403 1644
rect 369 1536 403 1570
rect 369 1462 403 1496
rect 369 1388 403 1422
rect 369 1314 403 1348
rect 369 1240 403 1274
rect 369 1166 403 1200
rect 369 1092 403 1126
rect 369 1018 403 1052
rect 369 944 403 978
rect 369 869 403 903
rect 369 794 403 828
rect 369 719 403 753
rect 369 644 403 678
rect 461 1758 495 1792
rect 461 1684 495 1718
rect 461 1610 495 1644
rect 461 1536 495 1570
rect 461 1462 495 1496
rect 461 1388 495 1422
rect 461 1314 495 1348
rect 461 1240 495 1274
rect 461 1166 495 1200
rect 461 1092 495 1126
rect 461 1018 495 1052
rect 461 944 495 978
rect 461 870 495 904
rect 461 796 495 830
rect 461 722 495 756
rect 461 648 495 682
rect 553 1758 587 1792
rect 553 1684 587 1718
rect 553 1610 587 1644
rect 553 1536 587 1570
rect 553 1462 587 1496
rect 553 1388 587 1422
rect 553 1314 587 1348
rect 553 1240 587 1274
rect 553 1166 587 1200
rect 553 1092 587 1126
rect 553 1018 587 1052
rect 553 944 587 978
rect 553 869 587 903
rect 553 794 587 828
rect 553 719 587 753
rect 553 644 587 678
rect 645 1758 679 1792
rect 645 1684 679 1718
rect 645 1610 679 1644
rect 645 1536 679 1570
rect 645 1462 679 1496
rect 645 1388 679 1422
rect 645 1314 679 1348
rect 645 1240 679 1274
rect 645 1166 679 1200
rect 645 1092 679 1126
rect 645 1018 679 1052
rect 645 944 679 978
rect 645 870 679 904
rect 645 796 679 830
rect 645 722 679 756
rect 645 648 679 682
rect 461 573 495 607
rect 461 498 495 532
rect 737 1758 771 1792
rect 737 1684 771 1718
rect 737 1610 771 1644
rect 737 1536 771 1570
rect 737 1462 771 1496
rect 737 1388 771 1422
rect 737 1314 771 1348
rect 737 1240 771 1274
rect 737 1166 771 1200
rect 737 1092 771 1126
rect 737 1018 771 1052
rect 737 944 771 978
rect 737 869 771 903
rect 737 794 771 828
rect 737 719 771 753
rect 737 644 771 678
rect 829 1758 863 1792
rect 829 1684 863 1718
rect 829 1610 863 1644
rect 829 1536 863 1570
rect 829 1462 863 1496
rect 829 1388 863 1422
rect 829 1314 863 1348
rect 829 1240 863 1274
rect 829 1166 863 1200
rect 829 1092 863 1126
rect 829 1018 863 1052
rect 829 944 863 978
rect 829 870 863 904
rect 829 796 863 830
rect 829 722 863 756
rect 829 648 863 682
rect 645 573 679 607
rect 645 498 679 532
rect 921 1758 955 1792
rect 921 1684 955 1718
rect 921 1610 955 1644
rect 921 1536 955 1570
rect 921 1462 955 1496
rect 921 1388 955 1422
rect 921 1314 955 1348
rect 921 1240 955 1274
rect 921 1166 955 1200
rect 921 1092 955 1126
rect 921 1018 955 1052
rect 921 944 955 978
rect 921 869 955 903
rect 921 794 955 828
rect 921 719 955 753
rect 921 644 955 678
rect 1013 1758 1047 1792
rect 1013 1684 1047 1718
rect 1013 1610 1047 1644
rect 1013 1536 1047 1570
rect 1013 1462 1047 1496
rect 1013 1388 1047 1422
rect 1013 1314 1047 1348
rect 1013 1240 1047 1274
rect 1013 1166 1047 1200
rect 1013 1092 1047 1126
rect 1013 1018 1047 1052
rect 1013 944 1047 978
rect 1013 870 1047 904
rect 1013 796 1047 830
rect 1013 722 1047 756
rect 1013 648 1047 682
rect 829 573 863 607
rect 829 498 863 532
rect 1105 1758 1139 1792
rect 1105 1684 1139 1718
rect 1105 1610 1139 1644
rect 1105 1536 1139 1570
rect 1105 1462 1139 1496
rect 1105 1388 1139 1422
rect 1105 1314 1139 1348
rect 1105 1240 1139 1274
rect 1105 1166 1139 1200
rect 1105 1092 1139 1126
rect 1105 1018 1139 1052
rect 1105 944 1139 978
rect 1105 869 1139 903
rect 1105 794 1139 828
rect 1105 719 1139 753
rect 1105 644 1139 678
rect 1197 1758 1231 1792
rect 1197 1684 1231 1718
rect 1197 1610 1231 1644
rect 1197 1536 1231 1570
rect 1197 1462 1231 1496
rect 1197 1388 1231 1422
rect 1197 1314 1231 1348
rect 1197 1240 1231 1274
rect 1197 1166 1231 1200
rect 1197 1092 1231 1126
rect 1197 1018 1231 1052
rect 1197 944 1231 978
rect 1197 870 1231 904
rect 1197 796 1231 830
rect 1197 722 1231 756
rect 1197 648 1231 682
rect 1013 573 1047 607
rect 1013 498 1047 532
rect 1197 573 1231 607
rect 1197 498 1231 532
rect 1289 1758 1323 1792
rect 1289 1684 1323 1718
rect 1289 1610 1323 1644
rect 1289 1536 1323 1570
rect 1289 1462 1323 1496
rect 1289 1387 1323 1421
rect 1289 1312 1323 1346
rect 1289 1237 1323 1271
rect 1289 1162 1323 1196
rect 1289 1087 1323 1121
rect 1289 1012 1323 1046
rect 1289 937 1323 971
rect 1289 862 1323 896
rect 1289 787 1323 821
rect 1289 712 1323 746
rect 1289 637 1323 671
rect 1289 562 1323 596
rect 1289 487 1323 521
rect 1289 412 1323 446
rect 1388 1768 1422 1785
rect 1388 1751 1422 1768
rect 1388 1700 1422 1712
rect 1388 1678 1422 1700
rect 1388 1632 1422 1639
rect 1388 1605 1422 1632
rect 1388 1564 1422 1566
rect 1388 1532 1422 1564
rect 1388 1462 1422 1493
rect 1388 1459 1422 1462
rect 1388 1394 1422 1420
rect 1388 1386 1422 1394
rect 1388 1326 1422 1347
rect 1388 1313 1422 1326
rect 1388 1258 1422 1274
rect 1388 1240 1422 1258
rect 1388 1190 1422 1201
rect 1388 1167 1422 1190
rect 1388 1122 1422 1128
rect 1388 1094 1422 1122
rect 1388 1054 1422 1055
rect 1388 1021 1422 1054
rect 1388 952 1422 982
rect 1388 948 1422 952
rect 1388 884 1422 909
rect 1388 875 1422 884
rect 1388 816 1422 836
rect 1388 802 1422 816
rect 1388 748 1422 763
rect 1388 729 1422 748
rect 1388 680 1422 690
rect 1388 656 1422 680
rect 426 322 430 356
rect 430 322 460 356
rect 500 322 503 356
rect 503 322 534 356
rect 574 322 576 356
rect 576 322 608 356
rect 648 322 649 356
rect 649 322 682 356
rect 721 322 722 356
rect 722 322 755 356
rect 794 322 795 356
rect 795 322 828 356
rect 867 322 868 356
rect 868 322 901 356
rect 940 322 974 356
rect 1013 322 1046 356
rect 1046 322 1047 356
rect 1086 322 1118 356
rect 1118 322 1120 356
rect 1159 322 1190 356
rect 1190 322 1193 356
rect 1232 322 1262 356
rect 1262 322 1266 356
rect 1677 3442 1711 3448
rect 1892 3442 1926 3461
rect 1967 3442 2001 3461
rect 2042 3442 2076 3461
rect 2117 3442 2151 3461
rect 2192 3442 2226 3461
rect 2266 3442 2300 3461
rect 2340 3442 2374 3461
rect 2414 3442 2448 3461
rect 2488 3442 2522 3461
rect 2562 3442 2596 3461
rect 2636 3442 2670 3461
rect 2710 3442 2744 3461
rect 2784 3442 2818 3461
rect 2858 3442 2892 3461
rect 2932 3442 2966 3461
rect 3006 3442 3040 3461
rect 3080 3442 3114 3461
rect 3154 3442 3188 3461
rect 3228 3442 3262 3461
rect 1677 3414 1711 3442
rect 1785 3408 1817 3412
rect 1817 3408 1819 3412
rect 1892 3427 1921 3442
rect 1921 3427 1926 3442
rect 1967 3427 1991 3442
rect 1991 3427 2001 3442
rect 2042 3427 2061 3442
rect 2061 3427 2076 3442
rect 2117 3427 2131 3442
rect 2131 3427 2151 3442
rect 2192 3427 2201 3442
rect 2201 3427 2226 3442
rect 2266 3427 2271 3442
rect 2271 3427 2300 3442
rect 2340 3427 2341 3442
rect 2341 3427 2374 3442
rect 2414 3427 2447 3442
rect 2447 3427 2448 3442
rect 2488 3427 2517 3442
rect 2517 3427 2522 3442
rect 2562 3427 2587 3442
rect 2587 3427 2596 3442
rect 2636 3427 2657 3442
rect 2657 3427 2670 3442
rect 2710 3427 2727 3442
rect 2727 3427 2744 3442
rect 2784 3427 2797 3442
rect 2797 3427 2818 3442
rect 2858 3427 2867 3442
rect 2867 3427 2892 3442
rect 2932 3427 2937 3442
rect 2937 3427 2966 3442
rect 3006 3427 3007 3442
rect 3007 3427 3040 3442
rect 3080 3427 3111 3442
rect 3111 3427 3114 3442
rect 3154 3427 3181 3442
rect 3181 3427 3188 3442
rect 3228 3427 3251 3442
rect 3251 3427 3262 3442
rect 1785 3378 1819 3408
rect 1677 3374 1711 3376
rect 1892 3374 1926 3389
rect 1967 3374 2001 3389
rect 2042 3374 2076 3389
rect 2117 3374 2151 3389
rect 2192 3374 2226 3389
rect 2266 3374 2300 3389
rect 2340 3374 2374 3389
rect 2414 3374 2448 3389
rect 2488 3374 2522 3389
rect 2562 3374 2596 3389
rect 2636 3374 2670 3389
rect 2710 3374 2744 3389
rect 2784 3374 2818 3389
rect 2858 3374 2892 3389
rect 2932 3374 2966 3389
rect 3006 3374 3040 3389
rect 3080 3374 3114 3389
rect 3154 3374 3188 3389
rect 3228 3374 3262 3389
rect 13623 3420 13655 3454
rect 13655 3420 13657 3454
rect 13747 3420 13757 3454
rect 13757 3420 13781 3454
rect 13821 3420 13825 3454
rect 13825 3420 13855 3454
rect 13895 3420 13927 3454
rect 13927 3420 13929 3454
rect 13969 3420 13995 3454
rect 13995 3420 14003 3454
rect 14044 3420 14063 3454
rect 14063 3420 14078 3454
rect 14119 3420 14131 3454
rect 14131 3420 14153 3454
rect 14194 3420 14199 3454
rect 14199 3420 14228 3454
rect 14269 3420 14301 3454
rect 14301 3420 14303 3454
rect 14344 3420 14369 3454
rect 14369 3420 14378 3454
rect 14419 3420 14437 3454
rect 14437 3420 14453 3454
rect 14494 3420 14505 3454
rect 14505 3420 14528 3454
rect 14569 3420 14573 3454
rect 14573 3420 14603 3454
rect 1677 3342 1711 3374
rect 1892 3355 1921 3374
rect 1921 3355 1926 3374
rect 1967 3355 1991 3374
rect 1991 3355 2001 3374
rect 2042 3355 2061 3374
rect 2061 3355 2076 3374
rect 2117 3355 2131 3374
rect 2131 3355 2151 3374
rect 2192 3355 2201 3374
rect 2201 3355 2226 3374
rect 2266 3355 2271 3374
rect 2271 3355 2300 3374
rect 2340 3355 2341 3374
rect 2341 3355 2374 3374
rect 2414 3355 2447 3374
rect 2447 3355 2448 3374
rect 2488 3355 2517 3374
rect 2517 3355 2522 3374
rect 2562 3355 2587 3374
rect 2587 3355 2596 3374
rect 2636 3355 2657 3374
rect 2657 3355 2670 3374
rect 2710 3355 2727 3374
rect 2727 3355 2744 3374
rect 2784 3355 2797 3374
rect 2797 3355 2818 3374
rect 2858 3355 2867 3374
rect 2867 3355 2892 3374
rect 2932 3355 2937 3374
rect 2937 3355 2966 3374
rect 3006 3355 3007 3374
rect 3007 3355 3040 3374
rect 3080 3355 3111 3374
rect 3111 3355 3114 3374
rect 3154 3355 3181 3374
rect 3181 3355 3188 3374
rect 3228 3355 3251 3374
rect 3251 3355 3262 3374
rect 1785 3306 1819 3340
rect 1892 3306 1926 3317
rect 1967 3306 2001 3317
rect 2042 3306 2076 3317
rect 2117 3306 2151 3317
rect 2192 3306 2226 3317
rect 2266 3306 2300 3317
rect 2340 3306 2374 3317
rect 2414 3306 2448 3317
rect 2488 3306 2522 3317
rect 2562 3306 2596 3317
rect 2636 3306 2670 3317
rect 2710 3306 2744 3317
rect 2784 3306 2818 3317
rect 2858 3306 2892 3317
rect 2932 3306 2966 3317
rect 3006 3306 3040 3317
rect 3080 3306 3114 3317
rect 3154 3306 3188 3317
rect 3228 3306 3262 3317
rect 1677 3272 1711 3304
rect 1892 3283 1921 3306
rect 1921 3283 1926 3306
rect 1967 3283 1991 3306
rect 1991 3283 2001 3306
rect 2042 3283 2061 3306
rect 2061 3283 2076 3306
rect 2117 3283 2131 3306
rect 2131 3283 2151 3306
rect 2192 3283 2201 3306
rect 2201 3283 2226 3306
rect 2266 3283 2271 3306
rect 2271 3283 2300 3306
rect 2340 3283 2341 3306
rect 2341 3283 2374 3306
rect 2414 3283 2447 3306
rect 2447 3283 2448 3306
rect 2488 3283 2517 3306
rect 2517 3283 2522 3306
rect 2562 3283 2587 3306
rect 2587 3283 2596 3306
rect 2636 3283 2657 3306
rect 2657 3283 2670 3306
rect 2710 3283 2727 3306
rect 2727 3283 2744 3306
rect 2784 3283 2797 3306
rect 2797 3283 2818 3306
rect 2858 3283 2867 3306
rect 2867 3283 2892 3306
rect 2932 3283 2937 3306
rect 2937 3283 2966 3306
rect 3006 3283 3007 3306
rect 3007 3283 3040 3306
rect 3080 3283 3111 3306
rect 3111 3283 3114 3306
rect 3154 3283 3181 3306
rect 3181 3283 3188 3306
rect 3228 3283 3251 3306
rect 3251 3283 3262 3306
rect 11396 3273 11502 3379
rect 13523 3352 13557 3382
rect 13523 3348 13557 3352
rect 14641 3378 14675 3382
rect 14641 3348 14675 3378
rect 13523 3284 13557 3309
rect 13523 3275 13557 3284
rect 1677 3270 1711 3272
rect 1785 3238 1819 3268
rect 1892 3238 1926 3245
rect 1967 3238 2001 3245
rect 2042 3238 2076 3245
rect 2117 3238 2151 3245
rect 2192 3238 2226 3245
rect 2266 3238 2300 3245
rect 2340 3238 2374 3245
rect 2414 3238 2448 3245
rect 2488 3238 2522 3245
rect 2562 3238 2596 3245
rect 2636 3238 2670 3245
rect 2710 3238 2744 3245
rect 2784 3238 2818 3245
rect 2858 3238 2892 3245
rect 2932 3238 2966 3245
rect 3006 3238 3040 3245
rect 3080 3238 3114 3245
rect 3154 3238 3188 3245
rect 3228 3238 3262 3245
rect 1677 3204 1711 3232
rect 1785 3234 1817 3238
rect 1817 3234 1819 3238
rect 1892 3211 1921 3238
rect 1921 3211 1926 3238
rect 1967 3211 1991 3238
rect 1991 3211 2001 3238
rect 2042 3211 2061 3238
rect 2061 3211 2076 3238
rect 2117 3211 2131 3238
rect 2131 3211 2151 3238
rect 2192 3211 2201 3238
rect 2201 3211 2226 3238
rect 2266 3211 2271 3238
rect 2271 3211 2300 3238
rect 2340 3211 2341 3238
rect 2341 3211 2374 3238
rect 2414 3211 2447 3238
rect 2447 3211 2448 3238
rect 2488 3211 2517 3238
rect 2517 3211 2522 3238
rect 2562 3211 2587 3238
rect 2587 3211 2596 3238
rect 2636 3211 2657 3238
rect 2657 3211 2670 3238
rect 2710 3211 2727 3238
rect 2727 3211 2744 3238
rect 2784 3211 2797 3238
rect 2797 3211 2818 3238
rect 2858 3211 2867 3238
rect 2867 3211 2892 3238
rect 2932 3211 2937 3238
rect 2937 3211 2966 3238
rect 3006 3211 3007 3238
rect 3007 3211 3040 3238
rect 3080 3211 3111 3238
rect 3111 3211 3114 3238
rect 3154 3211 3181 3238
rect 3181 3211 3188 3238
rect 3228 3211 3251 3238
rect 3251 3211 3262 3238
rect 1677 3198 1711 3204
rect 1785 3169 1819 3196
rect 1892 3169 1926 3173
rect 1967 3169 2001 3173
rect 2042 3169 2076 3173
rect 2117 3169 2151 3173
rect 2192 3169 2226 3173
rect 2266 3169 2300 3173
rect 2340 3169 2374 3173
rect 2414 3169 2448 3173
rect 2488 3169 2522 3173
rect 2562 3169 2596 3173
rect 2636 3169 2670 3173
rect 2710 3169 2744 3173
rect 2784 3169 2818 3173
rect 2858 3169 2892 3173
rect 2932 3169 2966 3173
rect 3006 3169 3040 3173
rect 3080 3169 3114 3173
rect 3154 3169 3188 3173
rect 3228 3169 3262 3173
rect 1677 3135 1711 3160
rect 1785 3162 1817 3169
rect 1817 3162 1819 3169
rect 1892 3139 1921 3169
rect 1921 3139 1926 3169
rect 1967 3139 1991 3169
rect 1991 3139 2001 3169
rect 2042 3139 2061 3169
rect 2061 3139 2076 3169
rect 2117 3139 2131 3169
rect 2131 3139 2151 3169
rect 2192 3139 2201 3169
rect 2201 3139 2226 3169
rect 2266 3139 2271 3169
rect 2271 3139 2300 3169
rect 2340 3139 2341 3169
rect 2341 3139 2374 3169
rect 2414 3139 2447 3169
rect 2447 3139 2448 3169
rect 2488 3139 2517 3169
rect 2517 3139 2522 3169
rect 2562 3139 2587 3169
rect 2587 3139 2596 3169
rect 2636 3139 2657 3169
rect 2657 3139 2670 3169
rect 2710 3139 2727 3169
rect 2727 3139 2744 3169
rect 2784 3139 2797 3169
rect 2797 3139 2818 3169
rect 2858 3139 2867 3169
rect 2867 3139 2892 3169
rect 2932 3139 2937 3169
rect 2937 3139 2966 3169
rect 3006 3139 3007 3169
rect 3007 3139 3040 3169
rect 3080 3139 3111 3169
rect 3111 3139 3114 3169
rect 3154 3139 3181 3169
rect 3181 3139 3188 3169
rect 3228 3139 3251 3169
rect 3251 3139 3262 3169
rect 1677 3126 1711 3135
rect 1785 3100 1819 3124
rect 1677 3066 1711 3088
rect 1785 3090 1817 3100
rect 1817 3090 1819 3100
rect 1677 3054 1711 3066
rect 1785 3031 1819 3052
rect 1677 2997 1711 3016
rect 1785 3018 1817 3031
rect 1817 3018 1819 3031
rect 1677 2982 1711 2997
rect 1785 2962 1819 2980
rect 1677 2928 1711 2944
rect 1785 2946 1817 2962
rect 1817 2946 1819 2962
rect 1677 2910 1711 2928
rect 1785 2893 1819 2908
rect 1677 2859 1711 2872
rect 1785 2874 1817 2893
rect 1817 2874 1819 2893
rect 1677 2838 1711 2859
rect 1785 2824 1819 2836
rect 1677 2790 1711 2800
rect 1785 2802 1817 2824
rect 1817 2802 1819 2824
rect 1677 2766 1711 2790
rect 1785 2755 1819 2764
rect 1677 2721 1711 2728
rect 1785 2730 1817 2755
rect 1817 2730 1819 2755
rect 1677 2694 1711 2721
rect 1785 2686 1819 2692
rect 1677 2652 1711 2656
rect 1785 2658 1817 2686
rect 1817 2658 1819 2686
rect 1677 2622 1711 2652
rect 1785 2617 1819 2620
rect 1677 2583 1711 2584
rect 1785 2586 1817 2617
rect 1817 2586 1819 2617
rect 1677 2550 1711 2583
rect 1785 2514 1817 2547
rect 1817 2514 1819 2547
rect 1785 2513 1819 2514
rect 1677 2479 1711 2511
rect 1677 2477 1711 2479
rect 1785 2445 1817 2474
rect 1817 2445 1819 2474
rect 1785 2440 1819 2445
rect 1677 2410 1711 2438
rect 1677 2404 1711 2410
rect 1785 2376 1817 2401
rect 1817 2376 1819 2401
rect 1785 2367 1819 2376
rect 1677 2341 1711 2365
rect 1677 2331 1711 2341
rect 1785 2307 1817 2328
rect 1817 2307 1819 2328
rect 1785 2294 1819 2307
rect 1677 2272 1711 2292
rect 1677 2258 1711 2272
rect 1785 2238 1817 2255
rect 1817 2238 1819 2255
rect 1785 2221 1819 2238
rect 1677 2203 1711 2219
rect 1677 2185 1711 2203
rect 1785 2169 1817 2182
rect 1817 2169 1819 2182
rect 1785 2148 1819 2169
rect 1677 2134 1711 2146
rect 1677 2112 1711 2134
rect 1785 2100 1817 2109
rect 1817 2100 1819 2109
rect 1785 2075 1819 2100
rect 1677 2065 1711 2073
rect 1677 2039 1711 2065
rect 1785 2031 1817 2036
rect 1817 2031 1819 2036
rect 1785 2002 1819 2031
rect 1677 1996 1711 2000
rect 1677 1966 1711 1996
rect 1785 1962 1817 1963
rect 1817 1962 1819 1963
rect 1785 1929 1819 1962
rect 1677 1893 1711 1927
rect 1785 1858 1819 1890
rect 1677 1824 1711 1854
rect 1785 1856 1817 1858
rect 1817 1856 1819 1858
rect 1677 1820 1711 1824
rect 1785 1789 1819 1817
rect 1677 1755 1711 1781
rect 1785 1783 1817 1789
rect 1817 1783 1819 1789
rect 1677 1747 1711 1755
rect 1785 1720 1819 1744
rect 1677 1686 1711 1708
rect 1785 1710 1817 1720
rect 1817 1710 1819 1720
rect 1677 1674 1711 1686
rect 1785 1651 1819 1671
rect 1677 1617 1711 1635
rect 1785 1637 1817 1651
rect 1817 1637 1819 1651
rect 1677 1601 1711 1617
rect 1785 1582 1819 1598
rect 1677 1548 1711 1562
rect 1785 1564 1817 1582
rect 1817 1564 1819 1582
rect 1677 1528 1711 1548
rect 1785 1513 1819 1525
rect 1677 1479 1711 1489
rect 1785 1491 1817 1513
rect 1817 1491 1819 1513
rect 1677 1455 1711 1479
rect 1785 1444 1819 1452
rect 1677 1410 1711 1416
rect 1785 1418 1817 1444
rect 1817 1418 1819 1444
rect 1677 1382 1711 1410
rect 1785 1375 1819 1379
rect 1677 1341 1711 1343
rect 1785 1345 1817 1375
rect 1817 1345 1819 1375
rect 1677 1309 1711 1341
rect 1785 1272 1817 1306
rect 1817 1272 1819 1306
rect 1677 1237 1711 1270
rect 1677 1236 1711 1237
rect 1785 1203 1817 1233
rect 1817 1203 1819 1233
rect 1785 1199 1819 1203
rect 1677 1168 1711 1197
rect 1677 1163 1711 1168
rect 1785 1134 1817 1160
rect 1817 1134 1819 1160
rect 1785 1126 1819 1134
rect 1677 1099 1711 1124
rect 1677 1090 1711 1099
rect 1785 1065 1817 1087
rect 1817 1065 1819 1087
rect 1785 1053 1819 1065
rect 1677 1030 1711 1051
rect 1677 1017 1711 1030
rect 1785 996 1817 1014
rect 1817 996 1819 1014
rect 1785 980 1819 996
rect 1677 961 1711 978
rect 1677 944 1711 961
rect 1785 927 1817 941
rect 1817 927 1819 941
rect 1785 907 1819 927
rect 1677 892 1711 905
rect 1677 871 1711 892
rect 1785 858 1817 868
rect 1817 858 1819 868
rect 1785 834 1819 858
rect 1677 823 1711 832
rect 1677 798 1711 823
rect 1785 789 1817 795
rect 1817 789 1819 795
rect 1785 761 1819 789
rect 1677 754 1711 759
rect 1677 725 1711 754
rect 1785 720 1817 722
rect 1817 720 1819 722
rect 1785 688 1819 720
rect 1677 685 1711 686
rect 1677 652 1711 685
rect 1785 616 1819 649
rect 1677 582 1711 613
rect 1785 615 1817 616
rect 1817 615 1819 616
rect 1677 579 1711 582
rect 1785 547 1819 576
rect 1892 548 1926 582
rect 1967 548 2001 582
rect 2042 548 2076 582
rect 2117 548 2151 582
rect 2192 548 2226 582
rect 2266 548 2300 582
rect 2340 548 2374 582
rect 2414 548 2448 582
rect 2488 548 2522 582
rect 2562 548 2596 582
rect 2636 548 2670 582
rect 2710 548 2744 582
rect 2784 548 2818 582
rect 2858 548 2892 582
rect 2932 548 2966 582
rect 3006 548 3040 582
rect 3080 548 3114 582
rect 3154 548 3188 582
rect 3228 548 3262 582
rect 1677 513 1711 540
rect 1785 542 1817 547
rect 1817 542 1819 547
rect 1677 506 1711 513
rect 1785 478 1819 503
rect 1892 478 1926 510
rect 1967 478 2001 510
rect 2042 478 2076 510
rect 2117 478 2151 510
rect 2192 478 2226 510
rect 2266 478 2300 510
rect 2340 478 2374 510
rect 2414 478 2448 510
rect 2488 478 2522 510
rect 2562 478 2596 510
rect 2636 478 2670 510
rect 2710 478 2744 510
rect 2784 478 2818 510
rect 2858 478 2892 510
rect 2932 478 2966 510
rect 3006 478 3040 510
rect 3080 478 3114 510
rect 3154 478 3188 510
rect 3228 478 3262 510
rect 1677 444 1711 467
rect 1785 469 1817 478
rect 1817 469 1819 478
rect 1892 476 1921 478
rect 1921 476 1926 478
rect 1967 476 1991 478
rect 1991 476 2001 478
rect 2042 476 2061 478
rect 2061 476 2076 478
rect 2117 476 2131 478
rect 2131 476 2151 478
rect 2192 476 2201 478
rect 2201 476 2226 478
rect 2266 476 2271 478
rect 2271 476 2300 478
rect 2340 476 2341 478
rect 2341 476 2374 478
rect 2414 476 2447 478
rect 2447 476 2448 478
rect 2488 476 2517 478
rect 2517 476 2522 478
rect 2562 476 2587 478
rect 2587 476 2596 478
rect 2636 476 2657 478
rect 2657 476 2670 478
rect 2710 476 2727 478
rect 2727 476 2744 478
rect 2784 476 2797 478
rect 2797 476 2818 478
rect 2858 476 2867 478
rect 2867 476 2892 478
rect 2932 476 2937 478
rect 2937 476 2966 478
rect 3006 476 3007 478
rect 3007 476 3040 478
rect 3080 476 3111 478
rect 3111 476 3114 478
rect 3154 476 3181 478
rect 3181 476 3188 478
rect 3228 476 3251 478
rect 3251 476 3262 478
rect 1677 433 1711 444
rect 1785 409 1819 430
rect 1860 409 1894 430
rect 1935 409 1969 430
rect 2010 409 2044 430
rect 2085 409 2119 430
rect 2160 409 2194 430
rect 2235 409 2269 430
rect 2310 409 2344 430
rect 2385 409 2419 430
rect 2460 409 2494 430
rect 2535 409 2569 430
rect 2610 409 2644 430
rect 2685 409 2719 430
rect 2760 409 2794 430
rect 2835 409 2869 430
rect 2910 409 2944 430
rect 2985 409 3019 430
rect 3060 409 3094 430
rect 3135 409 3169 430
rect 3210 409 3244 430
rect 1677 375 1711 394
rect 1785 396 1817 409
rect 1817 396 1819 409
rect 1860 396 1887 409
rect 1887 396 1894 409
rect 1935 396 1957 409
rect 1957 396 1969 409
rect 2010 396 2027 409
rect 2027 396 2044 409
rect 2085 396 2097 409
rect 2097 396 2119 409
rect 2160 396 2167 409
rect 2167 396 2194 409
rect 2235 396 2237 409
rect 2237 396 2269 409
rect 2310 396 2341 409
rect 2341 396 2344 409
rect 2385 396 2411 409
rect 2411 396 2419 409
rect 2460 396 2481 409
rect 2481 396 2494 409
rect 2535 396 2551 409
rect 2551 396 2569 409
rect 2610 396 2621 409
rect 2621 396 2644 409
rect 2685 396 2691 409
rect 2691 396 2719 409
rect 2760 396 2761 409
rect 2761 396 2794 409
rect 2835 396 2867 409
rect 2867 396 2869 409
rect 2910 396 2937 409
rect 2937 396 2944 409
rect 2985 396 3007 409
rect 3007 396 3019 409
rect 3060 396 3077 409
rect 3077 396 3094 409
rect 3135 396 3147 409
rect 3147 396 3169 409
rect 3210 396 3217 409
rect 3217 396 3244 409
rect 1677 360 1711 375
rect 13523 3216 13557 3236
rect 13523 3202 13557 3216
rect 13523 3148 13557 3163
rect 13523 3129 13557 3148
rect 13523 3080 13557 3090
rect 13523 3056 13557 3080
rect 13523 3012 13557 3017
rect 13523 2983 13557 3012
rect 13523 2910 13557 2944
rect 13523 2842 13557 2871
rect 13523 2837 13557 2842
rect 13523 2774 13557 2798
rect 13523 2764 13557 2774
rect 13523 2706 13557 2725
rect 13523 2691 13557 2706
rect 13523 2638 13557 2652
rect 13523 2618 13557 2638
rect 13523 2570 13557 2579
rect 13523 2545 13557 2570
rect 13523 2502 13557 2506
rect 13523 2472 13557 2502
rect 13523 2400 13557 2433
rect 13523 2399 13557 2400
rect 13523 2332 13557 2360
rect 13523 2326 13557 2332
rect 13523 2264 13557 2287
rect 13523 2253 13557 2264
rect 13523 2196 13557 2214
rect 13523 2180 13557 2196
rect 13523 2128 13557 2141
rect 13523 2107 13557 2128
rect 13523 2060 13557 2068
rect 13523 2034 13557 2060
rect 13523 1992 13557 1995
rect 13523 1961 13557 1992
rect 13622 3300 13656 3334
rect 13622 3226 13656 3260
rect 13622 3152 13656 3186
rect 13806 3300 13840 3334
rect 13806 3226 13840 3260
rect 13806 3152 13840 3186
rect 13622 3078 13656 3112
rect 13622 3004 13656 3038
rect 13622 2929 13656 2963
rect 13622 2854 13656 2888
rect 13622 2779 13656 2813
rect 13622 2704 13656 2738
rect 13622 2629 13656 2663
rect 13622 2554 13656 2588
rect 13622 2479 13656 2513
rect 13622 2404 13656 2438
rect 13622 2329 13656 2363
rect 13622 2254 13656 2288
rect 13622 2179 13656 2213
rect 13622 2104 13656 2138
rect 13622 2029 13656 2063
rect 13714 3098 13748 3132
rect 13714 3023 13748 3057
rect 13714 2948 13748 2982
rect 13714 2873 13748 2907
rect 13714 2798 13748 2832
rect 13714 2723 13748 2757
rect 13714 2648 13748 2682
rect 13714 2572 13748 2606
rect 13714 2496 13748 2530
rect 13714 2420 13748 2454
rect 13714 2344 13748 2378
rect 13714 2268 13748 2302
rect 13714 2192 13748 2226
rect 13714 2116 13748 2150
rect 13714 2040 13748 2074
rect 13990 3300 14024 3334
rect 13990 3226 14024 3260
rect 13990 3152 14024 3186
rect 13806 3078 13840 3112
rect 13806 3004 13840 3038
rect 13806 2929 13840 2963
rect 13806 2854 13840 2888
rect 13806 2779 13840 2813
rect 13806 2704 13840 2738
rect 13806 2629 13840 2663
rect 13806 2554 13840 2588
rect 13806 2479 13840 2513
rect 13806 2404 13840 2438
rect 13806 2329 13840 2363
rect 13806 2254 13840 2288
rect 13806 2179 13840 2213
rect 13806 2104 13840 2138
rect 13622 1954 13656 1988
rect 13806 2029 13840 2063
rect 13898 3098 13932 3132
rect 13898 3023 13932 3057
rect 13898 2948 13932 2982
rect 13898 2873 13932 2907
rect 13898 2798 13932 2832
rect 13898 2723 13932 2757
rect 13898 2648 13932 2682
rect 13898 2572 13932 2606
rect 13898 2496 13932 2530
rect 13898 2420 13932 2454
rect 13898 2344 13932 2378
rect 13898 2268 13932 2302
rect 13898 2192 13932 2226
rect 13898 2116 13932 2150
rect 13898 2040 13932 2074
rect 14174 3300 14208 3334
rect 14174 3226 14208 3260
rect 14174 3152 14208 3186
rect 13990 3078 14024 3112
rect 13990 3004 14024 3038
rect 13990 2929 14024 2963
rect 13990 2854 14024 2888
rect 13990 2779 14024 2813
rect 13990 2704 14024 2738
rect 13990 2629 14024 2663
rect 13990 2554 14024 2588
rect 13990 2479 14024 2513
rect 13990 2404 14024 2438
rect 13990 2329 14024 2363
rect 13990 2254 14024 2288
rect 13990 2179 14024 2213
rect 13990 2104 14024 2138
rect 13806 1954 13840 1988
rect 13990 2029 14024 2063
rect 14082 3098 14116 3132
rect 14082 3023 14116 3057
rect 14082 2948 14116 2982
rect 14082 2873 14116 2907
rect 14082 2798 14116 2832
rect 14082 2723 14116 2757
rect 14082 2648 14116 2682
rect 14082 2572 14116 2606
rect 14082 2496 14116 2530
rect 14082 2420 14116 2454
rect 14082 2344 14116 2378
rect 14082 2268 14116 2302
rect 14082 2192 14116 2226
rect 14082 2116 14116 2150
rect 14082 2040 14116 2074
rect 14358 3300 14392 3334
rect 14358 3226 14392 3260
rect 14358 3152 14392 3186
rect 14174 3078 14208 3112
rect 14174 3004 14208 3038
rect 14174 2929 14208 2963
rect 14174 2854 14208 2888
rect 14174 2779 14208 2813
rect 14174 2704 14208 2738
rect 14174 2629 14208 2663
rect 14174 2554 14208 2588
rect 14174 2479 14208 2513
rect 14174 2404 14208 2438
rect 14174 2329 14208 2363
rect 14174 2254 14208 2288
rect 14174 2179 14208 2213
rect 14174 2104 14208 2138
rect 13990 1954 14024 1988
rect 14174 2029 14208 2063
rect 14266 3098 14300 3132
rect 14266 3023 14300 3057
rect 14266 2948 14300 2982
rect 14266 2873 14300 2907
rect 14266 2798 14300 2832
rect 14266 2723 14300 2757
rect 14266 2648 14300 2682
rect 14266 2572 14300 2606
rect 14266 2496 14300 2530
rect 14266 2420 14300 2454
rect 14266 2344 14300 2378
rect 14266 2268 14300 2302
rect 14266 2192 14300 2226
rect 14266 2116 14300 2150
rect 14266 2040 14300 2074
rect 14542 3300 14576 3334
rect 14542 3226 14576 3260
rect 14542 3152 14576 3186
rect 14358 3078 14392 3112
rect 14358 3004 14392 3038
rect 14358 2929 14392 2963
rect 14358 2854 14392 2888
rect 14358 2779 14392 2813
rect 14358 2704 14392 2738
rect 14358 2629 14392 2663
rect 14358 2554 14392 2588
rect 14358 2479 14392 2513
rect 14358 2404 14392 2438
rect 14358 2329 14392 2363
rect 14358 2254 14392 2288
rect 14358 2179 14392 2213
rect 14358 2104 14392 2138
rect 14174 1954 14208 1988
rect 14358 2029 14392 2063
rect 14450 3098 14484 3132
rect 14450 3023 14484 3057
rect 14450 2948 14484 2982
rect 14450 2873 14484 2907
rect 14450 2798 14484 2832
rect 14450 2723 14484 2757
rect 14450 2648 14484 2682
rect 14450 2572 14484 2606
rect 14450 2496 14484 2530
rect 14450 2420 14484 2454
rect 14450 2344 14484 2378
rect 14450 2268 14484 2302
rect 14450 2192 14484 2226
rect 14450 2116 14484 2150
rect 14450 2040 14484 2074
rect 14542 3078 14576 3112
rect 14542 3004 14576 3038
rect 14542 2929 14576 2963
rect 14542 2854 14576 2888
rect 14542 2779 14576 2813
rect 14542 2704 14576 2738
rect 14542 2629 14576 2663
rect 14542 2554 14576 2588
rect 14542 2479 14576 2513
rect 14542 2404 14576 2438
rect 14542 2329 14576 2363
rect 14542 2254 14576 2288
rect 14542 2179 14576 2213
rect 14542 2104 14576 2138
rect 14358 1954 14392 1988
rect 14542 2029 14576 2063
rect 14542 1954 14576 1988
rect 14641 3276 14675 3310
rect 14641 3208 14675 3238
rect 14641 3204 14675 3208
rect 14641 3140 14675 3166
rect 14641 3132 14675 3140
rect 14641 3072 14675 3094
rect 14641 3060 14675 3072
rect 14641 3004 14675 3022
rect 14641 2988 14675 3004
rect 14641 2936 14675 2950
rect 14641 2916 14675 2936
rect 14641 2868 14675 2877
rect 14641 2843 14675 2868
rect 14641 2800 14675 2804
rect 14641 2770 14675 2800
rect 14641 2698 14675 2731
rect 14641 2697 14675 2698
rect 14641 2630 14675 2658
rect 14641 2624 14675 2630
rect 14641 2562 14675 2585
rect 14641 2551 14675 2562
rect 14641 2494 14675 2512
rect 14641 2478 14675 2494
rect 14641 2426 14675 2439
rect 14641 2405 14675 2426
rect 14641 2358 14675 2366
rect 14641 2332 14675 2358
rect 14641 2290 14675 2293
rect 14641 2259 14675 2290
rect 14641 2188 14675 2220
rect 14641 2186 14675 2188
rect 14641 2120 14675 2147
rect 14641 2113 14675 2120
rect 14641 2052 14675 2074
rect 14641 2040 14675 2052
rect 14641 1984 14675 2001
rect 14641 1967 14675 1984
rect 13523 1890 13557 1922
rect 14641 1916 14675 1928
rect 13523 1888 13557 1890
rect 14641 1894 14675 1916
rect 13523 1822 13557 1849
rect 13523 1815 13557 1822
rect 14641 1848 14675 1855
rect 14641 1821 14675 1848
rect 13523 1754 13557 1776
rect 13523 1742 13557 1754
rect 13523 1686 13557 1703
rect 13523 1669 13557 1686
rect 13523 1618 13557 1630
rect 13523 1596 13557 1618
rect 13523 1550 13557 1557
rect 13523 1523 13557 1550
rect 13523 1482 13557 1484
rect 13523 1450 13557 1482
rect 13523 1380 13557 1411
rect 13523 1377 13557 1380
rect 13523 1312 13557 1338
rect 13523 1304 13557 1312
rect 13523 1244 13557 1266
rect 13523 1232 13557 1244
rect 13523 1176 13557 1194
rect 13523 1160 13557 1176
rect 13523 1108 13557 1122
rect 13523 1088 13557 1108
rect 13523 1040 13557 1050
rect 13523 1016 13557 1040
rect 13523 972 13557 978
rect 13523 944 13557 972
rect 13523 904 13557 906
rect 13523 872 13557 904
rect 13523 802 13557 834
rect 13523 800 13557 802
rect 13523 734 13557 762
rect 13523 728 13557 734
rect 13523 666 13557 690
rect 13523 656 13557 666
rect 13622 1770 13656 1804
rect 13622 1696 13656 1730
rect 13622 1622 13656 1656
rect 13622 1548 13656 1582
rect 13622 1474 13656 1508
rect 13622 1400 13656 1434
rect 13622 1326 13656 1360
rect 13622 1252 13656 1286
rect 13622 1178 13656 1212
rect 13622 1104 13656 1138
rect 13622 1030 13656 1064
rect 13622 956 13656 990
rect 13622 881 13656 915
rect 13622 806 13656 840
rect 13622 731 13656 765
rect 13622 656 13656 690
rect 13714 1770 13748 1804
rect 13714 1696 13748 1730
rect 13714 1622 13748 1656
rect 13714 1548 13748 1582
rect 13714 1474 13748 1508
rect 13714 1400 13748 1434
rect 13714 1326 13748 1360
rect 13714 1252 13748 1286
rect 13714 1178 13748 1212
rect 13714 1104 13748 1138
rect 13714 1030 13748 1064
rect 13714 956 13748 990
rect 13714 882 13748 916
rect 13714 808 13748 842
rect 13714 734 13748 768
rect 13714 660 13748 694
rect 13806 1770 13840 1804
rect 13806 1696 13840 1730
rect 13806 1622 13840 1656
rect 13806 1548 13840 1582
rect 13806 1474 13840 1508
rect 13806 1400 13840 1434
rect 13806 1326 13840 1360
rect 13806 1252 13840 1286
rect 13806 1178 13840 1212
rect 13806 1104 13840 1138
rect 13806 1030 13840 1064
rect 13806 956 13840 990
rect 13806 881 13840 915
rect 13806 806 13840 840
rect 13806 731 13840 765
rect 13806 656 13840 690
rect 13898 1770 13932 1804
rect 13898 1696 13932 1730
rect 13898 1622 13932 1656
rect 13898 1548 13932 1582
rect 13898 1474 13932 1508
rect 13898 1400 13932 1434
rect 13898 1326 13932 1360
rect 13898 1252 13932 1286
rect 13898 1178 13932 1212
rect 13898 1104 13932 1138
rect 13898 1030 13932 1064
rect 13898 956 13932 990
rect 13898 882 13932 916
rect 13898 808 13932 842
rect 13898 734 13932 768
rect 13898 660 13932 694
rect 13714 585 13748 619
rect 13714 510 13748 544
rect 13990 1770 14024 1804
rect 13990 1696 14024 1730
rect 13990 1622 14024 1656
rect 13990 1548 14024 1582
rect 13990 1474 14024 1508
rect 13990 1400 14024 1434
rect 13990 1326 14024 1360
rect 13990 1252 14024 1286
rect 13990 1178 14024 1212
rect 13990 1104 14024 1138
rect 13990 1030 14024 1064
rect 13990 956 14024 990
rect 13990 881 14024 915
rect 13990 806 14024 840
rect 13990 731 14024 765
rect 13990 656 14024 690
rect 14082 1770 14116 1804
rect 14082 1696 14116 1730
rect 14082 1622 14116 1656
rect 14082 1548 14116 1582
rect 14082 1474 14116 1508
rect 14082 1400 14116 1434
rect 14082 1326 14116 1360
rect 14082 1252 14116 1286
rect 14082 1178 14116 1212
rect 14082 1104 14116 1138
rect 14082 1030 14116 1064
rect 14082 956 14116 990
rect 14082 882 14116 916
rect 14082 808 14116 842
rect 14082 734 14116 768
rect 14082 660 14116 694
rect 13898 585 13932 619
rect 13898 510 13932 544
rect 14174 1770 14208 1804
rect 14174 1696 14208 1730
rect 14174 1622 14208 1656
rect 14174 1548 14208 1582
rect 14174 1474 14208 1508
rect 14174 1400 14208 1434
rect 14174 1326 14208 1360
rect 14174 1252 14208 1286
rect 14174 1178 14208 1212
rect 14174 1104 14208 1138
rect 14174 1030 14208 1064
rect 14174 956 14208 990
rect 14174 881 14208 915
rect 14174 806 14208 840
rect 14174 731 14208 765
rect 14174 656 14208 690
rect 14266 1770 14300 1804
rect 14266 1696 14300 1730
rect 14266 1622 14300 1656
rect 14266 1548 14300 1582
rect 14266 1474 14300 1508
rect 14266 1400 14300 1434
rect 14266 1326 14300 1360
rect 14266 1252 14300 1286
rect 14266 1178 14300 1212
rect 14266 1104 14300 1138
rect 14266 1030 14300 1064
rect 14266 956 14300 990
rect 14266 882 14300 916
rect 14266 808 14300 842
rect 14266 734 14300 768
rect 14266 660 14300 694
rect 14082 585 14116 619
rect 14082 510 14116 544
rect 14358 1770 14392 1804
rect 14358 1696 14392 1730
rect 14358 1622 14392 1656
rect 14358 1548 14392 1582
rect 14358 1474 14392 1508
rect 14358 1400 14392 1434
rect 14358 1326 14392 1360
rect 14358 1252 14392 1286
rect 14358 1178 14392 1212
rect 14358 1104 14392 1138
rect 14358 1030 14392 1064
rect 14358 956 14392 990
rect 14358 881 14392 915
rect 14358 806 14392 840
rect 14358 731 14392 765
rect 14358 656 14392 690
rect 14450 1770 14484 1804
rect 14450 1696 14484 1730
rect 14450 1622 14484 1656
rect 14450 1548 14484 1582
rect 14450 1474 14484 1508
rect 14450 1400 14484 1434
rect 14450 1326 14484 1360
rect 14450 1252 14484 1286
rect 14450 1178 14484 1212
rect 14450 1104 14484 1138
rect 14450 1030 14484 1064
rect 14450 956 14484 990
rect 14450 882 14484 916
rect 14450 808 14484 842
rect 14450 734 14484 768
rect 14450 660 14484 694
rect 14266 585 14300 619
rect 14266 510 14300 544
rect 14450 585 14484 619
rect 14450 510 14484 544
rect 14542 1770 14576 1804
rect 14542 1696 14576 1730
rect 14542 1622 14576 1656
rect 14542 1548 14576 1582
rect 14542 1474 14576 1508
rect 14542 1399 14576 1433
rect 14542 1324 14576 1358
rect 14542 1249 14576 1283
rect 14542 1174 14576 1208
rect 14542 1099 14576 1133
rect 14542 1024 14576 1058
rect 14542 949 14576 983
rect 14542 874 14576 908
rect 14542 799 14576 833
rect 14542 724 14576 758
rect 14542 649 14576 683
rect 14542 574 14576 608
rect 14542 499 14576 533
rect 14542 424 14576 458
rect 14641 1780 14675 1782
rect 14641 1748 14675 1780
rect 14641 1678 14675 1709
rect 14641 1675 14675 1678
rect 14641 1610 14675 1636
rect 14641 1602 14675 1610
rect 14641 1542 14675 1563
rect 14641 1529 14675 1542
rect 14641 1474 14675 1490
rect 14641 1456 14675 1474
rect 14641 1406 14675 1417
rect 14641 1383 14675 1406
rect 14641 1338 14675 1344
rect 14641 1310 14675 1338
rect 14641 1270 14675 1271
rect 14641 1237 14675 1270
rect 14641 1168 14675 1198
rect 14641 1164 14675 1168
rect 14641 1100 14675 1125
rect 14641 1091 14675 1100
rect 14641 1032 14675 1052
rect 14641 1018 14675 1032
rect 14641 964 14675 979
rect 14641 945 14675 964
rect 14641 896 14675 906
rect 14641 872 14675 896
rect 14641 828 14675 833
rect 14641 799 14675 828
rect 14641 726 14675 760
rect 14641 658 14675 687
rect 14641 653 14675 658
rect 14641 590 14675 614
rect 14641 580 14675 590
rect 14641 522 14675 541
rect 14641 507 14675 522
rect 14641 454 14675 468
rect 14641 434 14675 454
rect 14641 386 14675 395
rect 1750 306 1781 322
rect 1781 306 1784 322
rect 1823 306 1851 322
rect 1851 306 1857 322
rect 1896 306 1921 322
rect 1921 306 1930 322
rect 1969 306 1991 322
rect 1991 306 2003 322
rect 2042 306 2061 322
rect 2061 306 2076 322
rect 2115 306 2131 322
rect 2131 306 2149 322
rect 2188 306 2201 322
rect 2201 306 2222 322
rect 2261 306 2271 322
rect 2271 306 2295 322
rect 2334 306 2341 322
rect 2341 306 2368 322
rect 2407 306 2411 322
rect 2411 306 2441 322
rect 2480 306 2481 322
rect 2481 306 2514 322
rect 1750 288 1784 306
rect 1823 288 1857 306
rect 1896 288 1930 306
rect 1969 288 2003 306
rect 2042 288 2076 306
rect 2115 288 2149 306
rect 2188 288 2222 306
rect 2261 288 2295 306
rect 2334 288 2368 306
rect 2407 288 2441 306
rect 2480 288 2514 306
rect 2553 288 2587 322
rect 2626 306 2657 322
rect 2657 306 2660 322
rect 2699 306 2727 322
rect 2727 306 2733 322
rect 2772 306 2797 322
rect 2797 306 2806 322
rect 2845 306 2867 322
rect 2867 306 2879 322
rect 2918 306 2937 322
rect 2937 306 2952 322
rect 2991 306 3007 322
rect 3007 306 3025 322
rect 3064 306 3077 322
rect 3077 306 3098 322
rect 3137 306 3147 322
rect 3147 306 3171 322
rect 3210 306 3217 322
rect 3217 306 3244 322
rect 2626 288 2660 306
rect 2699 288 2733 306
rect 2772 288 2806 306
rect 2845 288 2879 306
rect 2918 288 2952 306
rect 2991 288 3025 306
rect 3064 288 3098 306
rect 3137 288 3171 306
rect 3210 288 3244 306
rect 13340 241 13446 347
rect 13679 334 13683 368
rect 13683 334 13713 368
rect 13753 334 13756 368
rect 13756 334 13787 368
rect 13827 334 13829 368
rect 13829 334 13861 368
rect 13901 334 13902 368
rect 13902 334 13935 368
rect 13974 334 13975 368
rect 13975 334 14008 368
rect 14047 334 14048 368
rect 14048 334 14081 368
rect 14120 334 14121 368
rect 14121 334 14154 368
rect 14193 334 14227 368
rect 14266 334 14299 368
rect 14299 334 14300 368
rect 14339 334 14371 368
rect 14371 334 14373 368
rect 14412 334 14443 368
rect 14443 334 14446 368
rect 14485 334 14515 368
rect 14515 334 14519 368
rect 14641 361 14675 386
rect 14641 318 14675 322
rect 14641 288 14675 318
rect 13522 216 13556 250
rect 13597 216 13625 250
rect 13625 216 13631 250
rect 13672 216 13693 250
rect 13693 216 13706 250
rect 13747 216 13761 250
rect 13761 216 13781 250
rect 13822 216 13829 250
rect 13829 216 13856 250
rect 13897 216 13931 250
rect 13972 216 13999 250
rect 13999 216 14006 250
rect 14047 216 14067 250
rect 14067 216 14081 250
rect 14122 216 14135 250
rect 14135 216 14156 250
rect 14197 216 14203 250
rect 14203 216 14231 250
rect 14271 216 14305 250
rect 14345 216 14373 250
rect 14373 216 14379 250
rect 14419 216 14441 250
rect 14441 216 14453 250
rect 14493 216 14509 250
rect 14509 216 14527 250
rect 14567 216 14577 250
rect 14577 216 14601 250
<< metal1 >>
rect 13982 39556 14957 39568
rect 13982 39522 14775 39556
rect 14809 39522 14917 39556
rect 14951 39522 14957 39556
rect 1938 39476 13950 39482
rect 1938 39470 2163 39476
tri 1590 39284 1602 39296 se
rect 1602 39284 1734 39296
tri 1556 39250 1590 39284 se
rect 1590 39250 1684 39284
rect 1718 39250 1734 39284
tri 1520 39214 1556 39250 se
rect 1556 39214 1734 39250
rect 1520 39212 1734 39214
rect 1520 39178 1684 39212
rect 1718 39178 1734 39212
rect 1520 39166 1734 39178
rect 1520 28568 1638 39166
tri 1638 39106 1698 39166 nw
rect 1938 34108 1944 39470
rect 2050 39370 2163 39470
rect 10189 39442 10228 39476
rect 10262 39442 10301 39476
rect 10335 39442 10374 39476
rect 10408 39442 10447 39476
rect 10481 39442 10520 39476
rect 10554 39442 10593 39476
rect 10627 39442 10666 39476
rect 10700 39442 10739 39476
rect 10773 39442 10812 39476
rect 10846 39442 10885 39476
rect 10919 39442 10958 39476
rect 10992 39442 11031 39476
rect 11065 39442 11104 39476
rect 11138 39442 11177 39476
rect 11211 39442 11250 39476
rect 11284 39442 11323 39476
rect 11357 39442 11396 39476
rect 11430 39442 11469 39476
rect 11503 39442 11542 39476
rect 11576 39442 11615 39476
rect 11649 39442 11688 39476
rect 11722 39442 11761 39476
rect 11795 39442 11834 39476
rect 11868 39442 11907 39476
rect 11941 39442 11980 39476
rect 12014 39442 12053 39476
rect 12087 39442 12126 39476
rect 12160 39442 12199 39476
rect 12233 39442 12272 39476
rect 12306 39442 12345 39476
rect 12379 39442 12418 39476
rect 12452 39442 12491 39476
rect 12525 39442 12564 39476
rect 12598 39442 12637 39476
rect 12671 39442 12710 39476
rect 12744 39442 12783 39476
rect 12817 39442 12856 39476
rect 12890 39442 12929 39476
rect 12963 39442 13002 39476
rect 13036 39442 13075 39476
rect 13109 39442 13148 39476
rect 13182 39442 13221 39476
rect 13255 39442 13294 39476
rect 13328 39442 13367 39476
rect 13401 39442 13440 39476
rect 13474 39442 13513 39476
rect 13547 39442 13586 39476
rect 13620 39442 13659 39476
rect 13693 39442 13732 39476
rect 13766 39470 13950 39476
rect 13766 39442 13838 39470
rect 10189 39404 13838 39442
rect 10189 39370 10228 39404
rect 10262 39370 10301 39404
rect 10335 39370 10374 39404
rect 10408 39370 10447 39404
rect 10481 39370 10520 39404
rect 10554 39370 10593 39404
rect 10627 39370 10666 39404
rect 10700 39370 10739 39404
rect 10773 39370 10812 39404
rect 10846 39370 10885 39404
rect 10919 39370 10958 39404
rect 10992 39370 11031 39404
rect 11065 39370 11104 39404
rect 11138 39370 11177 39404
rect 11211 39370 11250 39404
rect 11284 39370 11323 39404
rect 11357 39370 11396 39404
rect 11430 39370 11469 39404
rect 11503 39370 11542 39404
rect 11576 39370 11615 39404
rect 11649 39370 11688 39404
rect 11722 39370 11761 39404
rect 11795 39370 11834 39404
rect 11868 39370 11907 39404
rect 11941 39370 11980 39404
rect 12014 39370 12053 39404
rect 12087 39370 12126 39404
rect 12160 39370 12199 39404
rect 12233 39370 12272 39404
rect 12306 39370 12345 39404
rect 12379 39370 12418 39404
rect 12452 39370 12491 39404
rect 12525 39370 12564 39404
rect 12598 39370 12637 39404
rect 12671 39370 12710 39404
rect 12744 39370 12783 39404
rect 12817 39370 12856 39404
rect 12890 39370 12929 39404
rect 12963 39370 13002 39404
rect 13036 39370 13075 39404
rect 13109 39370 13148 39404
rect 13182 39370 13221 39404
rect 13255 39370 13294 39404
rect 13328 39370 13367 39404
rect 13401 39370 13440 39404
rect 13474 39370 13513 39404
rect 13547 39370 13586 39404
rect 13620 39370 13659 39404
rect 13693 39370 13732 39404
rect 13766 39370 13838 39404
rect 2050 39364 13838 39370
rect 2050 34108 2056 39364
tri 2056 39330 2090 39364 nw
tri 13798 39330 13832 39364 ne
rect 1938 34069 2056 34108
rect 1938 34035 1944 34069
rect 1978 34035 2016 34069
rect 2050 34035 2056 34069
rect 1938 33996 2056 34035
rect 1938 33962 1944 33996
rect 1978 33962 2016 33996
rect 2050 33962 2056 33996
rect 1938 33923 2056 33962
rect 1938 33889 1944 33923
rect 1978 33889 2016 33923
rect 2050 33889 2056 33923
rect 1938 33850 2056 33889
rect 1938 33816 1944 33850
rect 1978 33816 2016 33850
rect 2050 33816 2056 33850
rect 1938 33777 2056 33816
rect 1938 33743 1944 33777
rect 1978 33743 2016 33777
rect 2050 33743 2056 33777
rect 1938 33704 2056 33743
rect 1938 33670 1944 33704
rect 1978 33670 2016 33704
rect 2050 33670 2056 33704
tri 1914 33537 1938 33561 se
rect 1938 33537 2056 33670
tri 1875 33498 1914 33537 se
rect 1914 33513 2056 33537
rect 1914 33498 2041 33513
tri 2041 33498 2056 33513 nw
rect 2213 39171 13705 39177
rect 2213 39099 2291 39171
rect 2213 39065 2219 39099
rect 2253 39065 2291 39099
rect 9957 39137 9996 39171
rect 10030 39137 10069 39171
rect 10103 39137 10142 39171
rect 10176 39137 10215 39171
rect 10249 39137 10288 39171
rect 10322 39137 10361 39171
rect 10395 39137 10434 39171
rect 10468 39137 10507 39171
rect 10541 39137 10580 39171
rect 10614 39137 10653 39171
rect 10687 39137 10726 39171
rect 10760 39137 10799 39171
rect 10833 39137 10872 39171
rect 10906 39137 10945 39171
rect 10979 39137 11018 39171
rect 11052 39137 11091 39171
rect 11125 39137 11164 39171
rect 11198 39137 11237 39171
rect 11271 39137 11310 39171
rect 11344 39137 11383 39171
rect 11417 39137 11456 39171
rect 11490 39137 11529 39171
rect 11563 39137 11602 39171
rect 11636 39137 11675 39171
rect 11709 39137 11748 39171
rect 11782 39137 11821 39171
rect 11855 39137 11894 39171
rect 11928 39137 11967 39171
rect 12001 39137 12040 39171
rect 12074 39137 12113 39171
rect 12147 39137 12186 39171
rect 12220 39137 12259 39171
rect 12293 39137 12332 39171
rect 12366 39137 12405 39171
rect 12439 39137 12478 39171
rect 12512 39137 12551 39171
rect 12585 39137 12624 39171
rect 12658 39137 12697 39171
rect 12731 39137 12770 39171
rect 12804 39137 12843 39171
rect 12877 39137 12916 39171
rect 12950 39137 12989 39171
rect 9957 39099 12989 39137
rect 9957 39065 9996 39099
rect 10030 39065 10069 39099
rect 10103 39065 10142 39099
rect 10176 39065 10215 39099
rect 10249 39065 10288 39099
rect 10322 39065 10361 39099
rect 10395 39065 10434 39099
rect 10468 39065 10507 39099
rect 10541 39065 10580 39099
rect 10614 39065 10653 39099
rect 10687 39065 10726 39099
rect 10760 39065 10799 39099
rect 10833 39065 10872 39099
rect 10906 39065 10945 39099
rect 10979 39065 11018 39099
rect 11052 39065 11091 39099
rect 11125 39065 11164 39099
rect 11198 39065 11237 39099
rect 11271 39065 11310 39099
rect 11344 39065 11383 39099
rect 11417 39065 11456 39099
rect 11490 39065 11529 39099
rect 11563 39065 11602 39099
rect 11636 39065 11675 39099
rect 11709 39065 11748 39099
rect 11782 39065 11821 39099
rect 11855 39065 11894 39099
rect 11928 39065 11967 39099
rect 12001 39065 12040 39099
rect 12074 39065 12113 39099
rect 12147 39065 12186 39099
rect 12220 39065 12259 39099
rect 12293 39065 12332 39099
rect 12366 39065 12405 39099
rect 12439 39065 12478 39099
rect 12512 39065 12551 39099
rect 12585 39065 12624 39099
rect 12658 39065 12697 39099
rect 12731 39065 12770 39099
rect 12804 39065 12843 39099
rect 12877 39065 12916 39099
rect 12950 39065 12989 39099
rect 2213 39026 2363 39065
rect 2213 38992 2219 39026
rect 2253 38992 2291 39026
rect 2325 38993 2363 39026
rect 9957 39027 12989 39065
rect 9957 38993 9996 39027
rect 10030 38993 10069 39027
rect 10103 38993 10142 39027
rect 10176 38993 10215 39027
rect 10249 38993 10288 39027
rect 10322 38993 10361 39027
rect 10395 38993 10434 39027
rect 10468 38993 10507 39027
rect 10541 38993 10580 39027
rect 10614 38993 10653 39027
rect 10687 38993 10726 39027
rect 10760 38993 10799 39027
rect 10833 38993 10872 39027
rect 10906 38993 10945 39027
rect 10979 38993 11018 39027
rect 11052 38993 11091 39027
rect 11125 38993 11164 39027
rect 11198 38993 11237 39027
rect 11271 38993 11310 39027
rect 11344 38993 11383 39027
rect 11417 38993 11456 39027
rect 11490 38993 11529 39027
rect 11563 38993 11602 39027
rect 11636 38993 11675 39027
rect 11709 38993 11748 39027
rect 11782 38993 11821 39027
rect 11855 38993 11894 39027
rect 11928 38993 11967 39027
rect 12001 38993 12040 39027
rect 12074 38993 12113 39027
rect 12147 38993 12186 39027
rect 12220 38993 12259 39027
rect 12293 38993 12332 39027
rect 12366 38993 12405 39027
rect 12439 38993 12478 39027
rect 12512 38993 12551 39027
rect 12585 38993 12624 39027
rect 12658 38993 12697 39027
rect 12731 38993 12770 39027
rect 12804 38993 12843 39027
rect 12877 38993 12916 39027
rect 12950 38993 12989 39027
rect 13095 39137 13137 39171
rect 13171 39137 13213 39171
rect 13247 39137 13289 39171
rect 13323 39137 13365 39171
rect 13399 39137 13441 39171
rect 13475 39137 13517 39171
rect 13551 39137 13593 39171
rect 13627 39137 13705 39171
rect 13095 39099 13705 39137
rect 13095 39065 13137 39099
rect 13171 39065 13213 39099
rect 13247 39065 13289 39099
rect 13323 39065 13365 39099
rect 13399 39065 13441 39099
rect 13475 39065 13517 39099
rect 13551 39065 13593 39099
rect 13095 39027 13593 39065
rect 13095 38993 13137 39027
rect 13171 38993 13213 39027
rect 13247 38993 13290 39027
rect 13324 38993 13367 39027
rect 13401 38993 13444 39027
rect 13478 38993 13521 39027
rect 2325 38992 13521 38993
rect 2213 38987 13521 38992
rect 2213 38954 2403 38987
rect 2213 38953 2363 38954
rect 2213 38919 2219 38953
rect 2253 38919 2291 38953
rect 2325 38920 2363 38953
rect 2397 38920 2403 38954
tri 2403 38953 2437 38987 nw
tri 13481 38953 13515 38987 ne
rect 2325 38919 2403 38920
rect 2213 38881 2403 38919
rect 2213 38880 2363 38881
rect 2213 38846 2219 38880
rect 2253 38846 2291 38880
rect 2325 38847 2363 38880
rect 2397 38847 2403 38881
rect 2325 38846 2403 38847
rect 2213 38808 2403 38846
rect 2213 38807 2363 38808
rect 2213 38773 2219 38807
rect 2253 38773 2291 38807
rect 2325 38774 2363 38807
rect 2397 38774 2403 38808
rect 2325 38773 2403 38774
rect 2213 38735 2403 38773
rect 2213 38734 2363 38735
rect 2213 38700 2219 38734
rect 2253 38720 2291 38734
rect 2325 38720 2363 38734
rect 2397 38701 2403 38735
rect 2213 38668 2249 38700
rect 2301 38668 2315 38700
rect 2367 38668 2403 38701
rect 2213 38662 2403 38668
rect 2213 38661 2363 38662
rect 2213 38627 2219 38661
rect 2253 38656 2291 38661
rect 2325 38656 2363 38661
rect 2397 38628 2403 38662
rect 2213 38604 2249 38627
rect 2301 38604 2315 38627
rect 2367 38604 2403 38628
rect 2213 38592 2403 38604
rect 2213 38588 2249 38592
rect 2301 38588 2315 38592
rect 2367 38589 2403 38592
rect 2213 38554 2219 38588
rect 2397 38555 2403 38589
rect 2213 38540 2249 38554
rect 2301 38540 2315 38554
rect 2367 38540 2403 38555
rect 2213 38528 2403 38540
rect 2213 38515 2249 38528
rect 2301 38515 2315 38528
rect 2367 38516 2403 38528
rect 2213 38481 2219 38515
rect 2397 38482 2403 38516
rect 2213 38476 2249 38481
rect 2301 38476 2315 38481
rect 2367 38476 2403 38482
rect 2213 38464 2403 38476
rect 2213 38442 2249 38464
rect 2301 38442 2315 38464
rect 2367 38443 2403 38464
rect 2213 38408 2219 38442
rect 2253 38408 2291 38412
rect 2325 38409 2363 38412
rect 2397 38409 2403 38443
rect 2325 38408 2403 38409
rect 2213 38400 2403 38408
rect 2213 38369 2249 38400
rect 2301 38369 2315 38400
rect 2367 38370 2403 38400
rect 2213 38335 2219 38369
rect 2253 38336 2291 38348
rect 2325 38336 2363 38348
rect 2397 38336 2403 38370
rect 2213 38296 2249 38335
rect 2301 38296 2315 38335
rect 2367 38297 2403 38336
rect 2213 38262 2219 38296
rect 2253 38272 2291 38284
rect 2325 38272 2363 38284
rect 2397 38263 2403 38297
rect 2213 38223 2249 38262
rect 2301 38223 2315 38262
rect 2367 38224 2403 38263
rect 2213 38189 2219 38223
rect 2253 38208 2291 38220
rect 2325 38208 2363 38220
rect 2397 38190 2403 38224
rect 2213 38156 2249 38189
rect 2301 38156 2315 38189
rect 2367 38156 2403 38190
rect 2213 38151 2403 38156
rect 2213 38150 2363 38151
rect 2213 38116 2219 38150
rect 2253 38144 2291 38150
rect 2325 38144 2363 38150
rect 2397 38117 2403 38151
rect 2213 38092 2249 38116
rect 2301 38092 2315 38116
rect 2367 38092 2403 38117
rect 2213 38080 2403 38092
rect 2213 38077 2249 38080
rect 2301 38077 2315 38080
rect 2367 38078 2403 38080
rect 2213 38043 2219 38077
rect 2397 38044 2403 38078
rect 2213 38028 2249 38043
rect 2301 38028 2315 38043
rect 2367 38028 2403 38044
rect 2213 38016 2403 38028
rect 2213 38004 2249 38016
rect 2301 38004 2315 38016
rect 2367 38005 2403 38016
rect 2213 37970 2219 38004
rect 2397 37971 2403 38005
rect 2213 37964 2249 37970
rect 2301 37964 2315 37970
rect 2367 37964 2403 37971
rect 2213 37952 2403 37964
rect 2213 37931 2249 37952
rect 2301 37931 2315 37952
rect 2367 37932 2403 37952
rect 2213 37897 2219 37931
rect 2253 37897 2291 37900
rect 2325 37898 2363 37900
rect 2397 37898 2403 37932
rect 2325 37897 2403 37898
rect 2213 37888 2403 37897
rect 2213 37858 2249 37888
rect 2301 37858 2315 37888
rect 2367 37859 2403 37888
rect 2213 37824 2219 37858
rect 2253 37824 2291 37836
rect 2325 37825 2363 37836
rect 2397 37825 2403 37859
rect 2325 37824 2403 37825
rect 2213 37785 2249 37824
rect 2301 37785 2315 37824
rect 2367 37786 2403 37824
rect 2213 37751 2219 37785
rect 2253 37760 2291 37772
rect 2325 37760 2363 37772
rect 2397 37752 2403 37786
rect 2213 37712 2249 37751
rect 2301 37712 2315 37751
rect 2367 37713 2403 37752
rect 2213 37678 2219 37712
rect 2253 37696 2291 37708
rect 2325 37696 2363 37708
rect 2397 37679 2403 37713
rect 2213 37644 2249 37678
rect 2301 37644 2315 37678
rect 2367 37644 2403 37679
rect 2213 37640 2403 37644
rect 2213 37639 2363 37640
rect 2213 37605 2219 37639
rect 2253 37632 2291 37639
rect 2325 37632 2363 37639
rect 2397 37606 2403 37640
rect 2213 37580 2249 37605
rect 2301 37580 2315 37605
rect 2367 37580 2403 37606
rect 2213 37568 2403 37580
rect 2213 37566 2249 37568
rect 2301 37566 2315 37568
rect 2367 37567 2403 37568
rect 2213 37532 2219 37566
rect 2397 37533 2403 37567
rect 2213 37516 2249 37532
rect 2301 37516 2315 37532
rect 2367 37516 2403 37533
rect 2213 37504 2403 37516
rect 2213 37493 2249 37504
rect 2301 37493 2315 37504
rect 2367 37494 2403 37504
rect 2213 37459 2219 37493
rect 2397 37460 2403 37494
rect 2213 37452 2249 37459
rect 2301 37452 2315 37459
rect 2367 37452 2403 37460
rect 2213 37440 2403 37452
rect 2213 37420 2249 37440
rect 2301 37420 2315 37440
rect 2367 37421 2403 37440
rect 2213 37386 2219 37420
rect 2253 37386 2291 37388
rect 2325 37387 2363 37388
rect 2397 37387 2403 37421
rect 2325 37386 2403 37387
rect 2213 37376 2403 37386
rect 2213 37347 2249 37376
rect 2301 37347 2315 37376
rect 2367 37348 2403 37376
rect 2213 37313 2219 37347
rect 2253 37313 2291 37324
rect 2325 37314 2363 37324
rect 2397 37314 2403 37348
rect 2325 37313 2403 37314
rect 2213 37312 2403 37313
rect 2213 37274 2249 37312
rect 2301 37274 2315 37312
rect 2367 37275 2403 37312
rect 2213 37240 2219 37274
rect 2253 37248 2291 37260
rect 2325 37248 2363 37260
rect 2397 37241 2403 37275
rect 2213 37201 2249 37240
rect 2301 37201 2315 37240
rect 2367 37202 2403 37241
rect 2213 37167 2219 37201
rect 2253 37184 2291 37196
rect 2325 37184 2363 37196
rect 2397 37168 2403 37202
rect 2213 37132 2249 37167
rect 2301 37132 2315 37167
rect 2367 37132 2403 37168
rect 2213 37129 2403 37132
rect 2213 37128 2363 37129
rect 2213 37094 2219 37128
rect 2253 37120 2291 37128
rect 2325 37120 2363 37128
rect 2397 37095 2403 37129
rect 2213 37068 2249 37094
rect 2301 37068 2315 37094
rect 2367 37068 2403 37095
rect 2213 37056 2403 37068
rect 2213 37055 2249 37056
rect 2301 37055 2315 37056
rect 2213 37021 2219 37055
rect 2397 37022 2403 37056
rect 2213 37004 2249 37021
rect 2301 37004 2315 37021
rect 2367 37004 2403 37022
rect 2213 36992 2403 37004
rect 2213 36982 2249 36992
rect 2301 36982 2315 36992
rect 2367 36983 2403 36992
rect 2213 36948 2219 36982
rect 2397 36949 2403 36983
rect 2213 36940 2249 36948
rect 2301 36940 2315 36948
rect 2367 36940 2403 36949
rect 2213 36928 2403 36940
rect 2213 36909 2249 36928
rect 2301 36909 2315 36928
rect 2367 36910 2403 36928
rect 2213 36875 2219 36909
rect 2397 36876 2403 36910
rect 2253 36875 2291 36876
rect 2325 36875 2403 36876
rect 2213 36864 2403 36875
rect 2213 36836 2249 36864
rect 2301 36836 2315 36864
rect 2367 36837 2403 36864
rect 2213 36802 2219 36836
rect 2253 36802 2291 36812
rect 2325 36803 2363 36812
rect 2397 36803 2403 36837
rect 2325 36802 2403 36803
rect 2213 36800 2403 36802
rect 2213 36763 2249 36800
rect 2301 36763 2315 36800
rect 2367 36764 2403 36800
rect 2213 36729 2219 36763
rect 2253 36736 2291 36748
rect 2325 36736 2363 36748
rect 2397 36730 2403 36764
rect 2213 36690 2249 36729
rect 2301 36690 2315 36729
rect 2367 36691 2403 36730
rect 2475 38834 2878 38886
rect 2930 38834 2943 38886
rect 2995 38834 3008 38886
rect 3060 38854 3073 38886
rect 3125 38854 3138 38886
rect 3190 38854 3203 38886
rect 3255 38854 3268 38886
rect 3320 38854 3332 38886
rect 3384 38854 3396 38886
rect 3064 38834 3073 38854
rect 3137 38834 3138 38854
rect 3320 38834 3322 38854
rect 3384 38834 3395 38854
rect 3448 38834 3460 38886
rect 3512 38834 3524 38886
rect 3576 38834 3588 38886
rect 3640 38854 3652 38886
rect 3704 38854 3716 38886
rect 3768 38854 3780 38886
rect 3832 38854 3844 38886
rect 3896 38854 3908 38886
rect 3648 38834 3652 38854
rect 3832 38834 3833 38854
rect 3896 38834 3906 38854
rect 3960 38834 3972 38886
rect 4024 38834 4036 38886
rect 4088 38834 4100 38886
rect 4152 38854 4164 38886
rect 4216 38854 4228 38886
rect 4280 38854 4292 38886
rect 4344 38854 4356 38886
rect 4408 38854 4420 38886
rect 4159 38834 4164 38854
rect 4408 38834 4417 38854
rect 4472 38834 4484 38886
rect 4536 38834 4548 38886
rect 4600 38834 4612 38886
rect 4664 38854 4676 38886
rect 4728 38854 4740 38886
rect 4792 38854 4804 38886
rect 4856 38854 4868 38886
rect 4920 38854 4932 38886
rect 4670 38834 4676 38854
rect 4920 38834 4928 38854
rect 4984 38834 4996 38886
rect 5048 38834 5060 38886
rect 5112 38834 5124 38886
rect 5176 38854 5188 38886
rect 5240 38854 5252 38886
rect 5304 38854 5316 38886
rect 5368 38854 5380 38886
rect 5432 38854 5444 38886
rect 5181 38834 5188 38854
rect 5432 38834 5439 38854
rect 5496 38834 5508 38886
rect 5560 38834 5572 38886
rect 5624 38834 5636 38886
rect 5688 38854 5700 38886
rect 5752 38854 5764 38886
rect 5816 38854 5828 38886
rect 5880 38854 5892 38886
rect 5944 38854 5956 38886
rect 6008 38854 6020 38886
rect 5690 38834 5700 38854
rect 5762 38834 5764 38854
rect 6008 38834 6016 38854
rect 6072 38834 6084 38886
rect 6136 38834 6148 38886
rect 6200 38834 6212 38886
rect 6264 38854 6276 38886
rect 6328 38854 6340 38886
rect 6392 38854 6404 38886
rect 6456 38854 6468 38886
rect 6520 38854 6532 38886
rect 6584 38854 6596 38886
rect 6266 38834 6276 38854
rect 6338 38834 6340 38854
rect 6584 38834 6592 38854
rect 6648 38834 6660 38886
rect 6712 38834 6724 38886
rect 6776 38834 6788 38886
rect 6840 38854 6852 38886
rect 6904 38854 6916 38886
rect 6968 38854 6980 38886
rect 7032 38854 7044 38886
rect 7096 38854 7108 38886
rect 7160 38854 7172 38886
rect 6842 38834 6852 38854
rect 6914 38834 6916 38854
rect 7160 38834 7168 38854
rect 7224 38834 7236 38886
rect 7288 38834 7300 38886
rect 7352 38834 7364 38886
rect 7416 38854 7428 38886
rect 7480 38854 7492 38886
rect 7544 38854 7556 38886
rect 7608 38854 7620 38886
rect 7672 38854 7684 38886
rect 7736 38854 7748 38886
rect 7418 38834 7428 38854
rect 7490 38834 7492 38854
rect 7736 38834 7744 38854
rect 7800 38834 7812 38886
rect 7864 38834 7876 38886
rect 7928 38834 7940 38886
rect 7992 38854 8004 38886
rect 8056 38854 8068 38886
rect 8120 38854 8132 38886
rect 8184 38854 8196 38886
rect 8248 38854 8260 38886
rect 8312 38854 8324 38886
rect 7994 38834 8004 38854
rect 8066 38834 8068 38854
rect 8312 38834 8320 38854
rect 8376 38834 8388 38886
rect 8440 38834 8452 38886
rect 8504 38834 8516 38886
rect 8568 38854 8580 38886
rect 8632 38854 8644 38886
rect 8696 38854 8708 38886
rect 8760 38854 8772 38886
rect 8824 38854 8836 38886
rect 8888 38854 8900 38886
rect 8570 38834 8580 38854
rect 8642 38834 8644 38854
rect 8888 38834 8896 38854
rect 8952 38834 8964 38886
rect 9016 38834 9028 38886
rect 9080 38834 9092 38886
rect 9144 38854 9156 38886
rect 9208 38854 9220 38886
rect 9272 38854 9284 38886
rect 9336 38854 9348 38886
rect 9400 38854 9412 38886
rect 9464 38854 9476 38886
rect 9146 38834 9156 38854
rect 9218 38834 9220 38854
rect 9464 38834 9472 38854
rect 9528 38834 9540 38886
rect 9592 38834 9604 38886
rect 9656 38834 9668 38886
rect 9720 38854 9732 38886
rect 9784 38854 9796 38886
rect 9848 38854 9860 38886
rect 9912 38854 9924 38886
rect 9976 38854 9988 38886
rect 10040 38854 10052 38886
rect 9722 38834 9732 38854
rect 9794 38834 9796 38854
rect 10040 38834 10048 38854
rect 10104 38834 10116 38886
rect 10168 38834 10180 38886
rect 10232 38834 10244 38886
rect 10296 38854 10308 38886
rect 10360 38854 10372 38886
rect 10424 38854 10436 38886
rect 10488 38854 10500 38886
rect 10552 38854 10564 38886
rect 10616 38854 10628 38886
rect 10298 38834 10308 38854
rect 10370 38834 10372 38854
rect 10616 38834 10624 38854
rect 10680 38834 10692 38886
rect 10744 38834 10756 38886
rect 10808 38834 10820 38886
rect 10872 38854 10884 38886
rect 10936 38854 10948 38886
rect 11000 38854 11012 38886
rect 11064 38854 11076 38886
rect 11128 38854 11140 38886
rect 11192 38854 11204 38886
rect 10874 38834 10884 38854
rect 10946 38834 10948 38854
rect 11192 38834 11200 38854
rect 11256 38834 11268 38886
rect 11320 38834 11332 38886
rect 11384 38834 11396 38886
rect 11448 38854 11460 38886
rect 11512 38854 11524 38886
rect 11576 38854 11588 38886
rect 11640 38854 11652 38886
rect 11704 38854 11716 38886
rect 11768 38854 11780 38886
rect 11450 38834 11460 38854
rect 11522 38834 11524 38854
rect 11768 38834 11776 38854
rect 11832 38834 11844 38886
rect 11896 38834 11908 38886
rect 11960 38834 11972 38886
rect 12024 38854 12036 38886
rect 12088 38854 12100 38886
rect 12152 38854 12164 38886
rect 12216 38854 12228 38886
rect 12280 38854 12292 38886
rect 12344 38854 12356 38886
rect 12026 38834 12036 38854
rect 12098 38834 12100 38854
rect 12344 38834 12352 38854
rect 12408 38834 12420 38886
rect 12472 38834 12484 38886
rect 12536 38834 12548 38886
rect 12600 38854 12612 38886
rect 12664 38854 12676 38886
rect 12728 38854 12740 38886
rect 12792 38854 12804 38886
rect 12856 38854 12868 38886
rect 12920 38854 12932 38886
rect 12602 38834 12612 38854
rect 12674 38834 12676 38854
rect 12920 38834 12928 38854
rect 12984 38834 12996 38886
rect 13048 38834 13060 38886
rect 13112 38834 13118 38886
rect 2475 38820 2884 38834
rect 2918 38820 2957 38834
rect 2991 38820 3030 38834
rect 3064 38820 3103 38834
rect 3137 38820 3176 38834
rect 3210 38820 3249 38834
rect 3283 38820 3322 38834
rect 3356 38820 3395 38834
rect 3429 38820 3468 38834
rect 3502 38820 3541 38834
rect 3575 38820 3614 38834
rect 3648 38820 3687 38834
rect 3721 38820 3760 38834
rect 3794 38820 3833 38834
rect 3867 38820 3906 38834
rect 3940 38820 3979 38834
rect 4013 38820 4052 38834
rect 4086 38820 4125 38834
rect 4159 38820 4198 38834
rect 4232 38820 4271 38834
rect 4305 38820 4344 38834
rect 4378 38820 4417 38834
rect 4451 38820 4490 38834
rect 4524 38820 4563 38834
rect 4597 38820 4636 38834
rect 4670 38820 4709 38834
rect 4743 38820 4782 38834
rect 4816 38820 4855 38834
rect 4889 38820 4928 38834
rect 4962 38820 5001 38834
rect 5035 38820 5074 38834
rect 5108 38820 5147 38834
rect 5181 38820 5220 38834
rect 5254 38820 5293 38834
rect 5327 38820 5366 38834
rect 5400 38820 5439 38834
rect 5473 38820 5512 38834
rect 5546 38820 5584 38834
rect 5618 38820 5656 38834
rect 5690 38820 5728 38834
rect 5762 38820 5800 38834
rect 5834 38820 5872 38834
rect 5906 38820 5944 38834
rect 5978 38820 6016 38834
rect 6050 38820 6088 38834
rect 6122 38820 6160 38834
rect 6194 38820 6232 38834
rect 6266 38820 6304 38834
rect 6338 38820 6376 38834
rect 6410 38820 6448 38834
rect 6482 38820 6520 38834
rect 6554 38820 6592 38834
rect 6626 38820 6664 38834
rect 6698 38820 6736 38834
rect 6770 38820 6808 38834
rect 6842 38820 6880 38834
rect 6914 38820 6952 38834
rect 6986 38820 7024 38834
rect 7058 38820 7096 38834
rect 7130 38820 7168 38834
rect 7202 38820 7240 38834
rect 7274 38820 7312 38834
rect 7346 38820 7384 38834
rect 7418 38820 7456 38834
rect 7490 38820 7528 38834
rect 7562 38820 7600 38834
rect 7634 38820 7672 38834
rect 7706 38820 7744 38834
rect 7778 38820 7816 38834
rect 7850 38820 7888 38834
rect 7922 38820 7960 38834
rect 7994 38820 8032 38834
rect 8066 38820 8104 38834
rect 8138 38820 8176 38834
rect 8210 38820 8248 38834
rect 8282 38820 8320 38834
rect 8354 38820 8392 38834
rect 8426 38820 8464 38834
rect 8498 38820 8536 38834
rect 8570 38820 8608 38834
rect 8642 38820 8680 38834
rect 8714 38820 8752 38834
rect 8786 38820 8824 38834
rect 8858 38820 8896 38834
rect 8930 38820 8968 38834
rect 9002 38820 9040 38834
rect 9074 38820 9112 38834
rect 9146 38820 9184 38834
rect 9218 38820 9256 38834
rect 9290 38820 9328 38834
rect 9362 38820 9400 38834
rect 9434 38820 9472 38834
rect 9506 38820 9544 38834
rect 9578 38820 9616 38834
rect 9650 38820 9688 38834
rect 9722 38820 9760 38834
rect 9794 38820 9832 38834
rect 9866 38820 9904 38834
rect 9938 38820 9976 38834
rect 10010 38820 10048 38834
rect 10082 38820 10120 38834
rect 10154 38820 10192 38834
rect 10226 38820 10264 38834
rect 10298 38820 10336 38834
rect 10370 38820 10408 38834
rect 10442 38820 10480 38834
rect 10514 38820 10552 38834
rect 10586 38820 10624 38834
rect 10658 38820 10696 38834
rect 10730 38820 10768 38834
rect 10802 38820 10840 38834
rect 10874 38820 10912 38834
rect 10946 38820 10984 38834
rect 11018 38820 11056 38834
rect 11090 38820 11128 38834
rect 11162 38820 11200 38834
rect 11234 38820 11272 38834
rect 11306 38820 11344 38834
rect 11378 38820 11416 38834
rect 11450 38820 11488 38834
rect 11522 38820 11560 38834
rect 11594 38820 11632 38834
rect 11666 38820 11704 38834
rect 11738 38820 11776 38834
rect 11810 38820 11848 38834
rect 11882 38820 11920 38834
rect 11954 38820 11992 38834
rect 12026 38820 12064 38834
rect 12098 38820 12136 38834
rect 12170 38820 12208 38834
rect 12242 38820 12280 38834
rect 12314 38820 12352 38834
rect 12386 38820 12424 38834
rect 12458 38820 12496 38834
rect 12530 38820 12568 38834
rect 12602 38820 12640 38834
rect 12674 38820 12712 38834
rect 12746 38820 12784 38834
rect 12818 38820 12856 38834
rect 12890 38820 12928 38834
rect 12962 38820 13000 38834
rect 13034 38820 13072 38834
rect 13106 38820 13118 38834
rect 2475 38814 13118 38820
rect 2475 37380 2532 38814
tri 2532 38783 2563 38814 nw
tri 13487 38726 13515 38754 se
rect 13515 38726 13521 38987
rect 2673 38720 2791 38726
rect 2725 38668 2739 38720
rect 2673 38656 2791 38668
rect 2725 38604 2739 38656
rect 2673 38592 2791 38604
rect 2725 38540 2739 38592
rect 2673 38534 2679 38540
rect 2713 38534 2751 38540
rect 2785 38534 2791 38540
rect 2673 38528 2791 38534
rect 2725 38476 2739 38528
rect 2673 38464 2679 38476
rect 2713 38464 2751 38476
rect 2785 38464 2791 38476
rect 2725 38422 2739 38464
rect 2673 38400 2679 38412
rect 2785 38400 2791 38412
rect 2673 38336 2679 38348
rect 2785 38336 2791 38348
rect 2673 38271 2679 38284
rect 2785 38271 2791 38284
rect 2673 38206 2679 38219
rect 2785 38206 2791 38219
rect 2673 38141 2679 38154
rect 2785 38141 2791 38154
rect 2673 38076 2679 38089
rect 2785 38076 2791 38089
rect 2673 38011 2679 38024
rect 2785 38011 2791 38024
rect 2673 37946 2679 37959
rect 2785 37946 2791 37959
rect 2673 37881 2679 37894
rect 2785 37881 2791 37894
rect 2673 37816 2679 37829
rect 2785 37816 2791 37829
rect 2673 37751 2679 37764
rect 2785 37751 2791 37764
rect 2673 37686 2679 37699
rect 2785 37686 2791 37699
rect 2673 37621 2679 37634
rect 2785 37621 2791 37634
rect 2673 37556 2679 37569
rect 2785 37556 2791 37569
rect 2673 37491 2679 37504
rect 2785 37491 2791 37504
rect 2673 37426 2679 37439
rect 2785 37426 2791 37439
tri 2532 37380 2537 37385 sw
rect 2475 37368 2537 37380
tri 2537 37368 2549 37380 sw
rect 2725 37374 2739 37380
rect 2673 37368 2791 37374
rect 2950 38714 3068 38726
rect 2950 38680 2956 38714
rect 2990 38680 3028 38714
rect 3062 38680 3068 38714
rect 2950 38641 3068 38680
rect 2950 38607 2956 38641
rect 2990 38607 3028 38641
rect 3062 38607 3068 38641
rect 2950 38568 3068 38607
rect 2950 38534 2956 38568
rect 2990 38534 3028 38568
rect 3062 38534 3068 38568
rect 2950 38495 3068 38534
rect 2950 38461 2956 38495
rect 2990 38461 3028 38495
rect 3062 38461 3068 38495
rect 2950 38422 3068 38461
rect 2950 37892 2956 38422
rect 3062 37892 3068 38422
rect 2950 37825 2956 37840
rect 3062 37825 3068 37840
rect 2950 37758 2956 37773
rect 3062 37758 3068 37773
rect 2950 37691 2956 37706
rect 3062 37691 3068 37706
rect 2950 37624 2956 37639
rect 3062 37624 3068 37639
rect 2950 37557 2956 37572
rect 3062 37557 3068 37572
rect 2950 37490 2956 37505
rect 3062 37490 3068 37505
rect 2950 37423 2956 37438
rect 3062 37423 3068 37438
rect 3002 37371 3016 37380
rect 2475 37336 2549 37368
tri 2549 37336 2581 37368 sw
rect 2950 37356 3068 37371
rect 2475 37324 2867 37336
rect 2475 37290 2482 37324
rect 2516 37290 2568 37324
rect 2602 37290 2654 37324
rect 2688 37290 2740 37324
rect 2774 37290 2826 37324
rect 2860 37290 2867 37324
rect 2475 37247 2867 37290
rect 2475 37213 2482 37247
rect 2516 37213 2568 37247
rect 2602 37213 2654 37247
rect 2688 37213 2740 37247
rect 2774 37213 2826 37247
rect 2860 37213 2867 37247
rect 2475 37170 2867 37213
rect 2475 37136 2482 37170
rect 2516 37136 2568 37170
rect 2602 37136 2654 37170
rect 2688 37136 2740 37170
rect 2774 37136 2826 37170
rect 2860 37136 2867 37170
rect 2475 37093 2867 37136
rect 2475 37059 2482 37093
rect 2516 37059 2568 37093
rect 2602 37059 2654 37093
rect 2688 37059 2740 37093
rect 2774 37059 2826 37093
rect 2860 37059 2867 37093
rect 2475 37016 2867 37059
rect 3002 37304 3016 37356
rect 2950 37289 3068 37304
rect 3002 37237 3016 37289
rect 2950 37222 3068 37237
rect 3002 37170 3016 37222
rect 2950 37155 3068 37170
rect 3002 37103 3016 37155
rect 2950 37088 3068 37103
rect 3002 37036 3016 37088
rect 2950 37030 3068 37036
rect 3227 38720 3345 38726
rect 3279 38668 3293 38720
rect 3227 38654 3345 38668
rect 3279 38602 3293 38654
rect 3227 38588 3345 38602
rect 3279 38536 3293 38588
rect 3227 38534 3233 38536
rect 3267 38534 3305 38536
rect 3339 38534 3345 38536
rect 3227 38522 3345 38534
rect 3279 38470 3293 38522
rect 3227 38461 3233 38470
rect 3267 38461 3305 38470
rect 3339 38461 3345 38470
rect 3227 38456 3345 38461
rect 3279 38422 3293 38456
rect 3227 38390 3233 38404
rect 3339 38390 3345 38404
rect 3227 38323 3233 38338
rect 3339 38323 3345 38338
rect 3227 38256 3233 38271
rect 3339 38256 3345 38271
rect 3227 37380 3233 38204
rect 3339 37380 3345 38204
rect 2475 36982 2482 37016
rect 2516 36982 2568 37016
rect 2602 36982 2654 37016
rect 2688 36982 2740 37016
rect 2774 36982 2826 37016
rect 2860 36982 2867 37016
rect 2475 36939 2867 36982
rect 2475 36905 2482 36939
rect 2516 36905 2568 36939
rect 2602 36905 2654 36939
rect 2688 36905 2740 36939
rect 2774 36905 2826 36939
rect 2860 36905 2867 36939
rect 2475 36862 2867 36905
rect 2475 36828 2482 36862
rect 2516 36828 2568 36862
rect 2602 36828 2654 36862
rect 2688 36828 2740 36862
rect 2774 36828 2826 36862
rect 2860 36828 2867 36862
rect 2475 36816 2867 36828
tri 2475 36714 2577 36816 ne
rect 2577 36714 2867 36816
rect 2213 36656 2219 36690
rect 2253 36672 2291 36684
rect 2325 36672 2363 36684
rect 2397 36657 2403 36691
tri 2577 36680 2611 36714 ne
rect 2611 36680 2867 36714
rect 2213 36620 2249 36656
rect 2301 36620 2315 36656
rect 2367 36620 2403 36657
tri 2611 36641 2650 36680 ne
rect 2650 36641 2867 36680
tri 2650 36624 2667 36641 ne
rect 2213 36618 2403 36620
rect 2213 36617 2363 36618
rect 2213 36583 2219 36617
rect 2253 36608 2291 36617
rect 2325 36608 2363 36617
rect 2397 36584 2403 36618
rect 2213 36556 2249 36583
rect 2301 36556 2315 36583
rect 2367 36556 2403 36584
rect 2213 36545 2403 36556
rect 2213 36544 2363 36545
rect 2213 36510 2219 36544
rect 2397 36511 2403 36545
rect 2213 36492 2249 36510
rect 2301 36492 2315 36510
rect 2367 36492 2403 36511
rect 2213 36480 2403 36492
rect 2213 36471 2249 36480
rect 2301 36471 2315 36480
rect 2367 36472 2403 36480
rect 2213 36437 2219 36471
rect 2397 36438 2403 36472
rect 2213 36428 2249 36437
rect 2301 36428 2315 36437
rect 2367 36428 2403 36438
rect 2213 36416 2403 36428
rect 2213 36398 2249 36416
rect 2301 36398 2315 36416
rect 2367 36399 2403 36416
rect 2213 36364 2219 36398
rect 2397 36365 2403 36399
rect 2367 36364 2403 36365
rect 2213 36352 2403 36364
rect 2213 36325 2249 36352
rect 2301 36325 2315 36352
rect 2367 36326 2403 36352
rect 2213 36291 2219 36325
rect 2253 36291 2291 36300
rect 2325 36292 2363 36300
rect 2397 36292 2403 36326
rect 2325 36291 2403 36292
rect 2213 36288 2403 36291
rect 2213 36252 2249 36288
rect 2301 36252 2315 36288
rect 2367 36253 2403 36288
rect 2213 36218 2219 36252
rect 2253 36224 2291 36236
rect 2325 36224 2363 36236
rect 2397 36219 2403 36253
rect 2213 36179 2249 36218
rect 2301 36179 2315 36218
rect 2367 36180 2403 36219
rect 2213 36145 2219 36179
rect 2253 36160 2291 36172
rect 2325 36160 2363 36172
rect 2397 36146 2403 36180
rect 2213 36108 2249 36145
rect 2301 36108 2315 36145
rect 2367 36108 2403 36146
rect 2213 36107 2403 36108
rect 2213 36106 2363 36107
rect 2213 36072 2219 36106
rect 2253 36096 2291 36106
rect 2325 36096 2363 36106
rect 2397 36073 2403 36107
rect 2213 36044 2249 36072
rect 2301 36044 2315 36072
rect 2367 36044 2403 36073
rect 2213 36034 2403 36044
rect 2213 36033 2363 36034
rect 2213 35999 2219 36033
rect 2253 36032 2291 36033
rect 2325 36032 2363 36033
rect 2397 36000 2403 36034
rect 2213 35980 2249 35999
rect 2301 35980 2315 35999
rect 2367 35980 2403 36000
rect 2213 35968 2403 35980
rect 2213 35960 2249 35968
rect 2301 35960 2315 35968
rect 2367 35961 2403 35968
rect 2213 35926 2219 35960
rect 2397 35927 2403 35961
rect 2213 35916 2249 35926
rect 2301 35916 2315 35926
rect 2367 35916 2403 35927
rect 2213 35904 2403 35916
rect 2213 35887 2249 35904
rect 2301 35887 2315 35904
rect 2367 35888 2403 35904
rect 2213 35853 2219 35887
rect 2397 35854 2403 35888
rect 2213 35852 2249 35853
rect 2301 35852 2315 35853
rect 2367 35852 2403 35854
rect 2213 35840 2403 35852
rect 2213 35814 2249 35840
rect 2301 35814 2315 35840
rect 2367 35815 2403 35840
rect 2213 35780 2219 35814
rect 2253 35780 2291 35788
rect 2325 35781 2363 35788
rect 2397 35781 2403 35815
rect 2325 35780 2403 35781
rect 2213 35776 2403 35780
rect 2213 35741 2249 35776
rect 2301 35741 2315 35776
rect 2367 35742 2403 35776
rect 2213 35707 2219 35741
rect 2253 35712 2291 35724
rect 2325 35712 2363 35724
rect 2397 35708 2403 35742
rect 2213 35668 2249 35707
rect 2301 35668 2315 35707
rect 2367 35669 2403 35708
rect 2213 35634 2219 35668
rect 2253 35648 2291 35660
rect 2325 35648 2363 35660
rect 2397 35635 2403 35669
rect 2213 35596 2249 35634
rect 2301 35596 2315 35634
rect 2367 35596 2403 35635
rect 2213 35595 2363 35596
rect 2213 35561 2219 35595
rect 2253 35584 2291 35595
rect 2325 35584 2363 35595
rect 2397 35562 2403 35596
rect 2213 35532 2249 35561
rect 2301 35532 2315 35561
rect 2367 35532 2403 35562
rect 2213 35523 2403 35532
rect 2213 35522 2363 35523
rect 2213 33688 2219 35522
rect 2325 35520 2363 35522
rect 2397 35489 2403 35523
rect 2367 35468 2403 35489
rect 2325 35456 2403 35468
rect 2367 35450 2403 35456
rect 2397 33688 2403 35450
rect 2213 33676 2249 33688
rect 2301 33676 2315 33688
rect 2367 33676 2403 33688
rect 2213 33664 2403 33676
rect 2213 33644 2249 33664
rect 2213 33610 2219 33644
rect 2301 33612 2315 33664
rect 2367 33656 2403 33664
tri 2367 33620 2403 33656 nw
rect 2667 35321 2867 36641
rect 3227 36720 3345 37380
rect 3279 36668 3293 36720
rect 3227 36654 3345 36668
rect 3279 36602 3293 36654
rect 3227 36588 3345 36602
rect 3279 36536 3293 36588
rect 3227 36534 3233 36536
rect 3267 36534 3305 36536
rect 3339 36534 3345 36536
rect 3227 36522 3345 36534
rect 3279 36470 3293 36522
rect 3227 36461 3233 36470
rect 3267 36461 3305 36470
rect 3339 36461 3345 36470
rect 3227 36456 3345 36461
rect 3279 36422 3293 36456
rect 3227 36390 3233 36404
rect 3339 36390 3345 36404
rect 3227 36323 3233 36338
rect 3339 36323 3345 36338
rect 3227 36256 3233 36271
rect 3339 36256 3345 36271
rect 3227 35380 3233 36204
rect 3339 35380 3345 36204
rect 3227 35368 3345 35380
rect 3504 38714 3622 38726
rect 3504 38680 3510 38714
rect 3544 38680 3582 38714
rect 3616 38680 3622 38714
rect 3504 38641 3622 38680
rect 3504 38607 3510 38641
rect 3544 38607 3582 38641
rect 3616 38607 3622 38641
rect 3504 38568 3622 38607
rect 3504 38534 3510 38568
rect 3544 38534 3582 38568
rect 3616 38534 3622 38568
rect 3504 38495 3622 38534
rect 3504 38461 3510 38495
rect 3544 38461 3582 38495
rect 3616 38461 3622 38495
rect 3504 38422 3622 38461
rect 3504 37892 3510 38422
rect 3616 37892 3622 38422
rect 3504 37825 3510 37840
rect 3616 37825 3622 37840
rect 3504 37758 3510 37773
rect 3616 37758 3622 37773
rect 3504 37691 3510 37706
rect 3616 37691 3622 37706
rect 3504 37624 3510 37639
rect 3616 37624 3622 37639
rect 3504 37557 3510 37572
rect 3616 37557 3622 37572
rect 3504 37490 3510 37505
rect 3616 37490 3622 37505
rect 3504 37423 3510 37438
rect 3616 37423 3622 37438
rect 3556 37371 3570 37380
rect 3504 37356 3622 37371
rect 3556 37304 3570 37356
rect 3504 37289 3622 37304
rect 3556 37237 3570 37289
rect 3504 37222 3622 37237
rect 3556 37170 3570 37222
rect 3504 37155 3622 37170
rect 3556 37103 3570 37155
rect 3504 37088 3622 37103
rect 3556 37036 3570 37088
rect 3504 36714 3622 37036
rect 3504 36680 3510 36714
rect 3544 36680 3582 36714
rect 3616 36680 3622 36714
rect 3504 36641 3622 36680
rect 3504 36607 3510 36641
rect 3544 36607 3582 36641
rect 3616 36607 3622 36641
rect 3504 36568 3622 36607
rect 3504 36534 3510 36568
rect 3544 36534 3582 36568
rect 3616 36534 3622 36568
rect 3504 36495 3622 36534
rect 3504 36461 3510 36495
rect 3544 36461 3582 36495
rect 3616 36461 3622 36495
rect 3504 36422 3622 36461
rect 3504 35892 3510 36422
rect 3616 35892 3622 36422
rect 3504 35826 3510 35840
rect 3616 35826 3622 35840
rect 3504 35760 3510 35774
rect 3616 35760 3622 35774
rect 3504 35694 3510 35708
rect 3616 35694 3622 35708
rect 3504 35627 3510 35642
rect 3616 35627 3622 35642
rect 3504 35560 3510 35575
rect 3616 35560 3622 35575
rect 3504 35493 3510 35508
rect 3616 35493 3622 35508
rect 3504 35426 3510 35441
rect 3616 35426 3622 35441
rect 3556 35374 3570 35380
rect 2667 35287 2674 35321
rect 2708 35287 2750 35321
rect 2784 35287 2826 35321
rect 2860 35287 2867 35321
rect 2667 35244 2867 35287
rect 2667 35210 2674 35244
rect 2708 35210 2750 35244
rect 2784 35210 2826 35244
rect 2860 35210 2867 35244
rect 2667 35167 2867 35210
rect 2667 35133 2674 35167
rect 2708 35133 2750 35167
rect 2784 35133 2826 35167
rect 2860 35133 2867 35167
rect 2667 35089 2867 35133
rect 2667 35055 2674 35089
rect 2708 35055 2750 35089
rect 2784 35055 2826 35089
rect 2860 35055 2867 35089
rect 2667 35011 2867 35055
rect 2667 34977 2674 35011
rect 2708 34977 2750 35011
rect 2784 34977 2826 35011
rect 2860 34977 2867 35011
rect 2667 34933 2867 34977
rect 2667 34899 2674 34933
rect 2708 34899 2750 34933
rect 2784 34899 2826 34933
rect 2860 34899 2867 34933
rect 2667 34855 2867 34899
rect 2667 34821 2674 34855
rect 2708 34821 2750 34855
rect 2784 34821 2826 34855
rect 2860 34821 2867 34855
rect 2253 33610 2325 33612
rect 2359 33610 2367 33612
rect 2213 33600 2367 33610
rect 2213 33571 2249 33600
rect 2213 33537 2219 33571
rect 2301 33548 2315 33600
rect 2253 33537 2325 33548
rect 2359 33537 2367 33548
rect 2213 33536 2367 33537
rect 2213 33498 2249 33536
tri 1841 33464 1875 33498 se
rect 1875 33464 2007 33498
tri 2007 33464 2041 33498 nw
rect 2213 33464 2219 33498
rect 2301 33484 2315 33536
rect 2253 33472 2325 33484
rect 2359 33472 2367 33484
tri 1831 33454 1841 33464 se
rect 1841 33454 1997 33464
tri 1997 33454 2007 33464 nw
rect 1831 33425 1968 33454
tri 1968 33425 1997 33454 nw
rect 2213 33425 2249 33464
rect 1831 33228 1949 33425
tri 1949 33406 1968 33425 nw
rect 2213 33391 2219 33425
rect 2301 33420 2315 33472
rect 2253 33408 2325 33420
rect 2359 33408 2367 33420
rect 2213 33356 2249 33391
rect 2301 33356 2315 33408
rect 2213 33352 2367 33356
rect 2213 33318 2219 33352
rect 2253 33344 2325 33352
rect 2359 33344 2367 33352
rect 2213 33292 2249 33318
rect 2301 33292 2315 33344
rect 2213 33280 2367 33292
rect 2213 33279 2249 33280
rect 2213 33245 2219 33279
rect 2213 33228 2249 33245
rect 2301 33228 2315 33280
rect 2213 33216 2367 33228
rect 2213 33206 2249 33216
rect 2213 33172 2219 33206
rect 2213 33164 2249 33172
rect 2301 33164 2315 33216
rect 2213 33152 2367 33164
rect 2213 33133 2249 33152
rect 2213 33099 2219 33133
rect 2301 33100 2315 33152
rect 2253 33099 2325 33100
rect 2359 33099 2367 33100
rect 2213 33088 2367 33099
rect 2213 33060 2249 33088
rect 2213 33026 2219 33060
rect 2301 33036 2315 33088
rect 2253 33026 2325 33036
rect 2359 33026 2367 33036
rect 2213 33024 2367 33026
rect 2213 32987 2249 33024
rect 2213 32953 2219 32987
rect 2301 32972 2315 33024
rect 2253 32960 2325 32972
rect 2359 32960 2367 32972
rect 2213 32914 2249 32953
rect 2213 32880 2219 32914
rect 2301 32908 2315 32960
rect 2253 32896 2325 32908
rect 2359 32896 2367 32908
rect 2213 32844 2249 32880
rect 2301 32844 2315 32896
rect 2213 32841 2367 32844
rect 2213 32807 2219 32841
rect 2253 32832 2325 32841
rect 2359 32832 2367 32841
rect 2213 32780 2249 32807
rect 2301 32780 2315 32832
rect 2213 32768 2367 32780
rect 2213 32734 2219 32768
rect 2213 32716 2249 32734
rect 2301 32716 2315 32768
rect 2213 32704 2367 32716
rect 2213 32695 2249 32704
rect 2213 32661 2219 32695
rect 2213 32652 2249 32661
rect 2301 32652 2315 32704
rect 2213 32640 2367 32652
rect 2213 32622 2249 32640
rect 2213 32588 2219 32622
rect 2301 32588 2315 32640
rect 2213 32576 2367 32588
rect 2213 32549 2249 32576
rect 2213 32515 2219 32549
rect 2301 32524 2315 32576
rect 2253 32515 2325 32524
rect 2359 32515 2367 32524
rect 2213 32512 2367 32515
rect 2213 32476 2249 32512
rect 2213 32442 2219 32476
rect 2301 32460 2315 32512
rect 2253 32448 2325 32460
rect 2359 32448 2367 32460
rect 2213 32403 2249 32442
rect 2213 32369 2219 32403
rect 2301 32396 2315 32448
rect 2253 32384 2325 32396
rect 2359 32384 2367 32396
rect 2213 32332 2249 32369
rect 2301 32332 2315 32384
rect 2213 32330 2367 32332
rect 2213 32296 2219 32330
rect 2253 32319 2325 32330
rect 2359 32319 2367 32330
rect 2213 32267 2249 32296
rect 2301 32267 2315 32319
rect 2213 32257 2367 32267
rect 2213 32223 2219 32257
rect 2253 32254 2325 32257
rect 2359 32254 2367 32257
rect 2213 32202 2249 32223
rect 2301 32202 2315 32254
rect 2213 32189 2367 32202
rect 2213 32184 2249 32189
rect 2213 32150 2219 32184
rect 2213 32137 2249 32150
rect 2301 32137 2315 32189
rect 2213 32124 2367 32137
rect 2213 32111 2249 32124
rect 2213 32077 2219 32111
rect 2213 32072 2249 32077
rect 2301 32072 2315 32124
rect 2213 32059 2367 32072
rect 2213 32038 2249 32059
rect 2213 32004 2219 32038
rect 2301 32007 2315 32059
rect 2253 32004 2325 32007
rect 2359 32004 2367 32007
rect 2213 31994 2367 32004
rect 2213 31965 2249 31994
rect 2213 31931 2219 31965
rect 2301 31942 2315 31994
rect 2253 31931 2325 31942
rect 2359 31931 2367 31942
rect 2213 31929 2367 31931
rect 2213 31892 2249 31929
rect 2213 31858 2219 31892
rect 2301 31877 2315 31929
rect 2253 31864 2325 31877
rect 2359 31864 2367 31877
rect 2213 31819 2249 31858
rect 2213 31785 2219 31819
rect 2301 31812 2315 31864
rect 2253 31799 2325 31812
rect 2359 31799 2367 31812
rect 2213 31747 2249 31785
rect 2301 31747 2315 31799
rect 2213 31746 2367 31747
rect 2213 31712 2219 31746
rect 2253 31734 2325 31746
rect 2359 31734 2367 31746
rect 2213 31682 2249 31712
rect 2301 31682 2315 31734
rect 2213 31673 2367 31682
rect 2213 31639 2219 31673
rect 2253 31669 2325 31673
rect 2359 31669 2367 31673
rect 2213 31617 2249 31639
rect 2301 31617 2315 31669
rect 2213 31604 2367 31617
rect 2213 31600 2249 31604
rect 2213 31566 2219 31600
rect 2213 31552 2249 31566
rect 2301 31552 2315 31604
rect 2213 31539 2367 31552
rect 2213 31527 2249 31539
rect 2213 31493 2219 31527
rect 2213 31487 2249 31493
rect 2301 31487 2315 31539
rect 2213 31474 2367 31487
rect 2213 31454 2249 31474
rect 2213 31420 2219 31454
rect 2301 31422 2315 31474
rect 2253 31420 2325 31422
rect 2359 31420 2367 31422
rect 2213 31409 2367 31420
rect 2213 31381 2249 31409
rect 2213 31347 2219 31381
rect 2301 31357 2315 31409
rect 2253 31347 2325 31357
rect 2359 31347 2367 31357
rect 2213 31344 2367 31347
rect 2213 31308 2249 31344
rect 2213 31274 2219 31308
rect 2301 31292 2315 31344
rect 2253 31279 2325 31292
rect 2359 31279 2367 31292
rect 2213 31235 2249 31274
rect 2213 31201 2219 31235
rect 2301 31227 2315 31279
rect 2253 31214 2325 31227
rect 2359 31214 2367 31227
rect 2213 31162 2249 31201
rect 2301 31162 2315 31214
rect 2213 31128 2219 31162
rect 2253 31149 2325 31162
rect 2359 31149 2367 31162
rect 2213 31097 2249 31128
rect 2301 31097 2315 31149
rect 2213 31089 2367 31097
rect 2213 31055 2219 31089
rect 2253 31084 2325 31089
rect 2359 31084 2367 31089
rect 2213 31032 2249 31055
rect 2301 31032 2315 31084
rect 2213 31019 2367 31032
rect 2213 31016 2249 31019
rect 2213 30982 2219 31016
rect 2213 30967 2249 30982
rect 2301 30967 2315 31019
rect 2213 30954 2367 30967
rect 2213 30943 2249 30954
rect 2213 30909 2219 30943
rect 2213 30902 2249 30909
rect 2301 30902 2315 30954
rect 2213 30889 2367 30902
rect 2213 30871 2249 30889
rect 2213 30837 2219 30871
rect 2301 30837 2315 30889
rect 2213 30824 2367 30837
rect 2213 30799 2249 30824
rect 2213 30765 2219 30799
rect 2301 30772 2315 30824
rect 2253 30765 2325 30772
rect 2359 30765 2367 30772
rect 2213 30759 2367 30765
rect 2213 30727 2249 30759
rect 2213 30693 2219 30727
rect 2301 30707 2315 30759
rect 2253 30694 2325 30707
rect 2359 30694 2367 30707
rect 2213 30655 2249 30693
rect 2213 30621 2219 30655
rect 2301 30642 2315 30694
rect 2253 30629 2325 30642
rect 2359 30629 2367 30642
rect 2213 30583 2249 30621
rect 2213 30549 2219 30583
rect 2301 30577 2315 30629
rect 2253 30564 2325 30577
rect 2359 30564 2367 30577
rect 2213 30512 2249 30549
rect 2301 30512 2315 30564
rect 2213 30511 2367 30512
rect 2213 30477 2219 30511
rect 2253 30499 2325 30511
rect 2359 30499 2367 30511
rect 2213 30447 2249 30477
rect 2301 30447 2315 30499
rect 2213 30439 2367 30447
rect 2213 30405 2219 30439
rect 2253 30434 2325 30439
rect 2359 30434 2367 30439
rect 2213 30382 2249 30405
rect 2301 30382 2315 30434
rect 2213 30369 2367 30382
rect 2213 30367 2249 30369
rect 2213 30333 2219 30367
rect 2213 30317 2249 30333
rect 2301 30317 2315 30369
rect 2213 30304 2367 30317
rect 2213 30295 2249 30304
rect 2213 30261 2219 30295
rect 2213 30252 2249 30261
rect 2301 30252 2315 30304
rect 2213 30239 2367 30252
rect 2213 30223 2249 30239
rect 2213 30189 2219 30223
rect 2213 30187 2249 30189
rect 2301 30187 2315 30239
rect 2213 30174 2367 30187
rect 2213 30151 2249 30174
rect 2213 30117 2219 30151
rect 2301 30122 2315 30174
rect 2253 30117 2325 30122
rect 2359 30117 2367 30122
rect 2213 30109 2367 30117
rect 2213 30079 2249 30109
rect 2213 30045 2219 30079
rect 2301 30057 2315 30109
rect 2253 30045 2325 30057
rect 2359 30045 2367 30057
rect 2213 30044 2367 30045
rect 2213 30007 2249 30044
rect 2213 29973 2219 30007
rect 2301 29992 2315 30044
rect 2253 29979 2325 29992
rect 2359 29979 2367 29992
rect 2213 29935 2249 29973
rect 2213 29901 2219 29935
rect 2301 29927 2315 29979
rect 2253 29914 2325 29927
rect 2359 29914 2367 29927
rect 2213 29863 2249 29901
rect 2213 29829 2219 29863
rect 2301 29862 2315 29914
rect 2253 29849 2325 29862
rect 2359 29849 2367 29862
rect 2213 29797 2249 29829
rect 2301 29797 2315 29849
rect 2213 29791 2367 29797
rect 2213 29757 2219 29791
rect 2253 29784 2325 29791
rect 2359 29784 2367 29791
rect 2213 29732 2249 29757
rect 2301 29732 2315 29784
rect 2213 29719 2367 29732
rect 2213 29685 2219 29719
rect 2213 29667 2249 29685
rect 2301 29667 2315 29719
rect 2213 29654 2367 29667
rect 2213 29647 2249 29654
rect 2213 29613 2219 29647
rect 2213 29602 2249 29613
rect 2301 29602 2315 29654
rect 2213 29589 2367 29602
rect 2213 29575 2249 29589
rect 2213 29541 2219 29575
rect 2213 29537 2249 29541
rect 2301 29537 2315 29589
rect 2213 29524 2367 29537
rect 2213 29503 2249 29524
rect 2213 29469 2219 29503
rect 2301 29472 2315 29524
rect 2253 29469 2325 29472
rect 2359 29469 2367 29472
rect 2213 29459 2367 29469
rect 2213 29431 2249 29459
rect 2213 29397 2219 29431
rect 2301 29407 2315 29459
rect 2253 29397 2325 29407
rect 2359 29397 2367 29407
rect 2213 29394 2367 29397
rect 2213 29359 2249 29394
rect 2213 29325 2219 29359
rect 2301 29342 2315 29394
rect 2253 29329 2325 29342
rect 2359 29329 2367 29342
rect 2213 29287 2249 29325
rect 2213 29253 2219 29287
rect 2301 29277 2315 29329
rect 2253 29264 2325 29277
rect 2359 29264 2367 29277
rect 2213 29215 2249 29253
rect 2213 29181 2219 29215
rect 2301 29212 2315 29264
rect 2253 29199 2325 29212
rect 2359 29199 2367 29212
rect 2213 29147 2249 29181
rect 2301 29147 2315 29199
rect 2213 29143 2367 29147
rect 2213 29109 2219 29143
rect 2253 29134 2325 29143
rect 2359 29134 2367 29143
rect 2213 29082 2249 29109
rect 2301 29082 2315 29134
rect 2213 29071 2367 29082
rect 2213 29037 2219 29071
rect 2253 29069 2325 29071
rect 2359 29069 2367 29071
rect 2213 29017 2249 29037
rect 2301 29017 2315 29069
rect 2213 29004 2367 29017
rect 2213 28999 2249 29004
rect 2213 28965 2219 28999
rect 2213 28952 2249 28965
rect 2301 28952 2315 29004
rect 2213 28939 2367 28952
rect 2213 28927 2249 28939
rect 2213 28893 2219 28927
rect 2213 28887 2249 28893
rect 2301 28887 2315 28939
rect 2213 28881 2367 28887
rect 2667 33322 2867 34821
rect 3504 35280 3622 35374
rect 3781 38720 3899 38726
rect 3833 38668 3847 38720
rect 3781 38654 3899 38668
rect 3833 38602 3847 38654
rect 3781 38588 3899 38602
rect 3833 38536 3847 38588
rect 3781 38534 3787 38536
rect 3821 38534 3859 38536
rect 3893 38534 3899 38536
rect 3781 38522 3899 38534
rect 3833 38470 3847 38522
rect 3781 38461 3787 38470
rect 3821 38461 3859 38470
rect 3893 38461 3899 38470
rect 3781 38456 3899 38461
rect 3833 38422 3847 38456
rect 3781 38390 3787 38404
rect 3893 38390 3899 38404
rect 3781 38323 3787 38338
rect 3893 38323 3899 38338
rect 3781 38256 3787 38271
rect 3893 38256 3899 38271
rect 3781 37380 3787 38204
rect 3893 37380 3899 38204
rect 3781 36720 3899 37380
rect 3833 36668 3847 36720
rect 3781 36654 3899 36668
rect 3833 36602 3847 36654
rect 3781 36588 3899 36602
rect 3833 36536 3847 36588
rect 3781 36534 3787 36536
rect 3821 36534 3859 36536
rect 3893 36534 3899 36536
rect 3781 36522 3899 36534
rect 3833 36470 3847 36522
rect 3781 36461 3787 36470
rect 3821 36461 3859 36470
rect 3893 36461 3899 36470
rect 3781 36456 3899 36461
rect 3833 36422 3847 36456
rect 3781 36390 3787 36404
rect 3893 36390 3899 36404
rect 3781 36323 3787 36338
rect 3893 36323 3899 36338
rect 3781 36256 3787 36271
rect 3893 36256 3899 36271
rect 3781 35380 3787 36204
rect 3893 35380 3899 36204
rect 3781 35368 3899 35380
rect 4058 38714 4176 38726
rect 4058 38680 4064 38714
rect 4098 38680 4136 38714
rect 4170 38680 4176 38714
rect 4058 38641 4176 38680
rect 4058 38607 4064 38641
rect 4098 38607 4136 38641
rect 4170 38607 4176 38641
rect 4058 38568 4176 38607
rect 4058 38534 4064 38568
rect 4098 38534 4136 38568
rect 4170 38534 4176 38568
rect 4058 38495 4176 38534
rect 4058 38461 4064 38495
rect 4098 38461 4136 38495
rect 4170 38461 4176 38495
rect 4058 38422 4176 38461
rect 4058 37892 4064 38422
rect 4170 37892 4176 38422
rect 4058 37825 4064 37840
rect 4170 37825 4176 37840
rect 4058 37758 4064 37773
rect 4170 37758 4176 37773
rect 4058 37691 4064 37706
rect 4170 37691 4176 37706
rect 4058 37624 4064 37639
rect 4170 37624 4176 37639
rect 4058 37557 4064 37572
rect 4170 37557 4176 37572
rect 4058 37490 4064 37505
rect 4170 37490 4176 37505
rect 4058 37423 4064 37438
rect 4170 37423 4176 37438
rect 4110 37371 4124 37380
rect 4058 37356 4176 37371
rect 4110 37304 4124 37356
rect 4058 37289 4176 37304
rect 4110 37237 4124 37289
rect 4058 37222 4176 37237
rect 4110 37170 4124 37222
rect 4058 37155 4176 37170
rect 4110 37103 4124 37155
rect 4058 37088 4176 37103
rect 4110 37036 4124 37088
rect 4058 36714 4176 37036
rect 4058 36680 4064 36714
rect 4098 36680 4136 36714
rect 4170 36680 4176 36714
rect 4058 36641 4176 36680
rect 4058 36607 4064 36641
rect 4098 36607 4136 36641
rect 4170 36607 4176 36641
rect 4058 36568 4176 36607
rect 4058 36534 4064 36568
rect 4098 36534 4136 36568
rect 4170 36534 4176 36568
rect 4058 36495 4176 36534
rect 4058 36461 4064 36495
rect 4098 36461 4136 36495
rect 4170 36461 4176 36495
rect 4058 36422 4176 36461
rect 4058 35892 4064 36422
rect 4170 35892 4176 36422
rect 4058 35826 4064 35840
rect 4170 35826 4176 35840
rect 4058 35760 4064 35774
rect 4170 35760 4176 35774
rect 4058 35694 4064 35708
rect 4170 35694 4176 35708
rect 4058 35627 4064 35642
rect 4170 35627 4176 35642
rect 4058 35560 4064 35575
rect 4170 35560 4176 35575
rect 4058 35493 4064 35508
rect 4170 35493 4176 35508
rect 4058 35426 4064 35441
rect 4170 35426 4176 35441
rect 4110 35374 4124 35380
tri 3622 35280 3666 35324 sw
tri 4014 35280 4058 35324 se
rect 4058 35280 4176 35374
rect 4335 38720 4453 38726
rect 4387 38668 4401 38720
rect 4335 38654 4453 38668
rect 4387 38602 4401 38654
rect 4335 38588 4453 38602
rect 4387 38536 4401 38588
rect 4335 38534 4341 38536
rect 4375 38534 4413 38536
rect 4447 38534 4453 38536
rect 4335 38522 4453 38534
rect 4387 38470 4401 38522
rect 4335 38461 4341 38470
rect 4375 38461 4413 38470
rect 4447 38461 4453 38470
rect 4335 38456 4453 38461
rect 4387 38422 4401 38456
rect 4335 38390 4341 38404
rect 4447 38390 4453 38404
rect 4335 38323 4341 38338
rect 4447 38323 4453 38338
rect 4335 38256 4341 38271
rect 4447 38256 4453 38271
rect 4335 37380 4341 38204
rect 4447 37380 4453 38204
rect 4335 36720 4453 37380
rect 4387 36668 4401 36720
rect 4335 36654 4453 36668
rect 4387 36602 4401 36654
rect 4335 36588 4453 36602
rect 4387 36536 4401 36588
rect 4335 36534 4341 36536
rect 4375 36534 4413 36536
rect 4447 36534 4453 36536
rect 4335 36522 4453 36534
rect 4387 36470 4401 36522
rect 4335 36461 4341 36470
rect 4375 36461 4413 36470
rect 4447 36461 4453 36470
rect 4335 36456 4453 36461
rect 4387 36422 4401 36456
rect 4335 36390 4341 36404
rect 4447 36390 4453 36404
rect 4335 36323 4341 36338
rect 4447 36323 4453 36338
rect 4335 36256 4341 36271
rect 4447 36256 4453 36271
rect 4335 35380 4341 36204
rect 4447 35380 4453 36204
rect 4335 35368 4453 35380
rect 4612 38714 4730 38726
rect 4612 38680 4618 38714
rect 4652 38680 4690 38714
rect 4724 38680 4730 38714
rect 4612 38641 4730 38680
rect 4612 38607 4618 38641
rect 4652 38607 4690 38641
rect 4724 38607 4730 38641
rect 4612 38568 4730 38607
rect 4612 38534 4618 38568
rect 4652 38534 4690 38568
rect 4724 38534 4730 38568
rect 4612 38495 4730 38534
rect 4612 38461 4618 38495
rect 4652 38461 4690 38495
rect 4724 38461 4730 38495
rect 4612 38422 4730 38461
rect 4612 37892 4618 38422
rect 4724 37892 4730 38422
rect 4612 37825 4618 37840
rect 4724 37825 4730 37840
rect 4612 37758 4618 37773
rect 4724 37758 4730 37773
rect 4612 37691 4618 37706
rect 4724 37691 4730 37706
rect 4612 37624 4618 37639
rect 4724 37624 4730 37639
rect 4612 37557 4618 37572
rect 4724 37557 4730 37572
rect 4612 37490 4618 37505
rect 4724 37490 4730 37505
rect 4612 37423 4618 37438
rect 4724 37423 4730 37438
rect 4664 37371 4678 37380
rect 4612 37356 4730 37371
rect 4664 37304 4678 37356
rect 4612 37289 4730 37304
rect 4664 37237 4678 37289
rect 4612 37222 4730 37237
rect 4664 37170 4678 37222
rect 4612 37155 4730 37170
rect 4664 37103 4678 37155
rect 4612 37088 4730 37103
rect 4664 37036 4678 37088
rect 4612 36714 4730 37036
rect 4612 36680 4618 36714
rect 4652 36680 4690 36714
rect 4724 36680 4730 36714
rect 4612 36641 4730 36680
rect 4612 36607 4618 36641
rect 4652 36607 4690 36641
rect 4724 36607 4730 36641
rect 4612 36568 4730 36607
rect 4612 36534 4618 36568
rect 4652 36534 4690 36568
rect 4724 36534 4730 36568
rect 4612 36495 4730 36534
rect 4612 36461 4618 36495
rect 4652 36461 4690 36495
rect 4724 36461 4730 36495
rect 4612 36422 4730 36461
rect 4612 35892 4618 36422
rect 4724 35892 4730 36422
rect 4612 35826 4618 35840
rect 4724 35826 4730 35840
rect 4612 35760 4618 35774
rect 4724 35760 4730 35774
rect 4612 35694 4618 35708
rect 4724 35694 4730 35708
rect 4612 35627 4618 35642
rect 4724 35627 4730 35642
rect 4612 35560 4618 35575
rect 4724 35560 4730 35575
rect 4612 35493 4618 35508
rect 4724 35493 4730 35508
rect 4612 35426 4618 35441
rect 4724 35426 4730 35441
rect 4664 35374 4678 35380
tri 4176 35280 4220 35324 sw
tri 4568 35280 4612 35324 se
rect 4612 35280 4730 35374
rect 4889 38720 5007 38726
rect 4941 38668 4955 38720
rect 4889 38654 5007 38668
rect 4941 38602 4955 38654
rect 4889 38588 5007 38602
rect 4941 38536 4955 38588
rect 4889 38534 4895 38536
rect 4929 38534 4967 38536
rect 5001 38534 5007 38536
rect 4889 38522 5007 38534
rect 4941 38470 4955 38522
rect 4889 38461 4895 38470
rect 4929 38461 4967 38470
rect 5001 38461 5007 38470
rect 4889 38456 5007 38461
rect 4941 38422 4955 38456
rect 4889 38390 4895 38404
rect 5001 38390 5007 38404
rect 4889 38323 4895 38338
rect 5001 38323 5007 38338
rect 4889 38256 4895 38271
rect 5001 38256 5007 38271
rect 4889 37380 4895 38204
rect 5001 37380 5007 38204
rect 4889 36720 5007 37380
rect 4941 36668 4955 36720
rect 4889 36654 5007 36668
rect 4941 36602 4955 36654
rect 4889 36588 5007 36602
rect 4941 36536 4955 36588
rect 4889 36534 4895 36536
rect 4929 36534 4967 36536
rect 5001 36534 5007 36536
rect 4889 36522 5007 36534
rect 4941 36470 4955 36522
rect 4889 36461 4895 36470
rect 4929 36461 4967 36470
rect 5001 36461 5007 36470
rect 4889 36456 5007 36461
rect 4941 36422 4955 36456
rect 4889 36390 4895 36404
rect 5001 36390 5007 36404
rect 4889 36323 4895 36338
rect 5001 36323 5007 36338
rect 4889 36256 4895 36271
rect 5001 36256 5007 36271
rect 4889 35380 4895 36204
rect 5001 35380 5007 36204
rect 4889 35368 5007 35380
rect 5166 38714 5284 38726
rect 5166 38680 5172 38714
rect 5206 38680 5244 38714
rect 5278 38680 5284 38714
rect 5166 38641 5284 38680
rect 5166 38607 5172 38641
rect 5206 38607 5244 38641
rect 5278 38607 5284 38641
rect 5166 38568 5284 38607
rect 5166 38534 5172 38568
rect 5206 38534 5244 38568
rect 5278 38534 5284 38568
rect 5166 38495 5284 38534
rect 5166 38461 5172 38495
rect 5206 38461 5244 38495
rect 5278 38461 5284 38495
rect 5166 38422 5284 38461
rect 5166 37892 5172 38422
rect 5278 37892 5284 38422
rect 5166 37825 5172 37840
rect 5278 37825 5284 37840
rect 5166 37758 5172 37773
rect 5278 37758 5284 37773
rect 5166 37691 5172 37706
rect 5278 37691 5284 37706
rect 5166 37624 5172 37639
rect 5278 37624 5284 37639
rect 5166 37557 5172 37572
rect 5278 37557 5284 37572
rect 5166 37490 5172 37505
rect 5278 37490 5284 37505
rect 5166 37423 5172 37438
rect 5278 37423 5284 37438
rect 5218 37371 5232 37380
rect 5166 37356 5284 37371
rect 5218 37304 5232 37356
rect 5166 37289 5284 37304
rect 5218 37237 5232 37289
rect 5166 37222 5284 37237
rect 5218 37170 5232 37222
rect 5166 37155 5284 37170
rect 5218 37103 5232 37155
rect 5166 37088 5284 37103
rect 5218 37036 5232 37088
rect 5166 36714 5284 37036
rect 5166 36680 5172 36714
rect 5206 36680 5244 36714
rect 5278 36680 5284 36714
rect 5166 36641 5284 36680
rect 5166 36607 5172 36641
rect 5206 36607 5244 36641
rect 5278 36607 5284 36641
rect 5166 36568 5284 36607
rect 5166 36534 5172 36568
rect 5206 36534 5244 36568
rect 5278 36534 5284 36568
rect 5166 36495 5284 36534
rect 5166 36461 5172 36495
rect 5206 36461 5244 36495
rect 5278 36461 5284 36495
rect 5166 36422 5284 36461
rect 5166 35892 5172 36422
rect 5278 35892 5284 36422
rect 5166 35826 5172 35840
rect 5278 35826 5284 35840
rect 5166 35760 5172 35774
rect 5278 35760 5284 35774
rect 5166 35694 5172 35708
rect 5278 35694 5284 35708
rect 5166 35627 5172 35642
rect 5278 35627 5284 35642
rect 5166 35560 5172 35575
rect 5278 35560 5284 35575
rect 5166 35493 5172 35508
rect 5278 35493 5284 35508
rect 5166 35426 5172 35441
rect 5278 35426 5284 35441
rect 5218 35374 5232 35380
tri 4730 35280 4774 35324 sw
tri 5122 35280 5166 35324 se
rect 5166 35280 5284 35374
rect 5443 38720 5561 38726
rect 5495 38668 5509 38720
rect 5443 38654 5561 38668
rect 5495 38602 5509 38654
rect 5443 38588 5561 38602
rect 5495 38536 5509 38588
rect 5443 38534 5449 38536
rect 5483 38534 5521 38536
rect 5555 38534 5561 38536
rect 5443 38522 5561 38534
rect 5495 38470 5509 38522
rect 5443 38461 5449 38470
rect 5483 38461 5521 38470
rect 5555 38461 5561 38470
rect 5443 38456 5561 38461
rect 5495 38422 5509 38456
rect 5443 38390 5449 38404
rect 5555 38390 5561 38404
rect 5443 38323 5449 38338
rect 5555 38323 5561 38338
rect 5443 38256 5449 38271
rect 5555 38256 5561 38271
rect 5443 37380 5449 38204
rect 5555 37380 5561 38204
rect 5443 36720 5561 37380
rect 5495 36668 5509 36720
rect 5443 36654 5561 36668
rect 5495 36602 5509 36654
rect 5443 36588 5561 36602
rect 5495 36536 5509 36588
rect 5443 36534 5449 36536
rect 5483 36534 5521 36536
rect 5555 36534 5561 36536
rect 5443 36522 5561 36534
rect 5495 36470 5509 36522
rect 5443 36461 5449 36470
rect 5483 36461 5521 36470
rect 5555 36461 5561 36470
rect 5443 36456 5561 36461
rect 5495 36422 5509 36456
rect 5443 36390 5449 36404
rect 5555 36390 5561 36404
rect 5443 36323 5449 36338
rect 5555 36323 5561 36338
rect 5443 36256 5449 36271
rect 5555 36256 5561 36271
rect 5443 35380 5449 36204
rect 5555 35380 5561 36204
rect 5443 35368 5561 35380
rect 5720 38714 5838 38726
rect 5720 38680 5726 38714
rect 5760 38680 5798 38714
rect 5832 38680 5838 38714
rect 5720 38641 5838 38680
rect 5720 38607 5726 38641
rect 5760 38607 5798 38641
rect 5832 38607 5838 38641
rect 5720 38568 5838 38607
rect 5720 38534 5726 38568
rect 5760 38534 5798 38568
rect 5832 38534 5838 38568
rect 5720 38495 5838 38534
rect 5720 38461 5726 38495
rect 5760 38461 5798 38495
rect 5832 38461 5838 38495
rect 5720 38422 5838 38461
rect 5720 37892 5726 38422
rect 5832 37892 5838 38422
rect 5720 37825 5726 37840
rect 5832 37825 5838 37840
rect 5720 37758 5726 37773
rect 5832 37758 5838 37773
rect 5720 37691 5726 37706
rect 5832 37691 5838 37706
rect 5720 37624 5726 37639
rect 5832 37624 5838 37639
rect 5720 37557 5726 37572
rect 5832 37557 5838 37572
rect 5720 37490 5726 37505
rect 5832 37490 5838 37505
rect 5720 37423 5726 37438
rect 5832 37423 5838 37438
rect 5772 37371 5786 37380
rect 5720 37356 5838 37371
rect 5772 37304 5786 37356
rect 5720 37289 5838 37304
rect 5772 37237 5786 37289
rect 5720 37222 5838 37237
rect 5772 37170 5786 37222
rect 5720 37155 5838 37170
rect 5772 37103 5786 37155
rect 5720 37088 5838 37103
rect 5772 37036 5786 37088
rect 5720 36714 5838 37036
rect 5720 36680 5726 36714
rect 5760 36680 5798 36714
rect 5832 36680 5838 36714
rect 5720 36641 5838 36680
rect 5720 36607 5726 36641
rect 5760 36607 5798 36641
rect 5832 36607 5838 36641
rect 5720 36568 5838 36607
rect 5720 36534 5726 36568
rect 5760 36534 5798 36568
rect 5832 36534 5838 36568
rect 5720 36495 5838 36534
rect 5720 36461 5726 36495
rect 5760 36461 5798 36495
rect 5832 36461 5838 36495
rect 5720 36422 5838 36461
rect 5720 35892 5726 36422
rect 5832 35892 5838 36422
rect 5720 35826 5726 35840
rect 5832 35826 5838 35840
rect 5720 35760 5726 35774
rect 5832 35760 5838 35774
rect 5720 35694 5726 35708
rect 5832 35694 5838 35708
rect 5720 35627 5726 35642
rect 5832 35627 5838 35642
rect 5720 35560 5726 35575
rect 5832 35560 5838 35575
rect 5720 35493 5726 35508
rect 5832 35493 5838 35508
rect 5720 35426 5726 35441
rect 5832 35426 5838 35441
rect 5772 35374 5786 35380
tri 5284 35280 5328 35324 sw
tri 5676 35280 5720 35324 se
rect 5720 35280 5838 35374
rect 5997 38720 6115 38726
rect 6049 38668 6063 38720
rect 5997 38654 6115 38668
rect 6049 38602 6063 38654
rect 5997 38588 6115 38602
rect 6049 38536 6063 38588
rect 5997 38534 6003 38536
rect 6037 38534 6075 38536
rect 6109 38534 6115 38536
rect 5997 38522 6115 38534
rect 6049 38470 6063 38522
rect 5997 38461 6003 38470
rect 6037 38461 6075 38470
rect 6109 38461 6115 38470
rect 5997 38456 6115 38461
rect 6049 38422 6063 38456
rect 5997 38390 6003 38404
rect 6109 38390 6115 38404
rect 5997 38323 6003 38338
rect 6109 38323 6115 38338
rect 5997 38256 6003 38271
rect 6109 38256 6115 38271
rect 5997 37380 6003 38204
rect 6109 37380 6115 38204
rect 5997 36720 6115 37380
rect 6049 36668 6063 36720
rect 5997 36654 6115 36668
rect 6049 36602 6063 36654
rect 5997 36588 6115 36602
rect 6049 36536 6063 36588
rect 5997 36534 6003 36536
rect 6037 36534 6075 36536
rect 6109 36534 6115 36536
rect 5997 36522 6115 36534
rect 6049 36470 6063 36522
rect 5997 36461 6003 36470
rect 6037 36461 6075 36470
rect 6109 36461 6115 36470
rect 5997 36456 6115 36461
rect 6049 36422 6063 36456
rect 5997 36390 6003 36404
rect 6109 36390 6115 36404
rect 5997 36323 6003 36338
rect 6109 36323 6115 36338
rect 5997 36256 6003 36271
rect 6109 36256 6115 36271
rect 5997 35380 6003 36204
rect 6109 35380 6115 36204
rect 5997 35368 6115 35380
rect 6274 38714 6392 38726
rect 6274 38680 6280 38714
rect 6314 38680 6352 38714
rect 6386 38680 6392 38714
rect 6274 38641 6392 38680
rect 6274 38607 6280 38641
rect 6314 38607 6352 38641
rect 6386 38607 6392 38641
rect 6274 38568 6392 38607
rect 6274 38534 6280 38568
rect 6314 38534 6352 38568
rect 6386 38534 6392 38568
rect 6274 38495 6392 38534
rect 6274 38461 6280 38495
rect 6314 38461 6352 38495
rect 6386 38461 6392 38495
rect 6274 38422 6392 38461
rect 6274 37892 6280 38422
rect 6386 37892 6392 38422
rect 6274 37825 6280 37840
rect 6386 37825 6392 37840
rect 6274 37758 6280 37773
rect 6386 37758 6392 37773
rect 6274 37691 6280 37706
rect 6386 37691 6392 37706
rect 6274 37624 6280 37639
rect 6386 37624 6392 37639
rect 6274 37557 6280 37572
rect 6386 37557 6392 37572
rect 6274 37490 6280 37505
rect 6386 37490 6392 37505
rect 6274 37423 6280 37438
rect 6386 37423 6392 37438
rect 6326 37371 6340 37380
rect 6274 37356 6392 37371
rect 6326 37304 6340 37356
rect 6274 37289 6392 37304
rect 6326 37237 6340 37289
rect 6274 37222 6392 37237
rect 6326 37170 6340 37222
rect 6274 37155 6392 37170
rect 6326 37103 6340 37155
rect 6274 37088 6392 37103
rect 6326 37036 6340 37088
rect 6274 36714 6392 37036
rect 6274 36680 6280 36714
rect 6314 36680 6352 36714
rect 6386 36680 6392 36714
rect 6274 36641 6392 36680
rect 6274 36607 6280 36641
rect 6314 36607 6352 36641
rect 6386 36607 6392 36641
rect 6274 36568 6392 36607
rect 6274 36534 6280 36568
rect 6314 36534 6352 36568
rect 6386 36534 6392 36568
rect 6274 36495 6392 36534
rect 6274 36461 6280 36495
rect 6314 36461 6352 36495
rect 6386 36461 6392 36495
rect 6274 36422 6392 36461
rect 6274 35892 6280 36422
rect 6386 35892 6392 36422
rect 6274 35826 6280 35840
rect 6386 35826 6392 35840
rect 6274 35760 6280 35774
rect 6386 35760 6392 35774
rect 6274 35694 6280 35708
rect 6386 35694 6392 35708
rect 6274 35627 6280 35642
rect 6386 35627 6392 35642
rect 6274 35560 6280 35575
rect 6386 35560 6392 35575
rect 6274 35493 6280 35508
rect 6386 35493 6392 35508
rect 6274 35426 6280 35441
rect 6386 35426 6392 35441
rect 6326 35374 6340 35380
tri 5838 35280 5882 35324 sw
tri 6230 35280 6274 35324 se
rect 6274 35280 6392 35374
rect 6551 38720 6669 38726
rect 6603 38668 6617 38720
rect 6551 38654 6669 38668
rect 6603 38602 6617 38654
rect 6551 38588 6669 38602
rect 6603 38536 6617 38588
rect 6551 38534 6557 38536
rect 6591 38534 6629 38536
rect 6663 38534 6669 38536
rect 6551 38522 6669 38534
rect 6603 38470 6617 38522
rect 6551 38461 6557 38470
rect 6591 38461 6629 38470
rect 6663 38461 6669 38470
rect 6551 38456 6669 38461
rect 6603 38422 6617 38456
rect 6551 38390 6557 38404
rect 6663 38390 6669 38404
rect 6551 38323 6557 38338
rect 6663 38323 6669 38338
rect 6551 38256 6557 38271
rect 6663 38256 6669 38271
rect 6551 37380 6557 38204
rect 6663 37380 6669 38204
rect 6551 36720 6669 37380
rect 6603 36668 6617 36720
rect 6551 36654 6669 36668
rect 6603 36602 6617 36654
rect 6551 36588 6669 36602
rect 6603 36536 6617 36588
rect 6551 36534 6557 36536
rect 6591 36534 6629 36536
rect 6663 36534 6669 36536
rect 6551 36522 6669 36534
rect 6603 36470 6617 36522
rect 6551 36461 6557 36470
rect 6591 36461 6629 36470
rect 6663 36461 6669 36470
rect 6551 36456 6669 36461
rect 6603 36422 6617 36456
rect 6551 36390 6557 36404
rect 6663 36390 6669 36404
rect 6551 36323 6557 36338
rect 6663 36323 6669 36338
rect 6551 36256 6557 36271
rect 6663 36256 6669 36271
rect 6551 35380 6557 36204
rect 6663 35380 6669 36204
rect 6551 35368 6669 35380
rect 6828 38714 6946 38726
rect 6828 38680 6834 38714
rect 6868 38680 6906 38714
rect 6940 38680 6946 38714
rect 6828 38641 6946 38680
rect 6828 38607 6834 38641
rect 6868 38607 6906 38641
rect 6940 38607 6946 38641
rect 6828 38568 6946 38607
rect 6828 38534 6834 38568
rect 6868 38534 6906 38568
rect 6940 38534 6946 38568
rect 6828 38495 6946 38534
rect 6828 38461 6834 38495
rect 6868 38461 6906 38495
rect 6940 38461 6946 38495
rect 6828 38422 6946 38461
rect 6828 37892 6834 38422
rect 6940 37892 6946 38422
rect 6828 37825 6834 37840
rect 6940 37825 6946 37840
rect 6828 37758 6834 37773
rect 6940 37758 6946 37773
rect 6828 37691 6834 37706
rect 6940 37691 6946 37706
rect 6828 37624 6834 37639
rect 6940 37624 6946 37639
rect 6828 37557 6834 37572
rect 6940 37557 6946 37572
rect 6828 37490 6834 37505
rect 6940 37490 6946 37505
rect 6828 37423 6834 37438
rect 6940 37423 6946 37438
rect 6880 37371 6894 37380
rect 6828 37356 6946 37371
rect 6880 37304 6894 37356
rect 6828 37289 6946 37304
rect 6880 37237 6894 37289
rect 6828 37222 6946 37237
rect 6880 37170 6894 37222
rect 6828 37155 6946 37170
rect 6880 37103 6894 37155
rect 6828 37088 6946 37103
rect 6880 37036 6894 37088
rect 6828 36714 6946 37036
rect 6828 36680 6834 36714
rect 6868 36680 6906 36714
rect 6940 36680 6946 36714
rect 6828 36641 6946 36680
rect 6828 36607 6834 36641
rect 6868 36607 6906 36641
rect 6940 36607 6946 36641
rect 6828 36568 6946 36607
rect 6828 36534 6834 36568
rect 6868 36534 6906 36568
rect 6940 36534 6946 36568
rect 6828 36495 6946 36534
rect 6828 36461 6834 36495
rect 6868 36461 6906 36495
rect 6940 36461 6946 36495
rect 6828 36422 6946 36461
rect 6828 35892 6834 36422
rect 6940 35892 6946 36422
rect 6828 35826 6834 35840
rect 6940 35826 6946 35840
rect 6828 35760 6834 35774
rect 6940 35760 6946 35774
rect 6828 35694 6834 35708
rect 6940 35694 6946 35708
rect 6828 35627 6834 35642
rect 6940 35627 6946 35642
rect 6828 35560 6834 35575
rect 6940 35560 6946 35575
rect 6828 35493 6834 35508
rect 6940 35493 6946 35508
rect 6828 35426 6834 35441
rect 6940 35426 6946 35441
rect 6880 35374 6894 35380
tri 6392 35280 6436 35324 sw
tri 6784 35280 6828 35324 se
rect 6828 35280 6946 35374
rect 7105 38720 7223 38726
rect 7157 38668 7171 38720
rect 7105 38654 7223 38668
rect 7157 38602 7171 38654
rect 7105 38588 7223 38602
rect 7157 38536 7171 38588
rect 7105 38534 7111 38536
rect 7145 38534 7183 38536
rect 7217 38534 7223 38536
rect 7105 38522 7223 38534
rect 7157 38470 7171 38522
rect 7105 38461 7111 38470
rect 7145 38461 7183 38470
rect 7217 38461 7223 38470
rect 7105 38456 7223 38461
rect 7157 38422 7171 38456
rect 7105 38390 7111 38404
rect 7217 38390 7223 38404
rect 7105 38323 7111 38338
rect 7217 38323 7223 38338
rect 7105 38256 7111 38271
rect 7217 38256 7223 38271
rect 7105 37380 7111 38204
rect 7217 37380 7223 38204
rect 7105 36720 7223 37380
rect 7157 36668 7171 36720
rect 7105 36654 7223 36668
rect 7157 36602 7171 36654
rect 7105 36588 7223 36602
rect 7157 36536 7171 36588
rect 7105 36534 7111 36536
rect 7145 36534 7183 36536
rect 7217 36534 7223 36536
rect 7105 36522 7223 36534
rect 7157 36470 7171 36522
rect 7105 36461 7111 36470
rect 7145 36461 7183 36470
rect 7217 36461 7223 36470
rect 7105 36456 7223 36461
rect 7157 36422 7171 36456
rect 7105 36390 7111 36404
rect 7217 36390 7223 36404
rect 7105 36323 7111 36338
rect 7217 36323 7223 36338
rect 7105 36256 7111 36271
rect 7217 36256 7223 36271
rect 7105 35380 7111 36204
rect 7217 35380 7223 36204
rect 7105 35368 7223 35380
rect 7382 38714 7500 38726
rect 7382 38680 7388 38714
rect 7422 38680 7460 38714
rect 7494 38680 7500 38714
rect 7382 38641 7500 38680
rect 7382 38607 7388 38641
rect 7422 38607 7460 38641
rect 7494 38607 7500 38641
rect 7382 38568 7500 38607
rect 7382 38534 7388 38568
rect 7422 38534 7460 38568
rect 7494 38534 7500 38568
rect 7382 38495 7500 38534
rect 7382 38461 7388 38495
rect 7422 38461 7460 38495
rect 7494 38461 7500 38495
rect 7382 38422 7500 38461
rect 7382 37892 7388 38422
rect 7494 37892 7500 38422
rect 7382 37825 7388 37840
rect 7494 37825 7500 37840
rect 7382 37758 7388 37773
rect 7494 37758 7500 37773
rect 7382 37691 7388 37706
rect 7494 37691 7500 37706
rect 7382 37624 7388 37639
rect 7494 37624 7500 37639
rect 7382 37557 7388 37572
rect 7494 37557 7500 37572
rect 7382 37490 7388 37505
rect 7494 37490 7500 37505
rect 7382 37423 7388 37438
rect 7494 37423 7500 37438
rect 7434 37371 7448 37380
rect 7382 37356 7500 37371
rect 7434 37304 7448 37356
rect 7382 37289 7500 37304
rect 7434 37237 7448 37289
rect 7382 37222 7500 37237
rect 7434 37170 7448 37222
rect 7382 37155 7500 37170
rect 7434 37103 7448 37155
rect 7382 37088 7500 37103
rect 7434 37036 7448 37088
rect 7382 36714 7500 37036
rect 7382 36680 7388 36714
rect 7422 36680 7460 36714
rect 7494 36680 7500 36714
rect 7382 36641 7500 36680
rect 7382 36607 7388 36641
rect 7422 36607 7460 36641
rect 7494 36607 7500 36641
rect 7382 36568 7500 36607
rect 7382 36534 7388 36568
rect 7422 36534 7460 36568
rect 7494 36534 7500 36568
rect 7382 36495 7500 36534
rect 7382 36461 7388 36495
rect 7422 36461 7460 36495
rect 7494 36461 7500 36495
rect 7382 36422 7500 36461
rect 7382 35892 7388 36422
rect 7494 35892 7500 36422
rect 7382 35826 7388 35840
rect 7494 35826 7500 35840
rect 7382 35760 7388 35774
rect 7494 35760 7500 35774
rect 7382 35694 7388 35708
rect 7494 35694 7500 35708
rect 7382 35627 7388 35642
rect 7494 35627 7500 35642
rect 7382 35560 7388 35575
rect 7494 35560 7500 35575
rect 7382 35493 7388 35508
rect 7494 35493 7500 35508
rect 7382 35426 7388 35441
rect 7494 35426 7500 35441
rect 7434 35374 7448 35380
tri 6946 35280 6990 35324 sw
tri 7338 35280 7382 35324 se
rect 7382 35280 7500 35374
rect 7659 38720 7777 38726
rect 7711 38668 7725 38720
rect 7659 38654 7777 38668
rect 7711 38602 7725 38654
rect 7659 38588 7777 38602
rect 7711 38536 7725 38588
rect 7659 38534 7665 38536
rect 7699 38534 7737 38536
rect 7771 38534 7777 38536
rect 7659 38522 7777 38534
rect 7711 38470 7725 38522
rect 7659 38461 7665 38470
rect 7699 38461 7737 38470
rect 7771 38461 7777 38470
rect 7659 38456 7777 38461
rect 7711 38422 7725 38456
rect 7659 38390 7665 38404
rect 7771 38390 7777 38404
rect 7659 38323 7665 38338
rect 7771 38323 7777 38338
rect 7659 38256 7665 38271
rect 7771 38256 7777 38271
rect 7659 37380 7665 38204
rect 7771 37380 7777 38204
rect 7659 36720 7777 37380
rect 7711 36668 7725 36720
rect 7659 36654 7777 36668
rect 7711 36602 7725 36654
rect 7659 36588 7777 36602
rect 7711 36536 7725 36588
rect 7659 36534 7665 36536
rect 7699 36534 7737 36536
rect 7771 36534 7777 36536
rect 7659 36522 7777 36534
rect 7711 36470 7725 36522
rect 7659 36461 7665 36470
rect 7699 36461 7737 36470
rect 7771 36461 7777 36470
rect 7659 36456 7777 36461
rect 7711 36422 7725 36456
rect 7659 36390 7665 36404
rect 7771 36390 7777 36404
rect 7659 36323 7665 36338
rect 7771 36323 7777 36338
rect 7659 36256 7665 36271
rect 7771 36256 7777 36271
rect 7659 35380 7665 36204
rect 7771 35380 7777 36204
rect 7659 35368 7777 35380
rect 7936 38714 8054 38726
rect 7936 38680 7942 38714
rect 7976 38680 8014 38714
rect 8048 38680 8054 38714
rect 7936 38641 8054 38680
rect 7936 38607 7942 38641
rect 7976 38607 8014 38641
rect 8048 38607 8054 38641
rect 7936 38568 8054 38607
rect 7936 38534 7942 38568
rect 7976 38534 8014 38568
rect 8048 38534 8054 38568
rect 7936 38495 8054 38534
rect 7936 38461 7942 38495
rect 7976 38461 8014 38495
rect 8048 38461 8054 38495
rect 7936 38422 8054 38461
rect 7936 37892 7942 38422
rect 8048 37892 8054 38422
rect 7936 37825 7942 37840
rect 8048 37825 8054 37840
rect 7936 37758 7942 37773
rect 8048 37758 8054 37773
rect 7936 37691 7942 37706
rect 8048 37691 8054 37706
rect 7936 37624 7942 37639
rect 8048 37624 8054 37639
rect 7936 37557 7942 37572
rect 8048 37557 8054 37572
rect 7936 37490 7942 37505
rect 8048 37490 8054 37505
rect 7936 37423 7942 37438
rect 8048 37423 8054 37438
rect 7988 37371 8002 37380
rect 7936 37356 8054 37371
rect 7988 37304 8002 37356
rect 7936 37289 8054 37304
rect 7988 37237 8002 37289
rect 7936 37222 8054 37237
rect 7988 37170 8002 37222
rect 7936 37155 8054 37170
rect 7988 37103 8002 37155
rect 7936 37088 8054 37103
rect 7988 37036 8002 37088
rect 7936 36714 8054 37036
rect 7936 36680 7942 36714
rect 7976 36680 8014 36714
rect 8048 36680 8054 36714
rect 7936 36641 8054 36680
rect 7936 36607 7942 36641
rect 7976 36607 8014 36641
rect 8048 36607 8054 36641
rect 7936 36568 8054 36607
rect 7936 36534 7942 36568
rect 7976 36534 8014 36568
rect 8048 36534 8054 36568
rect 7936 36495 8054 36534
rect 7936 36461 7942 36495
rect 7976 36461 8014 36495
rect 8048 36461 8054 36495
rect 7936 36422 8054 36461
rect 7936 35892 7942 36422
rect 8048 35892 8054 36422
rect 7936 35826 7942 35840
rect 8048 35826 8054 35840
rect 7936 35760 7942 35774
rect 8048 35760 8054 35774
rect 7936 35694 7942 35708
rect 8048 35694 8054 35708
rect 7936 35627 7942 35642
rect 8048 35627 8054 35642
rect 7936 35560 7942 35575
rect 8048 35560 8054 35575
rect 7936 35493 7942 35508
rect 8048 35493 8054 35508
rect 7936 35426 7942 35441
rect 8048 35426 8054 35441
rect 7988 35374 8002 35380
tri 7500 35280 7544 35324 sw
tri 7892 35280 7936 35324 se
rect 7936 35280 8054 35374
rect 8213 38720 8331 38726
rect 8265 38668 8279 38720
rect 8213 38654 8331 38668
rect 8265 38602 8279 38654
rect 8213 38588 8331 38602
rect 8265 38536 8279 38588
rect 8213 38534 8219 38536
rect 8253 38534 8291 38536
rect 8325 38534 8331 38536
rect 8213 38522 8331 38534
rect 8265 38470 8279 38522
rect 8213 38461 8219 38470
rect 8253 38461 8291 38470
rect 8325 38461 8331 38470
rect 8213 38456 8331 38461
rect 8265 38422 8279 38456
rect 8213 38390 8219 38404
rect 8325 38390 8331 38404
rect 8213 38323 8219 38338
rect 8325 38323 8331 38338
rect 8213 38256 8219 38271
rect 8325 38256 8331 38271
rect 8213 37380 8219 38204
rect 8325 37380 8331 38204
rect 8213 36720 8331 37380
rect 8265 36668 8279 36720
rect 8213 36654 8331 36668
rect 8265 36602 8279 36654
rect 8213 36588 8331 36602
rect 8265 36536 8279 36588
rect 8213 36534 8219 36536
rect 8253 36534 8291 36536
rect 8325 36534 8331 36536
rect 8213 36522 8331 36534
rect 8265 36470 8279 36522
rect 8213 36461 8219 36470
rect 8253 36461 8291 36470
rect 8325 36461 8331 36470
rect 8213 36456 8331 36461
rect 8265 36422 8279 36456
rect 8213 36390 8219 36404
rect 8325 36390 8331 36404
rect 8213 36323 8219 36338
rect 8325 36323 8331 36338
rect 8213 36256 8219 36271
rect 8325 36256 8331 36271
rect 8213 35380 8219 36204
rect 8325 35380 8331 36204
rect 8213 35368 8331 35380
rect 8490 38714 8608 38726
rect 8490 38680 8496 38714
rect 8530 38680 8568 38714
rect 8602 38680 8608 38714
rect 8490 38641 8608 38680
rect 8490 38607 8496 38641
rect 8530 38607 8568 38641
rect 8602 38607 8608 38641
rect 8490 38568 8608 38607
rect 8490 38534 8496 38568
rect 8530 38534 8568 38568
rect 8602 38534 8608 38568
rect 8490 38495 8608 38534
rect 8490 38461 8496 38495
rect 8530 38461 8568 38495
rect 8602 38461 8608 38495
rect 8490 38422 8608 38461
rect 8490 37892 8496 38422
rect 8602 37892 8608 38422
rect 8490 37825 8496 37840
rect 8602 37825 8608 37840
rect 8490 37758 8496 37773
rect 8602 37758 8608 37773
rect 8490 37691 8496 37706
rect 8602 37691 8608 37706
rect 8490 37624 8496 37639
rect 8602 37624 8608 37639
rect 8490 37557 8496 37572
rect 8602 37557 8608 37572
rect 8490 37490 8496 37505
rect 8602 37490 8608 37505
rect 8490 37423 8496 37438
rect 8602 37423 8608 37438
rect 8542 37371 8556 37380
rect 8490 37356 8608 37371
rect 8542 37304 8556 37356
rect 8490 37289 8608 37304
rect 8542 37237 8556 37289
rect 8490 37222 8608 37237
rect 8542 37170 8556 37222
rect 8490 37155 8608 37170
rect 8542 37103 8556 37155
rect 8490 37088 8608 37103
rect 8542 37036 8556 37088
rect 8490 36714 8608 37036
rect 8490 36680 8496 36714
rect 8530 36680 8568 36714
rect 8602 36680 8608 36714
rect 8490 36641 8608 36680
rect 8490 36607 8496 36641
rect 8530 36607 8568 36641
rect 8602 36607 8608 36641
rect 8490 36568 8608 36607
rect 8490 36534 8496 36568
rect 8530 36534 8568 36568
rect 8602 36534 8608 36568
rect 8490 36495 8608 36534
rect 8490 36461 8496 36495
rect 8530 36461 8568 36495
rect 8602 36461 8608 36495
rect 8490 36422 8608 36461
rect 8490 35892 8496 36422
rect 8602 35892 8608 36422
rect 8490 35826 8496 35840
rect 8602 35826 8608 35840
rect 8490 35760 8496 35774
rect 8602 35760 8608 35774
rect 8490 35694 8496 35708
rect 8602 35694 8608 35708
rect 8490 35627 8496 35642
rect 8602 35627 8608 35642
rect 8490 35560 8496 35575
rect 8602 35560 8608 35575
rect 8490 35493 8496 35508
rect 8602 35493 8608 35508
rect 8490 35426 8496 35441
rect 8602 35426 8608 35441
rect 8542 35374 8556 35380
tri 8054 35280 8098 35324 sw
tri 8446 35280 8490 35324 se
rect 8490 35280 8608 35374
rect 8767 38720 8885 38726
rect 8819 38668 8833 38720
rect 8767 38654 8885 38668
rect 8819 38602 8833 38654
rect 8767 38588 8885 38602
rect 8819 38536 8833 38588
rect 8767 38534 8773 38536
rect 8807 38534 8845 38536
rect 8879 38534 8885 38536
rect 8767 38522 8885 38534
rect 8819 38470 8833 38522
rect 8767 38461 8773 38470
rect 8807 38461 8845 38470
rect 8879 38461 8885 38470
rect 8767 38456 8885 38461
rect 8819 38422 8833 38456
rect 8767 38390 8773 38404
rect 8879 38390 8885 38404
rect 8767 38323 8773 38338
rect 8879 38323 8885 38338
rect 8767 38256 8773 38271
rect 8879 38256 8885 38271
rect 8767 37380 8773 38204
rect 8879 37380 8885 38204
rect 8767 36720 8885 37380
rect 8819 36668 8833 36720
rect 8767 36654 8885 36668
rect 8819 36602 8833 36654
rect 8767 36588 8885 36602
rect 8819 36536 8833 36588
rect 8767 36534 8773 36536
rect 8807 36534 8845 36536
rect 8879 36534 8885 36536
rect 8767 36522 8885 36534
rect 8819 36470 8833 36522
rect 8767 36461 8773 36470
rect 8807 36461 8845 36470
rect 8879 36461 8885 36470
rect 8767 36456 8885 36461
rect 8819 36422 8833 36456
rect 8767 36390 8773 36404
rect 8879 36390 8885 36404
rect 8767 36323 8773 36338
rect 8879 36323 8885 36338
rect 8767 36256 8773 36271
rect 8879 36256 8885 36271
rect 8767 35380 8773 36204
rect 8879 35380 8885 36204
rect 8767 35368 8885 35380
rect 9044 38714 9162 38726
rect 9044 38680 9050 38714
rect 9084 38680 9122 38714
rect 9156 38680 9162 38714
rect 9044 38641 9162 38680
rect 9044 38607 9050 38641
rect 9084 38607 9122 38641
rect 9156 38607 9162 38641
rect 9044 38568 9162 38607
rect 9044 38534 9050 38568
rect 9084 38534 9122 38568
rect 9156 38534 9162 38568
rect 9044 38495 9162 38534
rect 9044 38461 9050 38495
rect 9084 38461 9122 38495
rect 9156 38461 9162 38495
rect 9044 38422 9162 38461
rect 9044 37892 9050 38422
rect 9156 37892 9162 38422
rect 9044 37825 9050 37840
rect 9156 37825 9162 37840
rect 9044 37758 9050 37773
rect 9156 37758 9162 37773
rect 9044 37691 9050 37706
rect 9156 37691 9162 37706
rect 9044 37624 9050 37639
rect 9156 37624 9162 37639
rect 9044 37557 9050 37572
rect 9156 37557 9162 37572
rect 9044 37490 9050 37505
rect 9156 37490 9162 37505
rect 9044 37423 9050 37438
rect 9156 37423 9162 37438
rect 9096 37371 9110 37380
rect 9044 37356 9162 37371
rect 9096 37304 9110 37356
rect 9044 37289 9162 37304
rect 9096 37237 9110 37289
rect 9044 37222 9162 37237
rect 9096 37170 9110 37222
rect 9044 37155 9162 37170
rect 9096 37103 9110 37155
rect 9044 37088 9162 37103
rect 9096 37036 9110 37088
rect 9044 36714 9162 37036
rect 9044 36680 9050 36714
rect 9084 36680 9122 36714
rect 9156 36680 9162 36714
rect 9044 36641 9162 36680
rect 9044 36607 9050 36641
rect 9084 36607 9122 36641
rect 9156 36607 9162 36641
rect 9044 36568 9162 36607
rect 9044 36534 9050 36568
rect 9084 36534 9122 36568
rect 9156 36534 9162 36568
rect 9044 36495 9162 36534
rect 9044 36461 9050 36495
rect 9084 36461 9122 36495
rect 9156 36461 9162 36495
rect 9044 36422 9162 36461
rect 9044 35892 9050 36422
rect 9156 35892 9162 36422
rect 9044 35826 9050 35840
rect 9156 35826 9162 35840
rect 9044 35760 9050 35774
rect 9156 35760 9162 35774
rect 9044 35694 9050 35708
rect 9156 35694 9162 35708
rect 9044 35627 9050 35642
rect 9156 35627 9162 35642
rect 9044 35560 9050 35575
rect 9156 35560 9162 35575
rect 9044 35493 9050 35508
rect 9156 35493 9162 35508
rect 9044 35426 9050 35441
rect 9156 35426 9162 35441
rect 9096 35374 9110 35380
tri 8608 35280 8652 35324 sw
tri 9000 35280 9044 35324 se
rect 9044 35280 9162 35374
rect 9321 38720 9439 38726
rect 9373 38668 9387 38720
rect 9321 38654 9439 38668
rect 9373 38602 9387 38654
rect 9321 38588 9439 38602
rect 9373 38536 9387 38588
rect 9321 38534 9327 38536
rect 9361 38534 9399 38536
rect 9433 38534 9439 38536
rect 9321 38522 9439 38534
rect 9373 38470 9387 38522
rect 9321 38461 9327 38470
rect 9361 38461 9399 38470
rect 9433 38461 9439 38470
rect 9321 38456 9439 38461
rect 9373 38422 9387 38456
rect 9321 38390 9327 38404
rect 9433 38390 9439 38404
rect 9321 38323 9327 38338
rect 9433 38323 9439 38338
rect 9321 38256 9327 38271
rect 9433 38256 9439 38271
rect 9321 37380 9327 38204
rect 9433 37380 9439 38204
rect 9321 36720 9439 37380
rect 9373 36668 9387 36720
rect 9321 36654 9439 36668
rect 9373 36602 9387 36654
rect 9321 36588 9439 36602
rect 9373 36536 9387 36588
rect 9321 36534 9327 36536
rect 9361 36534 9399 36536
rect 9433 36534 9439 36536
rect 9321 36522 9439 36534
rect 9373 36470 9387 36522
rect 9321 36461 9327 36470
rect 9361 36461 9399 36470
rect 9433 36461 9439 36470
rect 9321 36456 9439 36461
rect 9373 36422 9387 36456
rect 9321 36390 9327 36404
rect 9433 36390 9439 36404
rect 9321 36323 9327 36338
rect 9433 36323 9439 36338
rect 9321 36256 9327 36271
rect 9433 36256 9439 36271
rect 9321 35380 9327 36204
rect 9433 35380 9439 36204
rect 9321 35368 9439 35380
rect 9598 38714 9716 38726
rect 9598 38680 9604 38714
rect 9638 38680 9676 38714
rect 9710 38680 9716 38714
rect 9598 38641 9716 38680
rect 9598 38607 9604 38641
rect 9638 38607 9676 38641
rect 9710 38607 9716 38641
rect 9598 38568 9716 38607
rect 9598 38534 9604 38568
rect 9638 38534 9676 38568
rect 9710 38534 9716 38568
rect 9598 38495 9716 38534
rect 9598 38461 9604 38495
rect 9638 38461 9676 38495
rect 9710 38461 9716 38495
rect 9598 38422 9716 38461
rect 9598 37892 9604 38422
rect 9710 37892 9716 38422
rect 9598 37825 9604 37840
rect 9710 37825 9716 37840
rect 9598 37758 9604 37773
rect 9710 37758 9716 37773
rect 9598 37691 9604 37706
rect 9710 37691 9716 37706
rect 9598 37624 9604 37639
rect 9710 37624 9716 37639
rect 9598 37557 9604 37572
rect 9710 37557 9716 37572
rect 9598 37490 9604 37505
rect 9710 37490 9716 37505
rect 9598 37423 9604 37438
rect 9710 37423 9716 37438
rect 9650 37371 9664 37380
rect 9598 37356 9716 37371
rect 9650 37304 9664 37356
rect 9598 37289 9716 37304
rect 9650 37237 9664 37289
rect 9598 37222 9716 37237
rect 9650 37170 9664 37222
rect 9598 37155 9716 37170
rect 9650 37103 9664 37155
rect 9598 37088 9716 37103
rect 9650 37036 9664 37088
rect 9598 36714 9716 37036
rect 9598 36680 9604 36714
rect 9638 36680 9676 36714
rect 9710 36680 9716 36714
rect 9598 36641 9716 36680
rect 9598 36607 9604 36641
rect 9638 36607 9676 36641
rect 9710 36607 9716 36641
rect 9598 36568 9716 36607
rect 9598 36534 9604 36568
rect 9638 36534 9676 36568
rect 9710 36534 9716 36568
rect 9598 36495 9716 36534
rect 9598 36461 9604 36495
rect 9638 36461 9676 36495
rect 9710 36461 9716 36495
rect 9598 36422 9716 36461
rect 9598 35892 9604 36422
rect 9710 35892 9716 36422
rect 9598 35826 9604 35840
rect 9710 35826 9716 35840
rect 9598 35760 9604 35774
rect 9710 35760 9716 35774
rect 9598 35694 9604 35708
rect 9710 35694 9716 35708
rect 9598 35627 9604 35642
rect 9710 35627 9716 35642
rect 9598 35560 9604 35575
rect 9710 35560 9716 35575
rect 9598 35493 9604 35508
rect 9710 35493 9716 35508
rect 9598 35426 9604 35441
rect 9710 35426 9716 35441
rect 9650 35374 9664 35380
tri 9162 35280 9206 35324 sw
tri 9554 35280 9598 35324 se
rect 9598 35280 9716 35374
rect 9875 38720 9993 38726
rect 9927 38668 9941 38720
rect 9875 38654 9993 38668
rect 9927 38602 9941 38654
rect 9875 38588 9993 38602
rect 9927 38536 9941 38588
rect 9875 38534 9881 38536
rect 9915 38534 9953 38536
rect 9987 38534 9993 38536
rect 9875 38522 9993 38534
rect 9927 38470 9941 38522
rect 9875 38461 9881 38470
rect 9915 38461 9953 38470
rect 9987 38461 9993 38470
rect 9875 38456 9993 38461
rect 9927 38422 9941 38456
rect 9875 38390 9881 38404
rect 9987 38390 9993 38404
rect 9875 38323 9881 38338
rect 9987 38323 9993 38338
rect 9875 38256 9881 38271
rect 9987 38256 9993 38271
rect 9875 37380 9881 38204
rect 9987 37380 9993 38204
rect 9875 36720 9993 37380
rect 9927 36668 9941 36720
rect 9875 36654 9993 36668
rect 9927 36602 9941 36654
rect 9875 36588 9993 36602
rect 9927 36536 9941 36588
rect 9875 36534 9881 36536
rect 9915 36534 9953 36536
rect 9987 36534 9993 36536
rect 9875 36522 9993 36534
rect 9927 36470 9941 36522
rect 9875 36461 9881 36470
rect 9915 36461 9953 36470
rect 9987 36461 9993 36470
rect 9875 36456 9993 36461
rect 9927 36422 9941 36456
rect 9875 36390 9881 36404
rect 9987 36390 9993 36404
rect 9875 36323 9881 36338
rect 9987 36323 9993 36338
rect 9875 36256 9881 36271
rect 9987 36256 9993 36271
rect 9875 35380 9881 36204
rect 9987 35380 9993 36204
rect 9875 35368 9993 35380
rect 10152 38714 10270 38726
rect 10152 38680 10158 38714
rect 10192 38680 10230 38714
rect 10264 38680 10270 38714
rect 10152 38641 10270 38680
rect 10152 38607 10158 38641
rect 10192 38607 10230 38641
rect 10264 38607 10270 38641
rect 10152 38568 10270 38607
rect 10152 38534 10158 38568
rect 10192 38534 10230 38568
rect 10264 38534 10270 38568
rect 10152 38495 10270 38534
rect 10152 38461 10158 38495
rect 10192 38461 10230 38495
rect 10264 38461 10270 38495
rect 10152 38422 10270 38461
rect 10152 37892 10158 38422
rect 10264 37892 10270 38422
rect 10152 37825 10158 37840
rect 10264 37825 10270 37840
rect 10152 37758 10158 37773
rect 10264 37758 10270 37773
rect 10152 37691 10158 37706
rect 10264 37691 10270 37706
rect 10152 37624 10158 37639
rect 10264 37624 10270 37639
rect 10152 37557 10158 37572
rect 10264 37557 10270 37572
rect 10152 37490 10158 37505
rect 10264 37490 10270 37505
rect 10152 37423 10158 37438
rect 10264 37423 10270 37438
rect 10204 37371 10218 37380
rect 10152 37356 10270 37371
rect 10204 37304 10218 37356
rect 10152 37289 10270 37304
rect 10204 37237 10218 37289
rect 10152 37222 10270 37237
rect 10204 37170 10218 37222
rect 10152 37155 10270 37170
rect 10204 37103 10218 37155
rect 10152 37088 10270 37103
rect 10204 37036 10218 37088
rect 10152 36714 10270 37036
rect 10152 36680 10158 36714
rect 10192 36680 10230 36714
rect 10264 36680 10270 36714
rect 10152 36641 10270 36680
rect 10152 36607 10158 36641
rect 10192 36607 10230 36641
rect 10264 36607 10270 36641
rect 10152 36568 10270 36607
rect 10152 36534 10158 36568
rect 10192 36534 10230 36568
rect 10264 36534 10270 36568
rect 10152 36495 10270 36534
rect 10152 36461 10158 36495
rect 10192 36461 10230 36495
rect 10264 36461 10270 36495
rect 10152 36422 10270 36461
rect 10152 35892 10158 36422
rect 10264 35892 10270 36422
rect 10152 35826 10158 35840
rect 10264 35826 10270 35840
rect 10152 35760 10158 35774
rect 10264 35760 10270 35774
rect 10152 35694 10158 35708
rect 10264 35694 10270 35708
rect 10152 35627 10158 35642
rect 10264 35627 10270 35642
rect 10152 35560 10158 35575
rect 10264 35560 10270 35575
rect 10152 35493 10158 35508
rect 10264 35493 10270 35508
rect 10152 35426 10158 35441
rect 10264 35426 10270 35441
rect 10204 35374 10218 35380
tri 9716 35280 9760 35324 sw
tri 10108 35280 10152 35324 se
rect 10152 35280 10270 35374
rect 10429 38720 10547 38726
rect 10481 38668 10495 38720
rect 10429 38654 10547 38668
rect 10481 38602 10495 38654
rect 10429 38588 10547 38602
rect 10481 38536 10495 38588
rect 10429 38534 10435 38536
rect 10469 38534 10507 38536
rect 10541 38534 10547 38536
rect 10429 38522 10547 38534
rect 10481 38470 10495 38522
rect 10429 38461 10435 38470
rect 10469 38461 10507 38470
rect 10541 38461 10547 38470
rect 10429 38456 10547 38461
rect 10481 38422 10495 38456
rect 10429 38390 10435 38404
rect 10541 38390 10547 38404
rect 10429 38323 10435 38338
rect 10541 38323 10547 38338
rect 10429 38256 10435 38271
rect 10541 38256 10547 38271
rect 10429 37380 10435 38204
rect 10541 37380 10547 38204
rect 10429 36720 10547 37380
rect 10481 36668 10495 36720
rect 10429 36654 10547 36668
rect 10481 36602 10495 36654
rect 10429 36588 10547 36602
rect 10481 36536 10495 36588
rect 10429 36534 10435 36536
rect 10469 36534 10507 36536
rect 10541 36534 10547 36536
rect 10429 36522 10547 36534
rect 10481 36470 10495 36522
rect 10429 36461 10435 36470
rect 10469 36461 10507 36470
rect 10541 36461 10547 36470
rect 10429 36456 10547 36461
rect 10481 36422 10495 36456
rect 10429 36390 10435 36404
rect 10541 36390 10547 36404
rect 10429 36323 10435 36338
rect 10541 36323 10547 36338
rect 10429 36256 10435 36271
rect 10541 36256 10547 36271
rect 10429 35380 10435 36204
rect 10541 35380 10547 36204
rect 10429 35368 10547 35380
rect 10706 38714 10824 38726
rect 10706 38680 10712 38714
rect 10746 38680 10784 38714
rect 10818 38680 10824 38714
rect 10706 38641 10824 38680
rect 10706 38607 10712 38641
rect 10746 38607 10784 38641
rect 10818 38607 10824 38641
rect 10706 38568 10824 38607
rect 10706 38534 10712 38568
rect 10746 38534 10784 38568
rect 10818 38534 10824 38568
rect 10706 38495 10824 38534
rect 10706 38461 10712 38495
rect 10746 38461 10784 38495
rect 10818 38461 10824 38495
rect 10706 38422 10824 38461
rect 10706 37892 10712 38422
rect 10818 37892 10824 38422
rect 10706 37825 10712 37840
rect 10818 37825 10824 37840
rect 10706 37758 10712 37773
rect 10818 37758 10824 37773
rect 10706 37691 10712 37706
rect 10818 37691 10824 37706
rect 10706 37624 10712 37639
rect 10818 37624 10824 37639
rect 10706 37557 10712 37572
rect 10818 37557 10824 37572
rect 10706 37490 10712 37505
rect 10818 37490 10824 37505
rect 10706 37423 10712 37438
rect 10818 37423 10824 37438
rect 10758 37371 10772 37380
rect 10706 37356 10824 37371
rect 10758 37304 10772 37356
rect 10706 37289 10824 37304
rect 10758 37237 10772 37289
rect 10706 37222 10824 37237
rect 10758 37170 10772 37222
rect 10706 37155 10824 37170
rect 10758 37103 10772 37155
rect 10706 37088 10824 37103
rect 10758 37036 10772 37088
rect 10706 36714 10824 37036
rect 10706 36680 10712 36714
rect 10746 36680 10784 36714
rect 10818 36680 10824 36714
rect 10706 36641 10824 36680
rect 10706 36607 10712 36641
rect 10746 36607 10784 36641
rect 10818 36607 10824 36641
rect 10706 36568 10824 36607
rect 10706 36534 10712 36568
rect 10746 36534 10784 36568
rect 10818 36534 10824 36568
rect 10706 36495 10824 36534
rect 10706 36461 10712 36495
rect 10746 36461 10784 36495
rect 10818 36461 10824 36495
rect 10706 36422 10824 36461
rect 10706 35892 10712 36422
rect 10818 35892 10824 36422
rect 10706 35826 10712 35840
rect 10818 35826 10824 35840
rect 10706 35760 10712 35774
rect 10818 35760 10824 35774
rect 10706 35694 10712 35708
rect 10818 35694 10824 35708
rect 10706 35627 10712 35642
rect 10818 35627 10824 35642
rect 10706 35560 10712 35575
rect 10818 35560 10824 35575
rect 10706 35493 10712 35508
rect 10818 35493 10824 35508
rect 10706 35426 10712 35441
rect 10818 35426 10824 35441
rect 10758 35374 10772 35380
tri 10270 35280 10314 35324 sw
tri 10662 35280 10706 35324 se
rect 10706 35280 10824 35374
rect 10983 38720 11101 38726
rect 11035 38668 11049 38720
rect 10983 38654 11101 38668
rect 11035 38602 11049 38654
rect 10983 38588 11101 38602
rect 11035 38536 11049 38588
rect 10983 38534 10989 38536
rect 11023 38534 11061 38536
rect 11095 38534 11101 38536
rect 10983 38522 11101 38534
rect 11035 38470 11049 38522
rect 10983 38461 10989 38470
rect 11023 38461 11061 38470
rect 11095 38461 11101 38470
rect 10983 38456 11101 38461
rect 11035 38422 11049 38456
rect 10983 38390 10989 38404
rect 11095 38390 11101 38404
rect 10983 38323 10989 38338
rect 11095 38323 11101 38338
rect 10983 38256 10989 38271
rect 11095 38256 11101 38271
rect 10983 37380 10989 38204
rect 11095 37380 11101 38204
rect 10983 36720 11101 37380
rect 11035 36668 11049 36720
rect 10983 36654 11101 36668
rect 11035 36602 11049 36654
rect 10983 36588 11101 36602
rect 11035 36536 11049 36588
rect 10983 36534 10989 36536
rect 11023 36534 11061 36536
rect 11095 36534 11101 36536
rect 10983 36522 11101 36534
rect 11035 36470 11049 36522
rect 10983 36461 10989 36470
rect 11023 36461 11061 36470
rect 11095 36461 11101 36470
rect 10983 36456 11101 36461
rect 11035 36422 11049 36456
rect 10983 36390 10989 36404
rect 11095 36390 11101 36404
rect 10983 36323 10989 36338
rect 11095 36323 11101 36338
rect 10983 36256 10989 36271
rect 11095 36256 11101 36271
rect 10983 35380 10989 36204
rect 11095 35380 11101 36204
rect 10983 35368 11101 35380
rect 11260 38714 11378 38726
rect 11260 38680 11266 38714
rect 11300 38680 11338 38714
rect 11372 38680 11378 38714
rect 11260 38641 11378 38680
rect 11260 38607 11266 38641
rect 11300 38607 11338 38641
rect 11372 38607 11378 38641
rect 11260 38568 11378 38607
rect 11260 38534 11266 38568
rect 11300 38534 11338 38568
rect 11372 38534 11378 38568
rect 11260 38495 11378 38534
rect 11260 38461 11266 38495
rect 11300 38461 11338 38495
rect 11372 38461 11378 38495
rect 11260 38422 11378 38461
rect 11260 37892 11266 38422
rect 11372 37892 11378 38422
rect 11260 37825 11266 37840
rect 11372 37825 11378 37840
rect 11260 37758 11266 37773
rect 11372 37758 11378 37773
rect 11260 37691 11266 37706
rect 11372 37691 11378 37706
rect 11260 37624 11266 37639
rect 11372 37624 11378 37639
rect 11260 37557 11266 37572
rect 11372 37557 11378 37572
rect 11260 37490 11266 37505
rect 11372 37490 11378 37505
rect 11260 37423 11266 37438
rect 11372 37423 11378 37438
rect 11312 37371 11326 37380
rect 11260 37356 11378 37371
rect 11312 37304 11326 37356
rect 11260 37289 11378 37304
rect 11312 37237 11326 37289
rect 11260 37222 11378 37237
rect 11312 37170 11326 37222
rect 11260 37155 11378 37170
rect 11312 37103 11326 37155
rect 11260 37088 11378 37103
rect 11312 37036 11326 37088
rect 11260 36714 11378 37036
rect 11260 36680 11266 36714
rect 11300 36680 11338 36714
rect 11372 36680 11378 36714
rect 11260 36641 11378 36680
rect 11260 36607 11266 36641
rect 11300 36607 11338 36641
rect 11372 36607 11378 36641
rect 11260 36568 11378 36607
rect 11260 36534 11266 36568
rect 11300 36534 11338 36568
rect 11372 36534 11378 36568
rect 11260 36495 11378 36534
rect 11260 36461 11266 36495
rect 11300 36461 11338 36495
rect 11372 36461 11378 36495
rect 11260 36422 11378 36461
rect 11260 35892 11266 36422
rect 11372 35892 11378 36422
rect 11260 35826 11266 35840
rect 11372 35826 11378 35840
rect 11260 35760 11266 35774
rect 11372 35760 11378 35774
rect 11260 35694 11266 35708
rect 11372 35694 11378 35708
rect 11260 35627 11266 35642
rect 11372 35627 11378 35642
rect 11260 35560 11266 35575
rect 11372 35560 11378 35575
rect 11260 35493 11266 35508
rect 11372 35493 11378 35508
rect 11260 35426 11266 35441
rect 11372 35426 11378 35441
rect 11312 35374 11326 35380
tri 10824 35280 10868 35324 sw
tri 11216 35280 11260 35324 se
rect 11260 35280 11378 35374
rect 11537 38720 11655 38726
rect 11589 38668 11603 38720
rect 11537 38654 11655 38668
rect 11589 38602 11603 38654
rect 11537 38588 11655 38602
rect 11589 38536 11603 38588
rect 11537 38534 11543 38536
rect 11577 38534 11615 38536
rect 11649 38534 11655 38536
rect 11537 38522 11655 38534
rect 11589 38470 11603 38522
rect 11537 38461 11543 38470
rect 11577 38461 11615 38470
rect 11649 38461 11655 38470
rect 11537 38456 11655 38461
rect 11589 38422 11603 38456
rect 11537 38390 11543 38404
rect 11649 38390 11655 38404
rect 11537 38323 11543 38338
rect 11649 38323 11655 38338
rect 11537 38256 11543 38271
rect 11649 38256 11655 38271
rect 11537 37380 11543 38204
rect 11649 37380 11655 38204
rect 11537 36720 11655 37380
rect 11589 36668 11603 36720
rect 11537 36654 11655 36668
rect 11589 36602 11603 36654
rect 11537 36588 11655 36602
rect 11589 36536 11603 36588
rect 11537 36534 11543 36536
rect 11577 36534 11615 36536
rect 11649 36534 11655 36536
rect 11537 36522 11655 36534
rect 11589 36470 11603 36522
rect 11537 36461 11543 36470
rect 11577 36461 11615 36470
rect 11649 36461 11655 36470
rect 11537 36456 11655 36461
rect 11589 36422 11603 36456
rect 11537 36390 11543 36404
rect 11649 36390 11655 36404
rect 11537 36323 11543 36338
rect 11649 36323 11655 36338
rect 11537 36256 11543 36271
rect 11649 36256 11655 36271
rect 11537 35380 11543 36204
rect 11649 35380 11655 36204
rect 11537 35368 11655 35380
rect 11814 38714 11932 38726
rect 11814 38680 11820 38714
rect 11854 38680 11892 38714
rect 11926 38680 11932 38714
rect 11814 38641 11932 38680
rect 11814 38607 11820 38641
rect 11854 38607 11892 38641
rect 11926 38607 11932 38641
rect 11814 38568 11932 38607
rect 11814 38534 11820 38568
rect 11854 38534 11892 38568
rect 11926 38534 11932 38568
rect 11814 38495 11932 38534
rect 11814 38461 11820 38495
rect 11854 38461 11892 38495
rect 11926 38461 11932 38495
rect 11814 38422 11932 38461
rect 11814 37892 11820 38422
rect 11926 37892 11932 38422
rect 11814 37825 11820 37840
rect 11926 37825 11932 37840
rect 11814 37758 11820 37773
rect 11926 37758 11932 37773
rect 11814 37691 11820 37706
rect 11926 37691 11932 37706
rect 11814 37624 11820 37639
rect 11926 37624 11932 37639
rect 11814 37557 11820 37572
rect 11926 37557 11932 37572
rect 11814 37490 11820 37505
rect 11926 37490 11932 37505
rect 11814 37423 11820 37438
rect 11926 37423 11932 37438
rect 11866 37371 11880 37380
rect 11814 37356 11932 37371
rect 11866 37304 11880 37356
rect 11814 37289 11932 37304
rect 11866 37237 11880 37289
rect 11814 37222 11932 37237
rect 11866 37170 11880 37222
rect 11814 37155 11932 37170
rect 11866 37103 11880 37155
rect 11814 37088 11932 37103
rect 11866 37036 11880 37088
rect 11814 36714 11932 37036
rect 11814 36680 11820 36714
rect 11854 36680 11892 36714
rect 11926 36680 11932 36714
rect 11814 36641 11932 36680
rect 11814 36607 11820 36641
rect 11854 36607 11892 36641
rect 11926 36607 11932 36641
rect 11814 36568 11932 36607
rect 11814 36534 11820 36568
rect 11854 36534 11892 36568
rect 11926 36534 11932 36568
rect 11814 36495 11932 36534
rect 11814 36461 11820 36495
rect 11854 36461 11892 36495
rect 11926 36461 11932 36495
rect 11814 36422 11932 36461
rect 11814 35892 11820 36422
rect 11926 35892 11932 36422
rect 11814 35826 11820 35840
rect 11926 35826 11932 35840
rect 11814 35760 11820 35774
rect 11926 35760 11932 35774
rect 11814 35694 11820 35708
rect 11926 35694 11932 35708
rect 11814 35627 11820 35642
rect 11926 35627 11932 35642
rect 11814 35560 11820 35575
rect 11926 35560 11932 35575
rect 11814 35493 11820 35508
rect 11926 35493 11932 35508
rect 11814 35426 11820 35441
rect 11926 35426 11932 35441
rect 11866 35374 11880 35380
tri 11378 35280 11422 35324 sw
tri 11770 35280 11814 35324 se
rect 11814 35280 11932 35374
rect 12091 38720 12209 38726
rect 12143 38668 12157 38720
rect 12091 38654 12209 38668
rect 12143 38602 12157 38654
rect 12091 38588 12209 38602
rect 12143 38536 12157 38588
rect 12091 38534 12097 38536
rect 12131 38534 12169 38536
rect 12203 38534 12209 38536
rect 12091 38522 12209 38534
rect 12143 38470 12157 38522
rect 12091 38461 12097 38470
rect 12131 38461 12169 38470
rect 12203 38461 12209 38470
rect 12091 38456 12209 38461
rect 12143 38422 12157 38456
rect 12091 38390 12097 38404
rect 12203 38390 12209 38404
rect 12091 38323 12097 38338
rect 12203 38323 12209 38338
rect 12091 38256 12097 38271
rect 12203 38256 12209 38271
rect 12091 37380 12097 38204
rect 12203 37380 12209 38204
rect 12091 36720 12209 37380
rect 12143 36668 12157 36720
rect 12091 36654 12209 36668
rect 12143 36602 12157 36654
rect 12091 36588 12209 36602
rect 12143 36536 12157 36588
rect 12091 36534 12097 36536
rect 12131 36534 12169 36536
rect 12203 36534 12209 36536
rect 12091 36522 12209 36534
rect 12143 36470 12157 36522
rect 12091 36461 12097 36470
rect 12131 36461 12169 36470
rect 12203 36461 12209 36470
rect 12091 36456 12209 36461
rect 12143 36422 12157 36456
rect 12091 36390 12097 36404
rect 12203 36390 12209 36404
rect 12091 36323 12097 36338
rect 12203 36323 12209 36338
rect 12091 36256 12097 36271
rect 12203 36256 12209 36271
rect 12091 35380 12097 36204
rect 12203 35380 12209 36204
rect 12091 35368 12209 35380
rect 12368 38714 12486 38726
rect 12368 38680 12374 38714
rect 12408 38680 12446 38714
rect 12480 38680 12486 38714
rect 12368 38641 12486 38680
rect 12368 38607 12374 38641
rect 12408 38607 12446 38641
rect 12480 38607 12486 38641
rect 12368 38568 12486 38607
rect 12368 38534 12374 38568
rect 12408 38534 12446 38568
rect 12480 38534 12486 38568
rect 12368 38495 12486 38534
rect 12368 38461 12374 38495
rect 12408 38461 12446 38495
rect 12480 38461 12486 38495
rect 12368 38422 12486 38461
rect 12368 37892 12374 38422
rect 12480 37892 12486 38422
rect 12368 37825 12374 37840
rect 12480 37825 12486 37840
rect 12368 37758 12374 37773
rect 12480 37758 12486 37773
rect 12368 37691 12374 37706
rect 12480 37691 12486 37706
rect 12368 37624 12374 37639
rect 12480 37624 12486 37639
rect 12368 37557 12374 37572
rect 12480 37557 12486 37572
rect 12368 37490 12374 37505
rect 12480 37490 12486 37505
rect 12368 37423 12374 37438
rect 12480 37423 12486 37438
rect 12420 37371 12434 37380
rect 12368 37356 12486 37371
rect 12420 37304 12434 37356
rect 12368 37289 12486 37304
rect 12420 37237 12434 37289
rect 12368 37222 12486 37237
rect 12420 37170 12434 37222
rect 12368 37155 12486 37170
rect 12420 37103 12434 37155
rect 12368 37088 12486 37103
rect 12420 37036 12434 37088
rect 12368 36714 12486 37036
rect 12368 36680 12374 36714
rect 12408 36680 12446 36714
rect 12480 36680 12486 36714
rect 12368 36641 12486 36680
rect 12368 36607 12374 36641
rect 12408 36607 12446 36641
rect 12480 36607 12486 36641
rect 12368 36568 12486 36607
rect 12368 36534 12374 36568
rect 12408 36534 12446 36568
rect 12480 36534 12486 36568
rect 12368 36495 12486 36534
rect 12368 36461 12374 36495
rect 12408 36461 12446 36495
rect 12480 36461 12486 36495
rect 12368 36422 12486 36461
rect 12368 35892 12374 36422
rect 12480 35892 12486 36422
rect 12368 35826 12374 35840
rect 12480 35826 12486 35840
rect 12368 35760 12374 35774
rect 12480 35760 12486 35774
rect 12368 35694 12374 35708
rect 12480 35694 12486 35708
rect 12368 35627 12374 35642
rect 12480 35627 12486 35642
rect 12368 35560 12374 35575
rect 12480 35560 12486 35575
rect 12368 35493 12374 35508
rect 12480 35493 12486 35508
rect 12368 35426 12374 35441
rect 12480 35426 12486 35441
rect 12420 35374 12434 35380
tri 11932 35280 11976 35324 sw
tri 12324 35280 12368 35324 se
rect 12368 35280 12486 35374
rect 12645 38720 12763 38726
rect 12697 38668 12711 38720
rect 12645 38654 12763 38668
rect 12697 38602 12711 38654
rect 12645 38588 12763 38602
rect 12697 38536 12711 38588
rect 12645 38534 12651 38536
rect 12685 38534 12723 38536
rect 12757 38534 12763 38536
rect 12645 38522 12763 38534
rect 12697 38470 12711 38522
rect 12645 38461 12651 38470
rect 12685 38461 12723 38470
rect 12757 38461 12763 38470
rect 12645 38456 12763 38461
rect 12697 38422 12711 38456
rect 12645 38390 12651 38404
rect 12757 38390 12763 38404
rect 12645 38323 12651 38338
rect 12757 38323 12763 38338
rect 12645 38256 12651 38271
rect 12757 38256 12763 38271
rect 12645 37380 12651 38204
rect 12757 37380 12763 38204
rect 12645 36720 12763 37380
rect 12697 36668 12711 36720
rect 12645 36654 12763 36668
rect 12697 36602 12711 36654
rect 12645 36588 12763 36602
rect 12697 36536 12711 36588
rect 12645 36534 12651 36536
rect 12685 36534 12723 36536
rect 12757 36534 12763 36536
rect 12645 36522 12763 36534
rect 12697 36470 12711 36522
rect 12645 36461 12651 36470
rect 12685 36461 12723 36470
rect 12757 36461 12763 36470
rect 12645 36456 12763 36461
rect 12697 36422 12711 36456
rect 12645 36390 12651 36404
rect 12757 36390 12763 36404
rect 12645 36323 12651 36338
rect 12757 36323 12763 36338
rect 12645 36256 12651 36271
rect 12757 36256 12763 36271
rect 12645 35380 12651 36204
rect 12757 35380 12763 36204
rect 12645 35368 12763 35380
rect 12922 38714 13040 38726
rect 12922 38680 12928 38714
rect 12962 38680 13000 38714
rect 13034 38680 13040 38714
rect 12922 38641 13040 38680
rect 12922 38607 12928 38641
rect 12962 38607 13000 38641
rect 13034 38607 13040 38641
rect 12922 38568 13040 38607
rect 12922 38534 12928 38568
rect 12962 38534 13000 38568
rect 13034 38534 13040 38568
rect 12922 38495 13040 38534
rect 12922 38461 12928 38495
rect 12962 38461 13000 38495
rect 13034 38461 13040 38495
rect 12922 38422 13040 38461
rect 12922 37892 12928 38422
rect 13034 37892 13040 38422
rect 12922 37825 12928 37840
rect 13034 37825 13040 37840
rect 12922 37758 12928 37773
rect 13034 37758 13040 37773
rect 12922 37691 12928 37706
rect 13034 37691 13040 37706
rect 12922 37624 12928 37639
rect 13034 37624 13040 37639
rect 12922 37557 12928 37572
rect 13034 37557 13040 37572
rect 12922 37490 12928 37505
rect 13034 37490 13040 37505
rect 12922 37423 12928 37438
rect 13034 37423 13040 37438
rect 12974 37371 12988 37380
rect 12922 37356 13040 37371
rect 12974 37304 12988 37356
rect 12922 37289 13040 37304
rect 12974 37237 12988 37289
rect 12922 37222 13040 37237
rect 12974 37170 12988 37222
rect 12922 37155 13040 37170
rect 12974 37103 12988 37155
rect 12922 37088 13040 37103
rect 12974 37036 12988 37088
rect 12922 36714 13040 37036
rect 12922 36680 12928 36714
rect 12962 36680 13000 36714
rect 13034 36680 13040 36714
rect 12922 36641 13040 36680
rect 12922 36607 12928 36641
rect 12962 36607 13000 36641
rect 13034 36607 13040 36641
rect 12922 36568 13040 36607
rect 12922 36534 12928 36568
rect 12962 36534 13000 36568
rect 13034 36534 13040 36568
rect 12922 36495 13040 36534
rect 12922 36461 12928 36495
rect 12962 36461 13000 36495
rect 13034 36461 13040 36495
rect 12922 36422 13040 36461
rect 12922 35892 12928 36422
rect 13034 35892 13040 36422
rect 12922 35826 12928 35840
rect 13034 35826 13040 35840
rect 12922 35760 12928 35774
rect 13034 35760 13040 35774
rect 12922 35694 12928 35708
rect 13034 35694 13040 35708
rect 12922 35627 12928 35642
rect 13034 35627 13040 35642
rect 12922 35560 12928 35575
rect 13034 35560 13040 35575
rect 12922 35493 12928 35508
rect 13034 35493 13040 35508
rect 12922 35426 12928 35441
rect 13034 35426 13040 35441
rect 12974 35374 12988 35380
tri 12486 35280 12530 35324 sw
tri 12878 35280 12922 35324 se
rect 12922 35280 13040 35374
rect 3504 34891 13040 35280
rect 13199 38720 13521 38726
rect 13199 38668 13200 38720
rect 13252 38668 13270 38720
rect 13322 38668 13340 38720
rect 13392 38668 13410 38720
rect 13462 38668 13480 38720
rect 13199 38654 13521 38668
rect 13199 38602 13200 38654
rect 13252 38602 13270 38654
rect 13322 38602 13340 38654
rect 13392 38602 13410 38654
rect 13462 38602 13480 38654
rect 13199 38588 13521 38602
rect 13199 38536 13200 38588
rect 13252 38536 13270 38588
rect 13322 38536 13340 38588
rect 13392 38536 13410 38588
rect 13462 38536 13480 38588
rect 13199 38534 13205 38536
rect 13239 38534 13277 38536
rect 13311 38534 13521 38536
rect 13199 38522 13521 38534
rect 13199 38470 13200 38522
rect 13252 38470 13270 38522
rect 13322 38470 13340 38522
rect 13392 38470 13410 38522
rect 13462 38470 13480 38522
rect 13199 38461 13205 38470
rect 13239 38461 13277 38470
rect 13311 38461 13521 38470
rect 13199 38456 13521 38461
rect 13199 38404 13200 38456
rect 13252 38422 13270 38456
rect 13322 38404 13340 38456
rect 13392 38404 13410 38456
rect 13462 38404 13480 38456
rect 13199 38390 13205 38404
rect 13311 38390 13521 38404
rect 13199 38338 13200 38390
rect 13322 38338 13340 38390
rect 13392 38338 13410 38390
rect 13462 38338 13480 38390
rect 13199 38323 13205 38338
rect 13311 38323 13521 38338
rect 13199 38271 13200 38323
rect 13322 38271 13340 38323
rect 13392 38271 13410 38323
rect 13462 38271 13480 38323
rect 13199 38256 13205 38271
rect 13311 38256 13521 38271
rect 13199 38204 13200 38256
rect 13322 38204 13340 38256
rect 13392 38204 13410 38256
rect 13462 38204 13480 38256
rect 13199 37380 13205 38204
rect 13311 37380 13521 38204
rect 13199 36720 13521 37380
rect 13199 36668 13200 36720
rect 13252 36668 13270 36720
rect 13322 36668 13340 36720
rect 13392 36668 13410 36720
rect 13462 36668 13480 36720
rect 13199 36654 13521 36668
rect 13199 36602 13200 36654
rect 13252 36602 13270 36654
rect 13322 36602 13340 36654
rect 13392 36602 13410 36654
rect 13462 36602 13480 36654
rect 13199 36588 13521 36602
rect 13199 36536 13200 36588
rect 13252 36536 13270 36588
rect 13322 36536 13340 36588
rect 13392 36536 13410 36588
rect 13462 36536 13480 36588
rect 13199 36534 13205 36536
rect 13239 36534 13277 36536
rect 13311 36534 13521 36536
rect 13199 36522 13521 36534
rect 13199 36470 13200 36522
rect 13252 36470 13270 36522
rect 13322 36470 13340 36522
rect 13392 36470 13410 36522
rect 13462 36470 13480 36522
rect 13199 36461 13205 36470
rect 13239 36461 13277 36470
rect 13311 36461 13521 36470
rect 13199 36456 13521 36461
rect 13199 36404 13200 36456
rect 13252 36422 13270 36456
rect 13322 36404 13340 36456
rect 13392 36404 13410 36456
rect 13462 36404 13480 36456
rect 13199 36390 13205 36404
rect 13311 36390 13521 36404
rect 13199 36338 13200 36390
rect 13322 36338 13340 36390
rect 13392 36338 13410 36390
rect 13462 36338 13480 36390
rect 13199 36323 13205 36338
rect 13311 36323 13521 36338
rect 13199 36271 13200 36323
rect 13322 36271 13340 36323
rect 13392 36271 13410 36323
rect 13462 36271 13480 36323
rect 13199 36256 13205 36271
rect 13311 36256 13521 36271
rect 13199 36204 13200 36256
rect 13322 36204 13340 36256
rect 13392 36204 13410 36256
rect 13462 36204 13480 36256
rect 13199 35380 13205 36204
rect 13311 35380 13521 36204
tri 3504 34810 3585 34891 ne
rect 2667 33288 2674 33322
rect 2708 33288 2750 33322
rect 2784 33288 2826 33322
rect 2860 33288 2867 33322
rect 2667 33245 2867 33288
rect 2667 33211 2674 33245
rect 2708 33211 2750 33245
rect 2784 33211 2826 33245
rect 2860 33211 2867 33245
rect 2667 33168 2867 33211
rect 2667 33134 2674 33168
rect 2708 33134 2750 33168
rect 2784 33134 2826 33168
rect 2860 33134 2867 33168
rect 2667 33090 2867 33134
rect 2667 33056 2674 33090
rect 2708 33056 2750 33090
rect 2784 33056 2826 33090
rect 2860 33056 2867 33090
rect 2667 33012 2867 33056
rect 2667 32978 2674 33012
rect 2708 32978 2750 33012
rect 2784 32978 2826 33012
rect 2860 32978 2867 33012
rect 2667 32934 2867 32978
rect 2667 32900 2674 32934
rect 2708 32900 2750 32934
rect 2784 32900 2826 32934
rect 2860 32900 2867 32934
rect 2667 32856 2867 32900
rect 2667 32822 2674 32856
rect 2708 32822 2750 32856
rect 2784 32822 2826 32856
rect 2860 32822 2867 32856
rect 2667 31323 2867 32822
rect 2667 31289 2674 31323
rect 2708 31289 2750 31323
rect 2784 31289 2826 31323
rect 2860 31289 2867 31323
rect 2667 31246 2867 31289
rect 2667 31212 2674 31246
rect 2708 31212 2750 31246
rect 2784 31212 2826 31246
rect 2860 31212 2867 31246
rect 2667 31169 2867 31212
rect 2667 31135 2674 31169
rect 2708 31135 2750 31169
rect 2784 31135 2826 31169
rect 2860 31135 2867 31169
rect 2667 31091 2867 31135
rect 2667 31057 2674 31091
rect 2708 31057 2750 31091
rect 2784 31057 2826 31091
rect 2860 31057 2867 31091
rect 2667 31013 2867 31057
rect 2667 30979 2674 31013
rect 2708 30979 2750 31013
rect 2784 30979 2826 31013
rect 2860 30979 2867 31013
rect 2667 30935 2867 30979
rect 2667 30901 2674 30935
rect 2708 30901 2750 30935
rect 2784 30901 2826 30935
rect 2860 30901 2867 30935
rect 2667 30857 2867 30901
rect 2667 30823 2674 30857
rect 2708 30823 2750 30857
rect 2784 30823 2826 30857
rect 2860 30823 2867 30857
rect 2667 29320 2867 30823
rect 3167 34720 3285 34726
rect 3219 34668 3233 34720
rect 3167 34654 3285 34668
rect 3219 34602 3233 34654
rect 3167 34588 3285 34602
rect 3219 34536 3233 34588
rect 3167 34534 3173 34536
rect 3207 34534 3245 34536
rect 3279 34534 3285 34536
rect 3167 34522 3285 34534
rect 3219 34470 3233 34522
rect 3167 34461 3173 34470
rect 3207 34461 3245 34470
rect 3279 34461 3285 34470
rect 3167 34456 3285 34461
rect 3219 34422 3233 34456
rect 3167 34390 3173 34404
rect 3279 34390 3285 34404
rect 3167 34323 3173 34338
rect 3279 34323 3285 34338
rect 3167 34256 3173 34271
rect 3279 34256 3285 34271
rect 3167 33380 3173 34204
rect 3279 33380 3285 34204
rect 3167 32720 3285 33380
rect 3219 32668 3233 32720
rect 3167 32654 3285 32668
rect 3219 32602 3233 32654
rect 3167 32588 3285 32602
rect 3219 32536 3233 32588
rect 3167 32534 3173 32536
rect 3207 32534 3245 32536
rect 3279 32534 3285 32536
rect 3167 32522 3285 32534
rect 3219 32470 3233 32522
rect 3167 32461 3173 32470
rect 3207 32461 3245 32470
rect 3279 32461 3285 32470
rect 3167 32456 3285 32461
rect 3219 32422 3233 32456
rect 3167 32390 3173 32404
rect 3279 32390 3285 32404
rect 3167 32323 3173 32338
rect 3279 32323 3285 32338
rect 3167 32256 3173 32271
rect 3279 32256 3285 32271
rect 3167 31380 3173 32204
rect 3279 31380 3285 32204
rect 3167 30720 3285 31380
rect 3219 30668 3233 30720
rect 3167 30654 3285 30668
rect 3219 30602 3233 30654
rect 3167 30588 3285 30602
rect 3219 30536 3233 30588
rect 3167 30534 3173 30536
rect 3207 30534 3245 30536
rect 3279 30534 3285 30536
rect 3167 30522 3285 30534
rect 3219 30470 3233 30522
rect 3167 30461 3173 30470
rect 3207 30461 3245 30470
rect 3279 30461 3285 30470
rect 3167 30456 3285 30461
rect 3219 30422 3233 30456
rect 3167 30390 3173 30404
rect 3279 30390 3285 30404
rect 3167 30323 3173 30338
rect 3279 30323 3285 30338
rect 3167 30256 3173 30271
rect 3279 30256 3285 30271
rect 3167 29380 3173 30204
rect 3279 29380 3285 30204
rect 3167 29368 3285 29380
rect 3585 34714 3703 34891
tri 3703 34821 3773 34891 nw
tri 4351 34821 4421 34891 ne
rect 3585 34680 3591 34714
rect 3625 34680 3663 34714
rect 3697 34680 3703 34714
rect 3585 34641 3703 34680
rect 3585 34607 3591 34641
rect 3625 34607 3663 34641
rect 3697 34607 3703 34641
rect 3585 34568 3703 34607
rect 3585 34534 3591 34568
rect 3625 34534 3663 34568
rect 3697 34534 3703 34568
rect 3585 34495 3703 34534
rect 3585 34461 3591 34495
rect 3625 34461 3663 34495
rect 3697 34461 3703 34495
rect 3585 34422 3703 34461
rect 3585 33892 3591 34422
rect 3697 33892 3703 34422
rect 3585 33826 3591 33840
rect 3697 33826 3703 33840
rect 3585 33760 3591 33774
rect 3697 33760 3703 33774
rect 3585 33694 3591 33708
rect 3697 33694 3703 33708
rect 3585 33627 3591 33642
rect 3697 33627 3703 33642
rect 3585 33560 3591 33575
rect 3697 33560 3703 33575
rect 3585 33493 3591 33508
rect 3697 33493 3703 33508
rect 3585 33426 3591 33441
rect 3697 33426 3703 33441
rect 3637 33374 3651 33380
rect 3585 32714 3703 33374
rect 3585 32680 3591 32714
rect 3625 32680 3663 32714
rect 3697 32680 3703 32714
rect 3585 32641 3703 32680
rect 3585 32607 3591 32641
rect 3625 32607 3663 32641
rect 3697 32607 3703 32641
rect 3585 32568 3703 32607
rect 3585 32534 3591 32568
rect 3625 32534 3663 32568
rect 3697 32534 3703 32568
rect 3585 32495 3703 32534
rect 3585 32461 3591 32495
rect 3625 32461 3663 32495
rect 3697 32461 3703 32495
rect 3585 32422 3703 32461
rect 3585 31892 3591 32422
rect 3697 31892 3703 32422
rect 3585 31826 3591 31840
rect 3697 31826 3703 31840
rect 3585 31760 3591 31774
rect 3697 31760 3703 31774
rect 3585 31694 3591 31708
rect 3697 31694 3703 31708
rect 3585 31627 3591 31642
rect 3697 31627 3703 31642
rect 3585 31560 3591 31575
rect 3697 31560 3703 31575
rect 3585 31493 3591 31508
rect 3697 31493 3703 31508
rect 3585 31426 3591 31441
rect 3697 31426 3703 31441
rect 3637 31374 3651 31380
rect 3585 30714 3703 31374
rect 3585 30680 3591 30714
rect 3625 30680 3663 30714
rect 3697 30680 3703 30714
rect 3585 30641 3703 30680
rect 3585 30607 3591 30641
rect 3625 30607 3663 30641
rect 3697 30607 3703 30641
rect 3585 30568 3703 30607
rect 3585 30534 3591 30568
rect 3625 30534 3663 30568
rect 3697 30534 3703 30568
rect 3585 30495 3703 30534
rect 3585 30461 3591 30495
rect 3625 30461 3663 30495
rect 3697 30461 3703 30495
rect 3585 30422 3703 30461
rect 3585 29892 3591 30422
rect 3697 29892 3703 30422
rect 3585 29826 3591 29840
rect 3697 29826 3703 29840
rect 3585 29760 3591 29774
rect 3697 29760 3703 29774
rect 3585 29694 3591 29708
rect 3697 29694 3703 29708
rect 3585 29627 3591 29642
rect 3697 29627 3703 29642
rect 3585 29560 3591 29575
rect 3697 29560 3703 29575
rect 3585 29493 3591 29508
rect 3697 29493 3703 29508
rect 3585 29426 3591 29441
rect 3697 29426 3703 29441
rect 3637 29374 3651 29380
rect 3585 29368 3703 29374
rect 4003 34720 4121 34726
rect 4055 34668 4069 34720
rect 4003 34654 4121 34668
rect 4055 34602 4069 34654
rect 4003 34588 4121 34602
rect 4055 34536 4069 34588
rect 4003 34534 4009 34536
rect 4043 34534 4081 34536
rect 4115 34534 4121 34536
rect 4003 34522 4121 34534
rect 4055 34470 4069 34522
rect 4003 34461 4009 34470
rect 4043 34461 4081 34470
rect 4115 34461 4121 34470
rect 4003 34456 4121 34461
rect 4055 34422 4069 34456
rect 4003 34390 4009 34404
rect 4115 34390 4121 34404
rect 4003 34323 4009 34338
rect 4115 34323 4121 34338
rect 4003 34256 4009 34271
rect 4115 34256 4121 34271
rect 4003 33380 4009 34204
rect 4115 33380 4121 34204
rect 4003 32720 4121 33380
rect 4055 32668 4069 32720
rect 4003 32654 4121 32668
rect 4055 32602 4069 32654
rect 4003 32588 4121 32602
rect 4055 32536 4069 32588
rect 4003 32534 4009 32536
rect 4043 32534 4081 32536
rect 4115 32534 4121 32536
rect 4003 32522 4121 32534
rect 4055 32470 4069 32522
rect 4003 32461 4009 32470
rect 4043 32461 4081 32470
rect 4115 32461 4121 32470
rect 4003 32456 4121 32461
rect 4055 32422 4069 32456
rect 4003 32390 4009 32404
rect 4115 32390 4121 32404
rect 4003 32323 4009 32338
rect 4115 32323 4121 32338
rect 4003 32256 4009 32271
rect 4115 32256 4121 32271
rect 4003 31380 4009 32204
rect 4115 31380 4121 32204
rect 4003 30720 4121 31380
rect 4055 30668 4069 30720
rect 4003 30654 4121 30668
rect 4055 30602 4069 30654
rect 4003 30588 4121 30602
rect 4055 30536 4069 30588
rect 4003 30534 4009 30536
rect 4043 30534 4081 30536
rect 4115 30534 4121 30536
rect 4003 30522 4121 30534
rect 4055 30470 4069 30522
rect 4003 30461 4009 30470
rect 4043 30461 4081 30470
rect 4115 30461 4121 30470
rect 4003 30456 4121 30461
rect 4055 30422 4069 30456
rect 4003 30390 4009 30404
rect 4115 30390 4121 30404
rect 4003 30323 4009 30338
rect 4115 30323 4121 30338
rect 4003 30256 4009 30271
rect 4115 30256 4121 30271
rect 4003 29380 4009 30204
rect 4115 29380 4121 30204
rect 4003 29368 4121 29380
rect 4421 34714 4539 34891
tri 4539 34821 4609 34891 nw
tri 5187 34821 5257 34891 ne
rect 4421 34680 4427 34714
rect 4461 34680 4499 34714
rect 4533 34680 4539 34714
rect 4421 34641 4539 34680
rect 4421 34607 4427 34641
rect 4461 34607 4499 34641
rect 4533 34607 4539 34641
rect 4421 34568 4539 34607
rect 4421 34534 4427 34568
rect 4461 34534 4499 34568
rect 4533 34534 4539 34568
rect 4421 34495 4539 34534
rect 4421 34461 4427 34495
rect 4461 34461 4499 34495
rect 4533 34461 4539 34495
rect 4421 34422 4539 34461
rect 4421 33892 4427 34422
rect 4533 33892 4539 34422
rect 4421 33826 4427 33840
rect 4533 33826 4539 33840
rect 4421 33760 4427 33774
rect 4533 33760 4539 33774
rect 4421 33694 4427 33708
rect 4533 33694 4539 33708
rect 4421 33627 4427 33642
rect 4533 33627 4539 33642
rect 4421 33560 4427 33575
rect 4533 33560 4539 33575
rect 4421 33493 4427 33508
rect 4533 33493 4539 33508
rect 4421 33426 4427 33441
rect 4533 33426 4539 33441
rect 4473 33374 4487 33380
rect 4421 32714 4539 33374
rect 4421 32680 4427 32714
rect 4461 32680 4499 32714
rect 4533 32680 4539 32714
rect 4421 32641 4539 32680
rect 4421 32607 4427 32641
rect 4461 32607 4499 32641
rect 4533 32607 4539 32641
rect 4421 32568 4539 32607
rect 4421 32534 4427 32568
rect 4461 32534 4499 32568
rect 4533 32534 4539 32568
rect 4421 32495 4539 32534
rect 4421 32461 4427 32495
rect 4461 32461 4499 32495
rect 4533 32461 4539 32495
rect 4421 32422 4539 32461
rect 4421 31892 4427 32422
rect 4533 31892 4539 32422
rect 4421 31826 4427 31840
rect 4533 31826 4539 31840
rect 4421 31760 4427 31774
rect 4533 31760 4539 31774
rect 4421 31694 4427 31708
rect 4533 31694 4539 31708
rect 4421 31627 4427 31642
rect 4533 31627 4539 31642
rect 4421 31560 4427 31575
rect 4533 31560 4539 31575
rect 4421 31493 4427 31508
rect 4533 31493 4539 31508
rect 4421 31426 4427 31441
rect 4533 31426 4539 31441
rect 4473 31374 4487 31380
rect 4421 30714 4539 31374
rect 4421 30680 4427 30714
rect 4461 30680 4499 30714
rect 4533 30680 4539 30714
rect 4421 30641 4539 30680
rect 4421 30607 4427 30641
rect 4461 30607 4499 30641
rect 4533 30607 4539 30641
rect 4421 30568 4539 30607
rect 4421 30534 4427 30568
rect 4461 30534 4499 30568
rect 4533 30534 4539 30568
rect 4421 30495 4539 30534
rect 4421 30461 4427 30495
rect 4461 30461 4499 30495
rect 4533 30461 4539 30495
rect 4421 30422 4539 30461
rect 4421 29892 4427 30422
rect 4533 29892 4539 30422
rect 4421 29826 4427 29840
rect 4533 29826 4539 29840
rect 4421 29760 4427 29774
rect 4533 29760 4539 29774
rect 4421 29694 4427 29708
rect 4533 29694 4539 29708
rect 4421 29627 4427 29642
rect 4533 29627 4539 29642
rect 4421 29560 4427 29575
rect 4533 29560 4539 29575
rect 4421 29493 4427 29508
rect 4533 29493 4539 29508
rect 4421 29426 4427 29441
rect 4533 29426 4539 29441
rect 4473 29374 4487 29380
rect 4421 29368 4539 29374
rect 4839 34720 4957 34726
rect 4891 34668 4905 34720
rect 4839 34654 4957 34668
rect 4891 34602 4905 34654
rect 4839 34588 4957 34602
rect 4891 34536 4905 34588
rect 4839 34534 4845 34536
rect 4879 34534 4917 34536
rect 4951 34534 4957 34536
rect 4839 34522 4957 34534
rect 4891 34470 4905 34522
rect 4839 34461 4845 34470
rect 4879 34461 4917 34470
rect 4951 34461 4957 34470
rect 4839 34456 4957 34461
rect 4891 34422 4905 34456
rect 4839 34390 4845 34404
rect 4951 34390 4957 34404
rect 4839 34323 4845 34338
rect 4951 34323 4957 34338
rect 4839 34256 4845 34271
rect 4951 34256 4957 34271
rect 4839 33380 4845 34204
rect 4951 33380 4957 34204
rect 4839 32720 4957 33380
rect 4891 32668 4905 32720
rect 4839 32654 4957 32668
rect 4891 32602 4905 32654
rect 4839 32588 4957 32602
rect 4891 32536 4905 32588
rect 4839 32534 4845 32536
rect 4879 32534 4917 32536
rect 4951 32534 4957 32536
rect 4839 32522 4957 32534
rect 4891 32470 4905 32522
rect 4839 32461 4845 32470
rect 4879 32461 4917 32470
rect 4951 32461 4957 32470
rect 4839 32456 4957 32461
rect 4891 32422 4905 32456
rect 4839 32390 4845 32404
rect 4951 32390 4957 32404
rect 4839 32323 4845 32338
rect 4951 32323 4957 32338
rect 4839 32256 4845 32271
rect 4951 32256 4957 32271
rect 4839 31380 4845 32204
rect 4951 31380 4957 32204
rect 4839 30720 4957 31380
rect 4891 30668 4905 30720
rect 4839 30654 4957 30668
rect 4891 30602 4905 30654
rect 4839 30588 4957 30602
rect 4891 30536 4905 30588
rect 4839 30534 4845 30536
rect 4879 30534 4917 30536
rect 4951 30534 4957 30536
rect 4839 30522 4957 30534
rect 4891 30470 4905 30522
rect 4839 30461 4845 30470
rect 4879 30461 4917 30470
rect 4951 30461 4957 30470
rect 4839 30456 4957 30461
rect 4891 30422 4905 30456
rect 4839 30390 4845 30404
rect 4951 30390 4957 30404
rect 4839 30323 4845 30338
rect 4951 30323 4957 30338
rect 4839 30256 4845 30271
rect 4951 30256 4957 30271
rect 4839 29380 4845 30204
rect 4951 29380 4957 30204
rect 2667 29286 2674 29320
rect 2708 29286 2750 29320
rect 2784 29286 2826 29320
rect 2860 29286 2867 29320
rect 2667 29239 2867 29286
rect 2667 29205 2674 29239
rect 2708 29205 2750 29239
rect 2784 29205 2826 29239
rect 2860 29205 2867 29239
rect 2667 29157 2867 29205
rect 2667 29123 2674 29157
rect 2708 29123 2750 29157
rect 2784 29123 2826 29157
rect 2860 29123 2867 29157
rect 2667 29068 2867 29123
tri 2867 29068 3012 29213 sw
rect 2667 28868 4532 29068
tri 4170 28714 4324 28868 ne
rect 4324 28714 4532 28868
tri 4324 28706 4332 28714 ne
tri 1638 28568 1672 28602 sw
rect 1520 28554 3760 28568
tri 1520 28534 1540 28554 ne
rect 1540 28534 3760 28554
tri 3760 28534 3794 28568 sw
tri 1540 28495 1579 28534 ne
rect 1579 28495 3794 28534
tri 3794 28495 3833 28534 sw
tri 1579 28461 1613 28495 ne
rect 1613 28461 3833 28495
tri 3833 28461 3867 28495 sw
tri 1613 28450 1624 28461 ne
rect 1624 28450 3867 28461
tri 3703 28444 3709 28450 ne
rect 3709 28444 3867 28450
tri 3867 28444 3884 28461 sw
tri 3709 28422 3731 28444 ne
rect 3731 28422 3884 28444
tri 3731 28397 3756 28422 ne
rect 3756 23697 3884 28422
rect 3756 23645 3757 23697
rect 3809 23645 3831 23697
rect 3883 23645 3884 23697
rect 3756 23625 3884 23645
rect 3756 23573 3757 23625
rect 3809 23573 3831 23625
rect 3883 23573 3884 23625
rect 3756 23553 3884 23573
rect 3756 23501 3757 23553
rect 3809 23501 3831 23553
rect 3883 23501 3884 23553
rect 3756 23480 3884 23501
rect 3756 23428 3757 23480
rect 3809 23428 3831 23480
rect 3883 23428 3884 23480
rect 3756 21775 3884 23428
rect 3756 21723 3762 21775
rect 3814 21723 3826 21775
rect 3878 21723 3884 21775
tri 3729 20465 3756 20492 se
rect 3756 20465 3884 21723
tri 3721 20457 3729 20465 se
rect 3729 20457 3884 20465
tri 420 20423 454 20457 se
rect 454 20445 3884 20457
rect 454 20423 3862 20445
tri 3862 20423 3884 20445 nw
rect 4332 27321 4532 28714
rect 4332 27287 4339 27321
rect 4373 27287 4415 27321
rect 4449 27287 4491 27321
rect 4525 27287 4532 27321
rect 4332 27244 4532 27287
rect 4332 27210 4339 27244
rect 4373 27210 4415 27244
rect 4449 27210 4491 27244
rect 4525 27210 4532 27244
rect 4332 27167 4532 27210
rect 4332 27133 4339 27167
rect 4373 27133 4415 27167
rect 4449 27133 4491 27167
rect 4525 27133 4532 27167
rect 4332 27089 4532 27133
rect 4332 27055 4339 27089
rect 4373 27055 4415 27089
rect 4449 27055 4491 27089
rect 4525 27055 4532 27089
rect 4332 27011 4532 27055
rect 4332 26977 4339 27011
rect 4373 26977 4415 27011
rect 4449 26977 4491 27011
rect 4525 26977 4532 27011
rect 4332 26933 4532 26977
rect 4332 26899 4339 26933
rect 4373 26899 4415 26933
rect 4449 26899 4491 26933
rect 4525 26899 4532 26933
rect 4332 26855 4532 26899
rect 4332 26821 4339 26855
rect 4373 26821 4415 26855
rect 4449 26821 4491 26855
rect 4525 26821 4532 26855
rect 4332 25670 4532 26821
rect 4839 28720 4957 29380
rect 4891 28668 4905 28720
rect 4839 28654 4957 28668
rect 4891 28602 4905 28654
rect 4839 28588 4957 28602
rect 4891 28536 4905 28588
rect 4839 28534 4845 28536
rect 4879 28534 4917 28536
rect 4951 28534 4957 28536
rect 4839 28522 4957 28534
rect 4891 28470 4905 28522
rect 4839 28461 4845 28470
rect 4879 28461 4917 28470
rect 4951 28461 4957 28470
rect 4839 28456 4957 28461
rect 4891 28422 4905 28456
rect 4839 28390 4845 28404
rect 4951 28390 4957 28404
rect 4839 28323 4845 28338
rect 4951 28323 4957 28338
rect 4839 28256 4845 28271
rect 4951 28256 4957 28271
rect 4839 27380 4845 28204
rect 4951 27380 4957 28204
rect 4839 26752 4957 27380
rect 4839 26720 4845 26752
rect 4879 26720 4917 26752
rect 4951 26720 4957 26752
rect 4891 26668 4905 26720
rect 4839 26654 4845 26668
rect 4879 26654 4917 26668
rect 4951 26654 4957 26668
rect 4891 26602 4905 26654
rect 4839 26588 4845 26602
rect 4879 26588 4917 26602
rect 4951 26588 4957 26602
rect 4891 26536 4905 26588
rect 4839 26527 4957 26536
rect 4839 26522 4845 26527
rect 4879 26522 4917 26527
rect 4951 26522 4957 26527
rect 4891 26470 4905 26522
rect 4839 26456 4957 26470
rect 4891 26404 4905 26456
rect 4839 26389 4957 26404
rect 4891 26337 4905 26389
rect 4839 26322 4957 26337
rect 4891 26270 4905 26322
rect 4839 26268 4845 26270
rect 4879 26268 4917 26270
rect 4951 26268 4957 26270
rect 4839 26255 4957 26268
rect 4891 26203 4905 26255
rect 4839 26193 4845 26203
rect 4879 26193 4917 26203
rect 4951 26193 4957 26203
rect 4839 26152 4957 26193
rect 4839 26118 4845 26152
rect 4879 26118 4917 26152
rect 4951 26118 4957 26152
rect 4839 26077 4957 26118
rect 4839 26043 4845 26077
rect 4879 26043 4917 26077
rect 4951 26043 4957 26077
rect 4839 26002 4957 26043
rect 4839 25968 4845 26002
rect 4879 25968 4917 26002
rect 4951 25968 4957 26002
rect 4839 25928 4957 25968
rect 4839 25894 4845 25928
rect 4879 25894 4917 25928
rect 4951 25894 4957 25928
rect 4839 25854 4957 25894
rect 4839 25820 4845 25854
rect 4879 25820 4917 25854
rect 4951 25820 4957 25854
rect 4839 25780 4957 25820
rect 4839 25746 4845 25780
rect 4879 25746 4917 25780
rect 4951 25746 4957 25780
rect 4839 25732 4957 25746
rect 5257 34714 5375 34891
tri 5375 34821 5445 34891 nw
tri 6023 34821 6093 34891 ne
rect 5257 34680 5263 34714
rect 5297 34680 5335 34714
rect 5369 34680 5375 34714
rect 5257 34641 5375 34680
rect 5257 34607 5263 34641
rect 5297 34607 5335 34641
rect 5369 34607 5375 34641
rect 5257 34568 5375 34607
rect 5257 34534 5263 34568
rect 5297 34534 5335 34568
rect 5369 34534 5375 34568
rect 5257 34495 5375 34534
rect 5257 34461 5263 34495
rect 5297 34461 5335 34495
rect 5369 34461 5375 34495
rect 5257 34422 5375 34461
rect 5257 33892 5263 34422
rect 5369 33892 5375 34422
rect 5257 33826 5263 33840
rect 5369 33826 5375 33840
rect 5257 33760 5263 33774
rect 5369 33760 5375 33774
rect 5257 33694 5263 33708
rect 5369 33694 5375 33708
rect 5257 33627 5263 33642
rect 5369 33627 5375 33642
rect 5257 33560 5263 33575
rect 5369 33560 5375 33575
rect 5257 33493 5263 33508
rect 5369 33493 5375 33508
rect 5257 33426 5263 33441
rect 5369 33426 5375 33441
rect 5309 33374 5323 33380
rect 5257 32714 5375 33374
rect 5257 32680 5263 32714
rect 5297 32680 5335 32714
rect 5369 32680 5375 32714
rect 5257 32641 5375 32680
rect 5257 32607 5263 32641
rect 5297 32607 5335 32641
rect 5369 32607 5375 32641
rect 5257 32568 5375 32607
rect 5257 32534 5263 32568
rect 5297 32534 5335 32568
rect 5369 32534 5375 32568
rect 5257 32495 5375 32534
rect 5257 32461 5263 32495
rect 5297 32461 5335 32495
rect 5369 32461 5375 32495
rect 5257 32422 5375 32461
rect 5257 31892 5263 32422
rect 5369 31892 5375 32422
rect 5257 31826 5263 31840
rect 5369 31826 5375 31840
rect 5257 31760 5263 31774
rect 5369 31760 5375 31774
rect 5257 31694 5263 31708
rect 5369 31694 5375 31708
rect 5257 31627 5263 31642
rect 5369 31627 5375 31642
rect 5257 31560 5263 31575
rect 5369 31560 5375 31575
rect 5257 31493 5263 31508
rect 5369 31493 5375 31508
rect 5257 31426 5263 31441
rect 5369 31426 5375 31441
rect 5309 31374 5323 31380
rect 5257 30714 5375 31374
rect 5257 30680 5263 30714
rect 5297 30680 5335 30714
rect 5369 30680 5375 30714
rect 5257 30641 5375 30680
rect 5257 30607 5263 30641
rect 5297 30607 5335 30641
rect 5369 30607 5375 30641
rect 5257 30568 5375 30607
rect 5257 30534 5263 30568
rect 5297 30534 5335 30568
rect 5369 30534 5375 30568
rect 5257 30495 5375 30534
rect 5257 30461 5263 30495
rect 5297 30461 5335 30495
rect 5369 30461 5375 30495
rect 5257 30422 5375 30461
rect 5257 29892 5263 30422
rect 5369 29892 5375 30422
rect 5257 29826 5263 29840
rect 5369 29826 5375 29840
rect 5257 29760 5263 29774
rect 5369 29760 5375 29774
rect 5257 29694 5263 29708
rect 5369 29694 5375 29708
rect 5257 29627 5263 29642
rect 5369 29627 5375 29642
rect 5257 29560 5263 29575
rect 5369 29560 5375 29575
rect 5257 29493 5263 29508
rect 5369 29493 5375 29508
rect 5257 29426 5263 29441
rect 5369 29426 5375 29441
rect 5309 29374 5323 29380
rect 5257 28714 5375 29374
rect 5257 28680 5263 28714
rect 5297 28680 5335 28714
rect 5369 28680 5375 28714
rect 5257 28641 5375 28680
rect 5257 28607 5263 28641
rect 5297 28607 5335 28641
rect 5369 28607 5375 28641
rect 5257 28568 5375 28607
rect 5257 28534 5263 28568
rect 5297 28534 5335 28568
rect 5369 28534 5375 28568
rect 5257 28495 5375 28534
rect 5257 28461 5263 28495
rect 5297 28461 5335 28495
rect 5369 28461 5375 28495
rect 5257 28422 5375 28461
rect 5257 27892 5263 28422
rect 5369 27892 5375 28422
rect 5257 27826 5263 27840
rect 5369 27826 5375 27840
rect 5257 27760 5263 27774
rect 5369 27760 5375 27774
rect 5257 27694 5263 27708
rect 5369 27694 5375 27708
rect 5257 27627 5263 27642
rect 5369 27627 5375 27642
rect 5257 27560 5263 27575
rect 5369 27560 5375 27575
rect 5257 27493 5263 27508
rect 5369 27493 5375 27508
rect 5257 27426 5263 27441
rect 5369 27426 5375 27441
rect 5309 27374 5323 27380
rect 5257 26743 5375 27374
rect 5257 26709 5263 26743
rect 5297 26709 5335 26743
rect 5369 26709 5375 26743
rect 5257 26668 5375 26709
rect 5257 26634 5263 26668
rect 5297 26634 5335 26668
rect 5369 26634 5375 26668
rect 5257 26594 5375 26634
rect 5257 26560 5263 26594
rect 5297 26560 5335 26594
rect 5369 26560 5375 26594
rect 5257 26520 5375 26560
rect 5257 26486 5263 26520
rect 5297 26486 5335 26520
rect 5369 26486 5375 26520
rect 5257 26446 5375 26486
rect 5257 26412 5263 26446
rect 5297 26412 5335 26446
rect 5369 26412 5375 26446
rect 5257 26372 5375 26412
rect 5257 26338 5263 26372
rect 5297 26338 5335 26372
rect 5369 26338 5375 26372
rect 5257 26298 5375 26338
rect 5257 26264 5263 26298
rect 5297 26264 5335 26298
rect 5369 26264 5375 26298
rect 5257 26224 5375 26264
rect 5257 26190 5263 26224
rect 5297 26190 5335 26224
rect 5369 26190 5375 26224
rect 5257 26150 5375 26190
rect 5257 26116 5263 26150
rect 5297 26116 5335 26150
rect 5369 26116 5375 26150
rect 5257 26076 5375 26116
rect 5257 26042 5263 26076
rect 5297 26042 5335 26076
rect 5369 26042 5375 26076
rect 5257 26002 5375 26042
rect 5257 25968 5263 26002
rect 5297 25968 5335 26002
rect 5369 25968 5375 26002
rect 5257 25928 5375 25968
rect 5257 25894 5263 25928
rect 5297 25894 5335 25928
rect 5369 25894 5375 25928
rect 5257 25891 5375 25894
rect 5309 25839 5323 25891
rect 5257 25825 5263 25839
rect 5297 25825 5335 25839
rect 5369 25825 5375 25839
rect 5309 25773 5323 25825
rect 5257 25759 5263 25773
rect 5297 25759 5335 25773
rect 5369 25759 5375 25773
rect 4332 25636 4344 25670
rect 4378 25636 4486 25670
rect 4520 25636 4532 25670
rect 4332 25071 4532 25636
rect 5309 25707 5323 25759
rect 5675 34720 5793 34726
rect 5727 34668 5741 34720
rect 5675 34654 5793 34668
rect 5727 34602 5741 34654
rect 5675 34588 5793 34602
rect 5727 34536 5741 34588
rect 5675 34534 5681 34536
rect 5715 34534 5753 34536
rect 5787 34534 5793 34536
rect 5675 34522 5793 34534
rect 5727 34470 5741 34522
rect 5675 34461 5681 34470
rect 5715 34461 5753 34470
rect 5787 34461 5793 34470
rect 5675 34456 5793 34461
rect 5727 34422 5741 34456
rect 5675 34390 5681 34404
rect 5787 34390 5793 34404
rect 5675 34323 5681 34338
rect 5787 34323 5793 34338
rect 5675 34256 5681 34271
rect 5787 34256 5793 34271
rect 5675 33380 5681 34204
rect 5787 33380 5793 34204
rect 5675 32720 5793 33380
rect 5727 32668 5741 32720
rect 5675 32654 5793 32668
rect 5727 32602 5741 32654
rect 5675 32588 5793 32602
rect 5727 32536 5741 32588
rect 5675 32534 5681 32536
rect 5715 32534 5753 32536
rect 5787 32534 5793 32536
rect 5675 32522 5793 32534
rect 5727 32470 5741 32522
rect 5675 32461 5681 32470
rect 5715 32461 5753 32470
rect 5787 32461 5793 32470
rect 5675 32456 5793 32461
rect 5727 32422 5741 32456
rect 5675 32390 5681 32404
rect 5787 32390 5793 32404
rect 5675 32323 5681 32338
rect 5787 32323 5793 32338
rect 5675 32256 5681 32271
rect 5787 32256 5793 32271
rect 5675 31380 5681 32204
rect 5787 31380 5793 32204
rect 5675 30720 5793 31380
rect 5727 30668 5741 30720
rect 5675 30654 5793 30668
rect 5727 30602 5741 30654
rect 5675 30588 5793 30602
rect 5727 30536 5741 30588
rect 5675 30534 5681 30536
rect 5715 30534 5753 30536
rect 5787 30534 5793 30536
rect 5675 30522 5793 30534
rect 5727 30470 5741 30522
rect 5675 30461 5681 30470
rect 5715 30461 5753 30470
rect 5787 30461 5793 30470
rect 5675 30456 5793 30461
rect 5727 30422 5741 30456
rect 5675 30390 5681 30404
rect 5787 30390 5793 30404
rect 5675 30323 5681 30338
rect 5787 30323 5793 30338
rect 5675 30256 5681 30271
rect 5787 30256 5793 30271
rect 5675 29380 5681 30204
rect 5787 29380 5793 30204
rect 5675 28720 5793 29380
rect 5727 28668 5741 28720
rect 5675 28654 5793 28668
rect 5727 28602 5741 28654
rect 5675 28588 5793 28602
rect 5727 28536 5741 28588
rect 5675 28534 5681 28536
rect 5715 28534 5753 28536
rect 5787 28534 5793 28536
rect 5675 28522 5793 28534
rect 5727 28470 5741 28522
rect 5675 28461 5681 28470
rect 5715 28461 5753 28470
rect 5787 28461 5793 28470
rect 5675 28456 5793 28461
rect 5727 28422 5741 28456
rect 5675 28390 5681 28404
rect 5787 28390 5793 28404
rect 5675 28323 5681 28338
rect 5787 28323 5793 28338
rect 5675 28256 5681 28271
rect 5787 28256 5793 28271
rect 5675 27380 5681 28204
rect 5787 27380 5793 28204
rect 5675 26752 5793 27380
rect 5675 26720 5681 26752
rect 5715 26720 5753 26752
rect 5787 26720 5793 26752
rect 5727 26668 5741 26720
rect 5675 26654 5681 26668
rect 5715 26654 5753 26668
rect 5787 26654 5793 26668
rect 5727 26602 5741 26654
rect 5675 26588 5681 26602
rect 5715 26588 5753 26602
rect 5787 26588 5793 26602
rect 5727 26536 5741 26588
rect 5675 26533 5793 26536
rect 5675 26522 5681 26533
rect 5715 26522 5753 26533
rect 5787 26522 5793 26533
rect 5727 26470 5741 26522
rect 5675 26460 5793 26470
rect 5675 26456 5681 26460
rect 5715 26456 5753 26460
rect 5787 26456 5793 26460
rect 5727 26404 5741 26456
rect 5675 26389 5793 26404
rect 5727 26337 5741 26389
rect 5675 26322 5793 26337
rect 5727 26270 5741 26322
rect 5675 26255 5793 26270
rect 5727 26203 5741 26255
rect 5675 26168 5793 26203
rect 5675 26134 5681 26168
rect 5715 26134 5753 26168
rect 5787 26134 5793 26168
rect 5675 26095 5793 26134
rect 5675 26061 5681 26095
rect 5715 26061 5753 26095
rect 5787 26061 5793 26095
rect 5675 26022 5793 26061
rect 5675 25772 5681 26022
rect 5787 25772 5793 26022
rect 5675 25732 5793 25772
rect 6093 34714 6211 34891
tri 6211 34821 6281 34891 nw
tri 6859 34821 6929 34891 ne
rect 6093 34680 6099 34714
rect 6133 34680 6171 34714
rect 6205 34680 6211 34714
rect 6093 34641 6211 34680
rect 6093 34607 6099 34641
rect 6133 34607 6171 34641
rect 6205 34607 6211 34641
rect 6093 34568 6211 34607
rect 6093 34534 6099 34568
rect 6133 34534 6171 34568
rect 6205 34534 6211 34568
rect 6093 34495 6211 34534
rect 6093 34461 6099 34495
rect 6133 34461 6171 34495
rect 6205 34461 6211 34495
rect 6093 34422 6211 34461
rect 6093 33892 6099 34422
rect 6205 33892 6211 34422
rect 6093 33826 6099 33840
rect 6205 33826 6211 33840
rect 6093 33760 6099 33774
rect 6205 33760 6211 33774
rect 6093 33694 6099 33708
rect 6205 33694 6211 33708
rect 6093 33627 6099 33642
rect 6205 33627 6211 33642
rect 6093 33560 6099 33575
rect 6205 33560 6211 33575
rect 6093 33493 6099 33508
rect 6205 33493 6211 33508
rect 6093 33426 6099 33441
rect 6205 33426 6211 33441
rect 6145 33374 6159 33380
rect 6093 32714 6211 33374
rect 6093 32680 6099 32714
rect 6133 32680 6171 32714
rect 6205 32680 6211 32714
rect 6093 32641 6211 32680
rect 6093 32607 6099 32641
rect 6133 32607 6171 32641
rect 6205 32607 6211 32641
rect 6093 32568 6211 32607
rect 6093 32534 6099 32568
rect 6133 32534 6171 32568
rect 6205 32534 6211 32568
rect 6093 32495 6211 32534
rect 6093 32461 6099 32495
rect 6133 32461 6171 32495
rect 6205 32461 6211 32495
rect 6093 32422 6211 32461
rect 6093 31892 6099 32422
rect 6205 31892 6211 32422
rect 6093 31826 6099 31840
rect 6205 31826 6211 31840
rect 6093 31760 6099 31774
rect 6205 31760 6211 31774
rect 6093 31694 6099 31708
rect 6205 31694 6211 31708
rect 6093 31627 6099 31642
rect 6205 31627 6211 31642
rect 6093 31560 6099 31575
rect 6205 31560 6211 31575
rect 6093 31493 6099 31508
rect 6205 31493 6211 31508
rect 6093 31426 6099 31441
rect 6205 31426 6211 31441
rect 6145 31374 6159 31380
rect 6093 30714 6211 31374
rect 6093 30680 6099 30714
rect 6133 30680 6171 30714
rect 6205 30680 6211 30714
rect 6093 30641 6211 30680
rect 6093 30607 6099 30641
rect 6133 30607 6171 30641
rect 6205 30607 6211 30641
rect 6093 30568 6211 30607
rect 6093 30534 6099 30568
rect 6133 30534 6171 30568
rect 6205 30534 6211 30568
rect 6093 30495 6211 30534
rect 6093 30461 6099 30495
rect 6133 30461 6171 30495
rect 6205 30461 6211 30495
rect 6093 30422 6211 30461
rect 6093 29892 6099 30422
rect 6205 29892 6211 30422
rect 6093 29826 6099 29840
rect 6205 29826 6211 29840
rect 6093 29760 6099 29774
rect 6205 29760 6211 29774
rect 6093 29694 6099 29708
rect 6205 29694 6211 29708
rect 6093 29627 6099 29642
rect 6205 29627 6211 29642
rect 6093 29560 6099 29575
rect 6205 29560 6211 29575
rect 6093 29493 6099 29508
rect 6205 29493 6211 29508
rect 6093 29426 6099 29441
rect 6205 29426 6211 29441
rect 6145 29374 6159 29380
rect 6093 28714 6211 29374
rect 6093 28680 6099 28714
rect 6133 28680 6171 28714
rect 6205 28680 6211 28714
rect 6093 28641 6211 28680
rect 6093 28607 6099 28641
rect 6133 28607 6171 28641
rect 6205 28607 6211 28641
rect 6093 28568 6211 28607
rect 6093 28534 6099 28568
rect 6133 28534 6171 28568
rect 6205 28534 6211 28568
rect 6093 28495 6211 28534
rect 6093 28461 6099 28495
rect 6133 28461 6171 28495
rect 6205 28461 6211 28495
rect 6093 28422 6211 28461
rect 6093 27892 6099 28422
rect 6205 27892 6211 28422
rect 6093 27826 6099 27840
rect 6205 27826 6211 27840
rect 6093 27760 6099 27774
rect 6205 27760 6211 27774
rect 6093 27694 6099 27708
rect 6205 27694 6211 27708
rect 6093 27627 6099 27642
rect 6205 27627 6211 27642
rect 6093 27560 6099 27575
rect 6205 27560 6211 27575
rect 6093 27493 6099 27508
rect 6205 27493 6211 27508
rect 6093 27426 6099 27441
rect 6205 27426 6211 27441
rect 6145 27374 6159 27380
rect 6093 26743 6211 27374
rect 6093 26709 6099 26743
rect 6133 26709 6171 26743
rect 6205 26709 6211 26743
rect 6093 26668 6211 26709
rect 6093 26634 6099 26668
rect 6133 26634 6171 26668
rect 6205 26634 6211 26668
rect 6093 26594 6211 26634
rect 6093 26560 6099 26594
rect 6133 26560 6171 26594
rect 6205 26560 6211 26594
rect 6093 26520 6211 26560
rect 6093 26486 6099 26520
rect 6133 26486 6171 26520
rect 6205 26486 6211 26520
rect 6093 26446 6211 26486
rect 6093 26412 6099 26446
rect 6133 26412 6171 26446
rect 6205 26412 6211 26446
rect 6093 26372 6211 26412
rect 6093 26338 6099 26372
rect 6133 26338 6171 26372
rect 6205 26338 6211 26372
rect 6093 26298 6211 26338
rect 6093 26264 6099 26298
rect 6133 26264 6171 26298
rect 6205 26264 6211 26298
rect 6093 26224 6211 26264
rect 6093 26190 6099 26224
rect 6133 26190 6171 26224
rect 6205 26190 6211 26224
rect 6093 26150 6211 26190
rect 6093 26116 6099 26150
rect 6133 26116 6171 26150
rect 6205 26116 6211 26150
rect 6093 26076 6211 26116
rect 6093 26042 6099 26076
rect 6133 26042 6171 26076
rect 6205 26042 6211 26076
rect 6093 26002 6211 26042
rect 6093 25968 6099 26002
rect 6133 25968 6171 26002
rect 6205 25968 6211 26002
rect 6093 25928 6211 25968
rect 6093 25894 6099 25928
rect 6133 25894 6171 25928
rect 6205 25894 6211 25928
rect 6093 25891 6211 25894
rect 6145 25839 6159 25891
rect 6093 25825 6099 25839
rect 6133 25825 6171 25839
rect 6205 25825 6211 25839
rect 6145 25773 6159 25825
rect 6093 25759 6099 25773
rect 6133 25759 6171 25773
rect 6205 25759 6211 25773
rect 5257 25693 5375 25707
rect 5309 25641 5323 25693
rect 5257 25626 5375 25641
rect 5309 25574 5323 25626
rect 5257 25559 5375 25574
rect 5309 25507 5323 25559
rect 5257 25492 5375 25507
rect 5309 25440 5323 25492
rect 5257 25425 5375 25440
rect 5309 25373 5323 25425
rect 5257 25367 5375 25373
rect 6145 25707 6159 25759
rect 6511 34720 6629 34726
rect 6563 34668 6577 34720
rect 6511 34654 6629 34668
rect 6563 34602 6577 34654
rect 6511 34588 6629 34602
rect 6563 34536 6577 34588
rect 6511 34534 6517 34536
rect 6551 34534 6589 34536
rect 6623 34534 6629 34536
rect 6511 34522 6629 34534
rect 6563 34470 6577 34522
rect 6511 34461 6517 34470
rect 6551 34461 6589 34470
rect 6623 34461 6629 34470
rect 6511 34456 6629 34461
rect 6563 34422 6577 34456
rect 6511 34390 6517 34404
rect 6623 34390 6629 34404
rect 6511 34323 6517 34338
rect 6623 34323 6629 34338
rect 6511 34256 6517 34271
rect 6623 34256 6629 34271
rect 6511 33380 6517 34204
rect 6623 33380 6629 34204
rect 6511 32720 6629 33380
rect 6563 32668 6577 32720
rect 6511 32654 6629 32668
rect 6563 32602 6577 32654
rect 6511 32588 6629 32602
rect 6563 32536 6577 32588
rect 6511 32534 6517 32536
rect 6551 32534 6589 32536
rect 6623 32534 6629 32536
rect 6511 32522 6629 32534
rect 6563 32470 6577 32522
rect 6511 32461 6517 32470
rect 6551 32461 6589 32470
rect 6623 32461 6629 32470
rect 6511 32456 6629 32461
rect 6563 32422 6577 32456
rect 6511 32390 6517 32404
rect 6623 32390 6629 32404
rect 6511 32323 6517 32338
rect 6623 32323 6629 32338
rect 6511 32256 6517 32271
rect 6623 32256 6629 32271
rect 6511 31380 6517 32204
rect 6623 31380 6629 32204
rect 6511 30720 6629 31380
rect 6563 30668 6577 30720
rect 6511 30654 6629 30668
rect 6563 30602 6577 30654
rect 6511 30588 6629 30602
rect 6563 30536 6577 30588
rect 6511 30534 6517 30536
rect 6551 30534 6589 30536
rect 6623 30534 6629 30536
rect 6511 30522 6629 30534
rect 6563 30470 6577 30522
rect 6511 30461 6517 30470
rect 6551 30461 6589 30470
rect 6623 30461 6629 30470
rect 6511 30456 6629 30461
rect 6563 30422 6577 30456
rect 6511 30390 6517 30404
rect 6623 30390 6629 30404
rect 6511 30323 6517 30338
rect 6623 30323 6629 30338
rect 6511 30256 6517 30271
rect 6623 30256 6629 30271
rect 6511 29380 6517 30204
rect 6623 29380 6629 30204
rect 6511 28720 6629 29380
rect 6563 28668 6577 28720
rect 6511 28654 6629 28668
rect 6563 28602 6577 28654
rect 6511 28588 6629 28602
rect 6563 28536 6577 28588
rect 6511 28534 6517 28536
rect 6551 28534 6589 28536
rect 6623 28534 6629 28536
rect 6511 28522 6629 28534
rect 6563 28470 6577 28522
rect 6511 28461 6517 28470
rect 6551 28461 6589 28470
rect 6623 28461 6629 28470
rect 6511 28456 6629 28461
rect 6563 28422 6577 28456
rect 6511 28390 6517 28404
rect 6623 28390 6629 28404
rect 6511 28323 6517 28338
rect 6623 28323 6629 28338
rect 6511 28256 6517 28271
rect 6623 28256 6629 28271
rect 6511 27380 6517 28204
rect 6623 27380 6629 28204
rect 6511 26751 6629 27380
rect 6511 26720 6517 26751
rect 6551 26720 6589 26751
rect 6623 26720 6629 26751
rect 6563 26668 6577 26720
rect 6511 26654 6517 26668
rect 6551 26654 6589 26668
rect 6623 26654 6629 26668
rect 6563 26602 6577 26654
rect 6511 26601 6629 26602
rect 6511 26588 6517 26601
rect 6551 26588 6589 26601
rect 6623 26588 6629 26601
rect 6563 26536 6577 26588
rect 6511 26526 6629 26536
rect 6511 26522 6517 26526
rect 6551 26522 6589 26526
rect 6623 26522 6629 26526
rect 6563 26470 6577 26522
rect 6511 26456 6629 26470
rect 6563 26404 6577 26456
rect 6511 26389 6629 26404
rect 6563 26337 6577 26389
rect 6511 26322 6629 26337
rect 6563 26270 6577 26322
rect 6511 26267 6517 26270
rect 6551 26267 6589 26270
rect 6623 26267 6629 26270
rect 6511 26255 6629 26267
rect 6563 26203 6577 26255
rect 6511 26192 6517 26203
rect 6551 26192 6589 26203
rect 6623 26192 6629 26203
rect 6511 26151 6629 26192
rect 6511 26117 6517 26151
rect 6551 26117 6589 26151
rect 6623 26117 6629 26151
rect 6511 26076 6629 26117
rect 6511 26042 6517 26076
rect 6551 26042 6589 26076
rect 6623 26042 6629 26076
rect 6511 26002 6629 26042
rect 6511 25968 6517 26002
rect 6551 25968 6589 26002
rect 6623 25968 6629 26002
rect 6511 25928 6629 25968
rect 6511 25894 6517 25928
rect 6551 25894 6589 25928
rect 6623 25894 6629 25928
rect 6511 25854 6629 25894
rect 6511 25820 6517 25854
rect 6551 25820 6589 25854
rect 6623 25820 6629 25854
rect 6511 25780 6629 25820
rect 6511 25746 6517 25780
rect 6551 25746 6589 25780
rect 6623 25746 6629 25780
rect 6511 25732 6629 25746
rect 6929 34714 7047 34891
tri 7047 34821 7117 34891 nw
tri 7695 34821 7765 34891 ne
rect 6929 34680 6935 34714
rect 6969 34680 7007 34714
rect 7041 34680 7047 34714
rect 6929 34641 7047 34680
rect 6929 34607 6935 34641
rect 6969 34607 7007 34641
rect 7041 34607 7047 34641
rect 6929 34568 7047 34607
rect 6929 34534 6935 34568
rect 6969 34534 7007 34568
rect 7041 34534 7047 34568
rect 6929 34495 7047 34534
rect 6929 34461 6935 34495
rect 6969 34461 7007 34495
rect 7041 34461 7047 34495
rect 6929 34422 7047 34461
rect 6929 33892 6935 34422
rect 7041 33892 7047 34422
rect 6929 33826 6935 33840
rect 7041 33826 7047 33840
rect 6929 33760 6935 33774
rect 7041 33760 7047 33774
rect 6929 33694 6935 33708
rect 7041 33694 7047 33708
rect 6929 33627 6935 33642
rect 7041 33627 7047 33642
rect 6929 33560 6935 33575
rect 7041 33560 7047 33575
rect 6929 33493 6935 33508
rect 7041 33493 7047 33508
rect 6929 33426 6935 33441
rect 7041 33426 7047 33441
rect 6981 33374 6995 33380
rect 6929 32714 7047 33374
rect 6929 32680 6935 32714
rect 6969 32680 7007 32714
rect 7041 32680 7047 32714
rect 6929 32641 7047 32680
rect 6929 32607 6935 32641
rect 6969 32607 7007 32641
rect 7041 32607 7047 32641
rect 6929 32568 7047 32607
rect 6929 32534 6935 32568
rect 6969 32534 7007 32568
rect 7041 32534 7047 32568
rect 6929 32495 7047 32534
rect 6929 32461 6935 32495
rect 6969 32461 7007 32495
rect 7041 32461 7047 32495
rect 6929 32422 7047 32461
rect 6929 31892 6935 32422
rect 7041 31892 7047 32422
rect 6929 31826 6935 31840
rect 7041 31826 7047 31840
rect 6929 31760 6935 31774
rect 7041 31760 7047 31774
rect 6929 31694 6935 31708
rect 7041 31694 7047 31708
rect 6929 31627 6935 31642
rect 7041 31627 7047 31642
rect 6929 31560 6935 31575
rect 7041 31560 7047 31575
rect 6929 31493 6935 31508
rect 7041 31493 7047 31508
rect 6929 31426 6935 31441
rect 7041 31426 7047 31441
rect 6981 31374 6995 31380
rect 6929 30714 7047 31374
rect 6929 30680 6935 30714
rect 6969 30680 7007 30714
rect 7041 30680 7047 30714
rect 6929 30641 7047 30680
rect 6929 30607 6935 30641
rect 6969 30607 7007 30641
rect 7041 30607 7047 30641
rect 6929 30568 7047 30607
rect 6929 30534 6935 30568
rect 6969 30534 7007 30568
rect 7041 30534 7047 30568
rect 6929 30495 7047 30534
rect 6929 30461 6935 30495
rect 6969 30461 7007 30495
rect 7041 30461 7047 30495
rect 6929 30422 7047 30461
rect 6929 29892 6935 30422
rect 7041 29892 7047 30422
rect 6929 29826 6935 29840
rect 7041 29826 7047 29840
rect 6929 29760 6935 29774
rect 7041 29760 7047 29774
rect 6929 29694 6935 29708
rect 7041 29694 7047 29708
rect 6929 29627 6935 29642
rect 7041 29627 7047 29642
rect 6929 29560 6935 29575
rect 7041 29560 7047 29575
rect 6929 29493 6935 29508
rect 7041 29493 7047 29508
rect 6929 29426 6935 29441
rect 7041 29426 7047 29441
rect 6981 29374 6995 29380
rect 6929 28714 7047 29374
rect 6929 28680 6935 28714
rect 6969 28680 7007 28714
rect 7041 28680 7047 28714
rect 6929 28641 7047 28680
rect 6929 28607 6935 28641
rect 6969 28607 7007 28641
rect 7041 28607 7047 28641
rect 6929 28568 7047 28607
rect 6929 28534 6935 28568
rect 6969 28534 7007 28568
rect 7041 28534 7047 28568
rect 6929 28495 7047 28534
rect 6929 28461 6935 28495
rect 6969 28461 7007 28495
rect 7041 28461 7047 28495
rect 6929 28422 7047 28461
rect 6929 27892 6935 28422
rect 7041 27892 7047 28422
rect 6929 27826 6935 27840
rect 7041 27826 7047 27840
rect 6929 27760 6935 27774
rect 7041 27760 7047 27774
rect 6929 27694 6935 27708
rect 7041 27694 7047 27708
rect 6929 27627 6935 27642
rect 7041 27627 7047 27642
rect 6929 27560 6935 27575
rect 7041 27560 7047 27575
rect 6929 27493 6935 27508
rect 7041 27493 7047 27508
rect 6929 27426 6935 27441
rect 7041 27426 7047 27441
rect 6981 27374 6995 27380
rect 6929 26768 7047 27374
rect 6929 26734 6935 26768
rect 6969 26734 7007 26768
rect 7041 26734 7047 26768
rect 6929 26692 7047 26734
rect 6929 26658 6935 26692
rect 6969 26658 7007 26692
rect 7041 26658 7047 26692
rect 6929 26616 7047 26658
rect 6929 26582 6935 26616
rect 6969 26582 7007 26616
rect 7041 26582 7047 26616
rect 6929 26540 7047 26582
rect 6929 26506 6935 26540
rect 6969 26506 7007 26540
rect 7041 26506 7047 26540
rect 6929 26464 7047 26506
rect 6929 26430 6935 26464
rect 6969 26430 7007 26464
rect 7041 26430 7047 26464
rect 6929 26388 7047 26430
rect 6929 26354 6935 26388
rect 6969 26354 7007 26388
rect 7041 26354 7047 26388
rect 6929 26312 7047 26354
rect 6929 26278 6935 26312
rect 6969 26278 7007 26312
rect 7041 26278 7047 26312
rect 6929 26236 7047 26278
rect 6929 26202 6935 26236
rect 6969 26202 7007 26236
rect 7041 26202 7047 26236
rect 6929 26160 7047 26202
rect 6929 26126 6935 26160
rect 6969 26126 7007 26160
rect 7041 26126 7047 26160
rect 6929 26084 7047 26126
rect 6929 26050 6935 26084
rect 6969 26050 7007 26084
rect 7041 26050 7047 26084
rect 6929 26008 7047 26050
rect 6929 25974 6935 26008
rect 6969 25974 7007 26008
rect 7041 25974 7047 26008
rect 6929 25932 7047 25974
rect 6929 25898 6935 25932
rect 6969 25898 7007 25932
rect 7041 25898 7047 25932
rect 6929 25891 7047 25898
rect 6981 25839 6995 25891
rect 6929 25825 6935 25839
rect 6969 25825 7007 25839
rect 7041 25825 7047 25839
rect 6981 25773 6995 25825
rect 6929 25759 6935 25773
rect 6969 25759 7007 25773
rect 7041 25759 7047 25773
rect 6093 25693 6211 25707
rect 6145 25641 6159 25693
rect 6093 25626 6211 25641
rect 6145 25574 6159 25626
rect 6093 25559 6211 25574
rect 6145 25507 6159 25559
rect 6093 25492 6211 25507
rect 6145 25440 6159 25492
rect 6093 25425 6211 25440
rect 6145 25373 6159 25425
rect 6093 25367 6211 25373
rect 6981 25707 6995 25759
rect 7347 34720 7465 34726
rect 7399 34668 7413 34720
rect 7347 34654 7465 34668
rect 7399 34602 7413 34654
rect 7347 34588 7465 34602
rect 7399 34536 7413 34588
rect 7347 34534 7353 34536
rect 7387 34534 7425 34536
rect 7459 34534 7465 34536
rect 7347 34522 7465 34534
rect 7399 34470 7413 34522
rect 7347 34461 7353 34470
rect 7387 34461 7425 34470
rect 7459 34461 7465 34470
rect 7347 34456 7465 34461
rect 7399 34422 7413 34456
rect 7347 34390 7353 34404
rect 7459 34390 7465 34404
rect 7347 34323 7353 34338
rect 7459 34323 7465 34338
rect 7347 34256 7353 34271
rect 7459 34256 7465 34271
rect 7347 33380 7353 34204
rect 7459 33380 7465 34204
rect 7347 32720 7465 33380
rect 7399 32668 7413 32720
rect 7347 32654 7465 32668
rect 7399 32602 7413 32654
rect 7347 32588 7465 32602
rect 7399 32536 7413 32588
rect 7347 32534 7353 32536
rect 7387 32534 7425 32536
rect 7459 32534 7465 32536
rect 7347 32522 7465 32534
rect 7399 32470 7413 32522
rect 7347 32461 7353 32470
rect 7387 32461 7425 32470
rect 7459 32461 7465 32470
rect 7347 32456 7465 32461
rect 7399 32422 7413 32456
rect 7347 32390 7353 32404
rect 7459 32390 7465 32404
rect 7347 32323 7353 32338
rect 7459 32323 7465 32338
rect 7347 32256 7353 32271
rect 7459 32256 7465 32271
rect 7347 31380 7353 32204
rect 7459 31380 7465 32204
rect 7347 30720 7465 31380
rect 7399 30668 7413 30720
rect 7347 30654 7465 30668
rect 7399 30602 7413 30654
rect 7347 30588 7465 30602
rect 7399 30536 7413 30588
rect 7347 30534 7353 30536
rect 7387 30534 7425 30536
rect 7459 30534 7465 30536
rect 7347 30522 7465 30534
rect 7399 30470 7413 30522
rect 7347 30461 7353 30470
rect 7387 30461 7425 30470
rect 7459 30461 7465 30470
rect 7347 30456 7465 30461
rect 7399 30422 7413 30456
rect 7347 30390 7353 30404
rect 7459 30390 7465 30404
rect 7347 30323 7353 30338
rect 7459 30323 7465 30338
rect 7347 30256 7353 30271
rect 7459 30256 7465 30271
rect 7347 29380 7353 30204
rect 7459 29380 7465 30204
rect 7347 28720 7465 29380
rect 7399 28668 7413 28720
rect 7347 28654 7465 28668
rect 7399 28602 7413 28654
rect 7347 28588 7465 28602
rect 7399 28536 7413 28588
rect 7347 28534 7353 28536
rect 7387 28534 7425 28536
rect 7459 28534 7465 28536
rect 7347 28522 7465 28534
rect 7399 28470 7413 28522
rect 7347 28461 7353 28470
rect 7387 28461 7425 28470
rect 7459 28461 7465 28470
rect 7347 28456 7465 28461
rect 7399 28422 7413 28456
rect 7347 28390 7353 28404
rect 7459 28390 7465 28404
rect 7347 28323 7353 28338
rect 7459 28323 7465 28338
rect 7347 28256 7353 28271
rect 7459 28256 7465 28271
rect 7347 27380 7353 28204
rect 7459 27380 7465 28204
rect 7347 26751 7465 27380
rect 7347 26720 7353 26751
rect 7387 26720 7425 26751
rect 7459 26720 7465 26751
rect 7399 26668 7413 26720
rect 7347 26654 7353 26668
rect 7387 26654 7425 26668
rect 7459 26654 7465 26668
rect 7399 26602 7413 26654
rect 7347 26601 7465 26602
rect 7347 26588 7353 26601
rect 7387 26588 7425 26601
rect 7459 26588 7465 26601
rect 7399 26536 7413 26588
rect 7347 26526 7465 26536
rect 7347 26522 7353 26526
rect 7387 26522 7425 26526
rect 7459 26522 7465 26526
rect 7399 26470 7413 26522
rect 7347 26456 7465 26470
rect 7399 26404 7413 26456
rect 7347 26389 7465 26404
rect 7399 26337 7413 26389
rect 7347 26322 7465 26337
rect 7399 26270 7413 26322
rect 7347 26267 7353 26270
rect 7387 26267 7425 26270
rect 7459 26267 7465 26270
rect 7347 26255 7465 26267
rect 7399 26203 7413 26255
rect 7347 26192 7353 26203
rect 7387 26192 7425 26203
rect 7459 26192 7465 26203
rect 7347 26151 7465 26192
rect 7347 26117 7353 26151
rect 7387 26117 7425 26151
rect 7459 26117 7465 26151
rect 7347 26076 7465 26117
rect 7347 26042 7353 26076
rect 7387 26042 7425 26076
rect 7459 26042 7465 26076
rect 7347 26002 7465 26042
rect 7347 25968 7353 26002
rect 7387 25968 7425 26002
rect 7459 25968 7465 26002
rect 7347 25928 7465 25968
rect 7347 25894 7353 25928
rect 7387 25894 7425 25928
rect 7459 25894 7465 25928
rect 7347 25854 7465 25894
rect 7347 25820 7353 25854
rect 7387 25820 7425 25854
rect 7459 25820 7465 25854
rect 7347 25780 7465 25820
rect 7347 25746 7353 25780
rect 7387 25746 7425 25780
rect 7459 25746 7465 25780
rect 7347 25732 7465 25746
rect 7765 34714 7883 34891
tri 7883 34821 7953 34891 nw
tri 8531 34821 8601 34891 ne
rect 7765 34680 7771 34714
rect 7805 34680 7843 34714
rect 7877 34680 7883 34714
rect 7765 34641 7883 34680
rect 7765 34607 7771 34641
rect 7805 34607 7843 34641
rect 7877 34607 7883 34641
rect 7765 34568 7883 34607
rect 7765 34534 7771 34568
rect 7805 34534 7843 34568
rect 7877 34534 7883 34568
rect 7765 34495 7883 34534
rect 7765 34461 7771 34495
rect 7805 34461 7843 34495
rect 7877 34461 7883 34495
rect 7765 34422 7883 34461
rect 7765 33892 7771 34422
rect 7877 33892 7883 34422
rect 7765 33826 7771 33840
rect 7877 33826 7883 33840
rect 7765 33760 7771 33774
rect 7877 33760 7883 33774
rect 7765 33694 7771 33708
rect 7877 33694 7883 33708
rect 7765 33627 7771 33642
rect 7877 33627 7883 33642
rect 7765 33560 7771 33575
rect 7877 33560 7883 33575
rect 7765 33493 7771 33508
rect 7877 33493 7883 33508
rect 7765 33426 7771 33441
rect 7877 33426 7883 33441
rect 7817 33374 7831 33380
rect 7765 32714 7883 33374
rect 7765 32680 7771 32714
rect 7805 32680 7843 32714
rect 7877 32680 7883 32714
rect 7765 32641 7883 32680
rect 7765 32607 7771 32641
rect 7805 32607 7843 32641
rect 7877 32607 7883 32641
rect 7765 32568 7883 32607
rect 7765 32534 7771 32568
rect 7805 32534 7843 32568
rect 7877 32534 7883 32568
rect 7765 32495 7883 32534
rect 7765 32461 7771 32495
rect 7805 32461 7843 32495
rect 7877 32461 7883 32495
rect 7765 32422 7883 32461
rect 7765 31892 7771 32422
rect 7877 31892 7883 32422
rect 7765 31826 7771 31840
rect 7877 31826 7883 31840
rect 7765 31760 7771 31774
rect 7877 31760 7883 31774
rect 7765 31694 7771 31708
rect 7877 31694 7883 31708
rect 7765 31627 7771 31642
rect 7877 31627 7883 31642
rect 7765 31560 7771 31575
rect 7877 31560 7883 31575
rect 7765 31493 7771 31508
rect 7877 31493 7883 31508
rect 7765 31426 7771 31441
rect 7877 31426 7883 31441
rect 7817 31374 7831 31380
rect 7765 30714 7883 31374
rect 7765 30680 7771 30714
rect 7805 30680 7843 30714
rect 7877 30680 7883 30714
rect 7765 30641 7883 30680
rect 7765 30607 7771 30641
rect 7805 30607 7843 30641
rect 7877 30607 7883 30641
rect 7765 30568 7883 30607
rect 7765 30534 7771 30568
rect 7805 30534 7843 30568
rect 7877 30534 7883 30568
rect 7765 30495 7883 30534
rect 7765 30461 7771 30495
rect 7805 30461 7843 30495
rect 7877 30461 7883 30495
rect 7765 30422 7883 30461
rect 7765 29892 7771 30422
rect 7877 29892 7883 30422
rect 7765 29826 7771 29840
rect 7877 29826 7883 29840
rect 7765 29760 7771 29774
rect 7877 29760 7883 29774
rect 7765 29694 7771 29708
rect 7877 29694 7883 29708
rect 7765 29627 7771 29642
rect 7877 29627 7883 29642
rect 7765 29560 7771 29575
rect 7877 29560 7883 29575
rect 7765 29493 7771 29508
rect 7877 29493 7883 29508
rect 7765 29426 7771 29441
rect 7877 29426 7883 29441
rect 7817 29374 7831 29380
rect 7765 28714 7883 29374
rect 7765 28680 7771 28714
rect 7805 28680 7843 28714
rect 7877 28680 7883 28714
rect 7765 28641 7883 28680
rect 7765 28607 7771 28641
rect 7805 28607 7843 28641
rect 7877 28607 7883 28641
rect 7765 28568 7883 28607
rect 7765 28534 7771 28568
rect 7805 28534 7843 28568
rect 7877 28534 7883 28568
rect 7765 28495 7883 28534
rect 7765 28461 7771 28495
rect 7805 28461 7843 28495
rect 7877 28461 7883 28495
rect 7765 28422 7883 28461
rect 7765 27892 7771 28422
rect 7877 27892 7883 28422
rect 7765 27826 7771 27840
rect 7877 27826 7883 27840
rect 7765 27760 7771 27774
rect 7877 27760 7883 27774
rect 7765 27694 7771 27708
rect 7877 27694 7883 27708
rect 7765 27627 7771 27642
rect 7877 27627 7883 27642
rect 7765 27560 7771 27575
rect 7877 27560 7883 27575
rect 7765 27493 7771 27508
rect 7877 27493 7883 27508
rect 7765 27426 7771 27441
rect 7877 27426 7883 27441
rect 7817 27374 7831 27380
rect 7765 26785 7883 27374
rect 7765 26751 7771 26785
rect 7805 26751 7843 26785
rect 7877 26751 7883 26785
rect 7765 26707 7883 26751
rect 7765 26673 7771 26707
rect 7805 26673 7843 26707
rect 7877 26673 7883 26707
rect 7765 26629 7883 26673
rect 7765 26595 7771 26629
rect 7805 26595 7843 26629
rect 7877 26595 7883 26629
rect 7765 26551 7883 26595
rect 7765 26517 7771 26551
rect 7805 26517 7843 26551
rect 7877 26517 7883 26551
rect 7765 26473 7883 26517
rect 7765 26439 7771 26473
rect 7805 26439 7843 26473
rect 7877 26439 7883 26473
rect 7765 26396 7883 26439
rect 7765 26362 7771 26396
rect 7805 26362 7843 26396
rect 7877 26362 7883 26396
rect 7765 26319 7883 26362
rect 7765 26285 7771 26319
rect 7805 26285 7843 26319
rect 7877 26285 7883 26319
rect 7765 26242 7883 26285
rect 7765 26208 7771 26242
rect 7805 26208 7843 26242
rect 7877 26208 7883 26242
rect 7765 26165 7883 26208
rect 7765 26131 7771 26165
rect 7805 26131 7843 26165
rect 7877 26131 7883 26165
rect 7765 26088 7883 26131
rect 7765 26054 7771 26088
rect 7805 26054 7843 26088
rect 7877 26054 7883 26088
rect 7765 26011 7883 26054
rect 7765 25977 7771 26011
rect 7805 25977 7843 26011
rect 7877 25977 7883 26011
rect 7765 25934 7883 25977
rect 7765 25900 7771 25934
rect 7805 25900 7843 25934
rect 7877 25900 7883 25934
rect 7765 25891 7883 25900
rect 7817 25839 7831 25891
rect 7765 25825 7771 25839
rect 7805 25825 7843 25839
rect 7877 25825 7883 25839
rect 7817 25773 7831 25825
rect 7765 25759 7771 25773
rect 7805 25759 7843 25773
rect 7877 25759 7883 25773
rect 6929 25693 7047 25707
rect 6981 25641 6995 25693
rect 6929 25626 7047 25641
rect 6981 25574 6995 25626
rect 6929 25559 7047 25574
rect 6981 25507 6995 25559
rect 6929 25492 7047 25507
rect 6981 25440 6995 25492
rect 6929 25425 7047 25440
rect 6981 25373 6995 25425
rect 6929 25367 7047 25373
rect 7817 25707 7831 25759
rect 8183 34720 8301 34726
rect 8235 34668 8249 34720
rect 8183 34654 8301 34668
rect 8235 34602 8249 34654
rect 8183 34588 8301 34602
rect 8235 34536 8249 34588
rect 8183 34534 8189 34536
rect 8223 34534 8261 34536
rect 8295 34534 8301 34536
rect 8183 34522 8301 34534
rect 8235 34470 8249 34522
rect 8183 34461 8189 34470
rect 8223 34461 8261 34470
rect 8295 34461 8301 34470
rect 8183 34456 8301 34461
rect 8235 34422 8249 34456
rect 8183 34390 8189 34404
rect 8295 34390 8301 34404
rect 8183 34323 8189 34338
rect 8295 34323 8301 34338
rect 8183 34256 8189 34271
rect 8295 34256 8301 34271
rect 8183 33380 8189 34204
rect 8295 33380 8301 34204
rect 8183 32720 8301 33380
rect 8235 32668 8249 32720
rect 8183 32654 8301 32668
rect 8235 32602 8249 32654
rect 8183 32588 8301 32602
rect 8235 32536 8249 32588
rect 8183 32534 8189 32536
rect 8223 32534 8261 32536
rect 8295 32534 8301 32536
rect 8183 32522 8301 32534
rect 8235 32470 8249 32522
rect 8183 32461 8189 32470
rect 8223 32461 8261 32470
rect 8295 32461 8301 32470
rect 8183 32456 8301 32461
rect 8235 32422 8249 32456
rect 8183 32390 8189 32404
rect 8295 32390 8301 32404
rect 8183 32323 8189 32338
rect 8295 32323 8301 32338
rect 8183 32256 8189 32271
rect 8295 32256 8301 32271
rect 8183 31380 8189 32204
rect 8295 31380 8301 32204
rect 8183 30720 8301 31380
rect 8235 30668 8249 30720
rect 8183 30654 8301 30668
rect 8235 30602 8249 30654
rect 8183 30588 8301 30602
rect 8235 30536 8249 30588
rect 8183 30534 8189 30536
rect 8223 30534 8261 30536
rect 8295 30534 8301 30536
rect 8183 30522 8301 30534
rect 8235 30470 8249 30522
rect 8183 30461 8189 30470
rect 8223 30461 8261 30470
rect 8295 30461 8301 30470
rect 8183 30456 8301 30461
rect 8235 30422 8249 30456
rect 8183 30390 8189 30404
rect 8295 30390 8301 30404
rect 8183 30323 8189 30338
rect 8295 30323 8301 30338
rect 8183 30256 8189 30271
rect 8295 30256 8301 30271
rect 8183 29380 8189 30204
rect 8295 29380 8301 30204
rect 8183 28720 8301 29380
rect 8235 28668 8249 28720
rect 8183 28654 8301 28668
rect 8235 28602 8249 28654
rect 8183 28588 8301 28602
rect 8235 28536 8249 28588
rect 8183 28534 8189 28536
rect 8223 28534 8261 28536
rect 8295 28534 8301 28536
rect 8183 28522 8301 28534
rect 8235 28470 8249 28522
rect 8183 28461 8189 28470
rect 8223 28461 8261 28470
rect 8295 28461 8301 28470
rect 8183 28456 8301 28461
rect 8235 28422 8249 28456
rect 8183 28390 8189 28404
rect 8295 28390 8301 28404
rect 8183 28323 8189 28338
rect 8295 28323 8301 28338
rect 8183 28256 8189 28271
rect 8295 28256 8301 28271
rect 8183 27380 8189 28204
rect 8295 27380 8301 28204
rect 8183 26751 8301 27380
rect 8183 26720 8189 26751
rect 8223 26720 8261 26751
rect 8295 26720 8301 26751
rect 8235 26668 8249 26720
rect 8183 26654 8189 26668
rect 8223 26654 8261 26668
rect 8295 26654 8301 26668
rect 8235 26602 8249 26654
rect 8183 26601 8301 26602
rect 8183 26588 8189 26601
rect 8223 26588 8261 26601
rect 8295 26588 8301 26601
rect 8235 26536 8249 26588
rect 8183 26526 8301 26536
rect 8183 26522 8189 26526
rect 8223 26522 8261 26526
rect 8295 26522 8301 26526
rect 8235 26470 8249 26522
rect 8183 26456 8301 26470
rect 8235 26404 8249 26456
rect 8183 26389 8301 26404
rect 8235 26337 8249 26389
rect 8183 26322 8301 26337
rect 8235 26270 8249 26322
rect 8183 26267 8189 26270
rect 8223 26267 8261 26270
rect 8295 26267 8301 26270
rect 8183 26255 8301 26267
rect 8235 26203 8249 26255
rect 8183 26192 8189 26203
rect 8223 26192 8261 26203
rect 8295 26192 8301 26203
rect 8183 26151 8301 26192
rect 8183 26117 8189 26151
rect 8223 26117 8261 26151
rect 8295 26117 8301 26151
rect 8183 26076 8301 26117
rect 8183 26042 8189 26076
rect 8223 26042 8261 26076
rect 8295 26042 8301 26076
rect 8183 26002 8301 26042
rect 8183 25968 8189 26002
rect 8223 25968 8261 26002
rect 8295 25968 8301 26002
rect 8183 25928 8301 25968
rect 8183 25894 8189 25928
rect 8223 25894 8261 25928
rect 8295 25894 8301 25928
rect 8183 25854 8301 25894
rect 8183 25820 8189 25854
rect 8223 25820 8261 25854
rect 8295 25820 8301 25854
rect 8183 25780 8301 25820
rect 8183 25746 8189 25780
rect 8223 25746 8261 25780
rect 8295 25746 8301 25780
rect 8183 25732 8301 25746
rect 8601 34714 8719 34891
tri 8719 34821 8789 34891 nw
tri 9367 34821 9437 34891 ne
rect 8601 34680 8607 34714
rect 8641 34680 8679 34714
rect 8713 34680 8719 34714
rect 8601 34641 8719 34680
rect 8601 34607 8607 34641
rect 8641 34607 8679 34641
rect 8713 34607 8719 34641
rect 8601 34568 8719 34607
rect 8601 34534 8607 34568
rect 8641 34534 8679 34568
rect 8713 34534 8719 34568
rect 8601 34495 8719 34534
rect 8601 34461 8607 34495
rect 8641 34461 8679 34495
rect 8713 34461 8719 34495
rect 8601 34422 8719 34461
rect 8601 33892 8607 34422
rect 8713 33892 8719 34422
rect 8601 33826 8607 33840
rect 8713 33826 8719 33840
rect 8601 33760 8607 33774
rect 8713 33760 8719 33774
rect 8601 33694 8607 33708
rect 8713 33694 8719 33708
rect 8601 33627 8607 33642
rect 8713 33627 8719 33642
rect 8601 33560 8607 33575
rect 8713 33560 8719 33575
rect 8601 33493 8607 33508
rect 8713 33493 8719 33508
rect 8601 33426 8607 33441
rect 8713 33426 8719 33441
rect 8653 33374 8667 33380
rect 8601 32714 8719 33374
rect 8601 32680 8607 32714
rect 8641 32680 8679 32714
rect 8713 32680 8719 32714
rect 8601 32641 8719 32680
rect 8601 32607 8607 32641
rect 8641 32607 8679 32641
rect 8713 32607 8719 32641
rect 8601 32568 8719 32607
rect 8601 32534 8607 32568
rect 8641 32534 8679 32568
rect 8713 32534 8719 32568
rect 8601 32495 8719 32534
rect 8601 32461 8607 32495
rect 8641 32461 8679 32495
rect 8713 32461 8719 32495
rect 8601 32422 8719 32461
rect 8601 31892 8607 32422
rect 8713 31892 8719 32422
rect 8601 31826 8607 31840
rect 8713 31826 8719 31840
rect 8601 31760 8607 31774
rect 8713 31760 8719 31774
rect 8601 31694 8607 31708
rect 8713 31694 8719 31708
rect 8601 31627 8607 31642
rect 8713 31627 8719 31642
rect 8601 31560 8607 31575
rect 8713 31560 8719 31575
rect 8601 31493 8607 31508
rect 8713 31493 8719 31508
rect 8601 31426 8607 31441
rect 8713 31426 8719 31441
rect 8653 31374 8667 31380
rect 8601 30714 8719 31374
rect 8601 30680 8607 30714
rect 8641 30680 8679 30714
rect 8713 30680 8719 30714
rect 8601 30641 8719 30680
rect 8601 30607 8607 30641
rect 8641 30607 8679 30641
rect 8713 30607 8719 30641
rect 8601 30568 8719 30607
rect 8601 30534 8607 30568
rect 8641 30534 8679 30568
rect 8713 30534 8719 30568
rect 8601 30495 8719 30534
rect 8601 30461 8607 30495
rect 8641 30461 8679 30495
rect 8713 30461 8719 30495
rect 8601 30422 8719 30461
rect 8601 29892 8607 30422
rect 8713 29892 8719 30422
rect 8601 29826 8607 29840
rect 8713 29826 8719 29840
rect 8601 29760 8607 29774
rect 8713 29760 8719 29774
rect 8601 29694 8607 29708
rect 8713 29694 8719 29708
rect 8601 29627 8607 29642
rect 8713 29627 8719 29642
rect 8601 29560 8607 29575
rect 8713 29560 8719 29575
rect 8601 29493 8607 29508
rect 8713 29493 8719 29508
rect 8601 29426 8607 29441
rect 8713 29426 8719 29441
rect 8653 29374 8667 29380
rect 8601 28714 8719 29374
rect 8601 28680 8607 28714
rect 8641 28680 8679 28714
rect 8713 28680 8719 28714
rect 8601 28641 8719 28680
rect 8601 28607 8607 28641
rect 8641 28607 8679 28641
rect 8713 28607 8719 28641
rect 8601 28568 8719 28607
rect 8601 28534 8607 28568
rect 8641 28534 8679 28568
rect 8713 28534 8719 28568
rect 8601 28495 8719 28534
rect 8601 28461 8607 28495
rect 8641 28461 8679 28495
rect 8713 28461 8719 28495
rect 8601 28422 8719 28461
rect 8601 27892 8607 28422
rect 8713 27892 8719 28422
rect 8601 27826 8607 27840
rect 8713 27826 8719 27840
rect 8601 27760 8607 27774
rect 8713 27760 8719 27774
rect 8601 27694 8607 27708
rect 8713 27694 8719 27708
rect 8601 27627 8607 27642
rect 8713 27627 8719 27642
rect 8601 27560 8607 27575
rect 8713 27560 8719 27575
rect 8601 27493 8607 27508
rect 8713 27493 8719 27508
rect 8601 27426 8607 27441
rect 8713 27426 8719 27441
rect 8653 27374 8667 27380
rect 8601 26785 8719 27374
rect 8601 26751 8607 26785
rect 8641 26751 8679 26785
rect 8713 26751 8719 26785
rect 8601 26707 8719 26751
rect 8601 26673 8607 26707
rect 8641 26673 8679 26707
rect 8713 26673 8719 26707
rect 8601 26629 8719 26673
rect 8601 26595 8607 26629
rect 8641 26595 8679 26629
rect 8713 26595 8719 26629
rect 8601 26551 8719 26595
rect 8601 26517 8607 26551
rect 8641 26517 8679 26551
rect 8713 26517 8719 26551
rect 8601 26473 8719 26517
rect 8601 26439 8607 26473
rect 8641 26439 8679 26473
rect 8713 26439 8719 26473
rect 8601 26396 8719 26439
rect 8601 26362 8607 26396
rect 8641 26362 8679 26396
rect 8713 26362 8719 26396
rect 8601 26319 8719 26362
rect 8601 26285 8607 26319
rect 8641 26285 8679 26319
rect 8713 26285 8719 26319
rect 8601 26242 8719 26285
rect 8601 26208 8607 26242
rect 8641 26208 8679 26242
rect 8713 26208 8719 26242
rect 8601 26165 8719 26208
rect 8601 26131 8607 26165
rect 8641 26131 8679 26165
rect 8713 26131 8719 26165
rect 8601 26088 8719 26131
rect 8601 26054 8607 26088
rect 8641 26054 8679 26088
rect 8713 26054 8719 26088
rect 8601 26011 8719 26054
rect 8601 25977 8607 26011
rect 8641 25977 8679 26011
rect 8713 25977 8719 26011
rect 8601 25934 8719 25977
rect 8601 25900 8607 25934
rect 8641 25900 8679 25934
rect 8713 25900 8719 25934
rect 8601 25891 8719 25900
rect 8653 25839 8667 25891
rect 8601 25825 8607 25839
rect 8641 25825 8679 25839
rect 8713 25825 8719 25839
rect 8653 25773 8667 25825
rect 8601 25759 8607 25773
rect 8641 25759 8679 25773
rect 8713 25759 8719 25773
rect 7765 25693 7883 25707
rect 7817 25641 7831 25693
rect 7765 25626 7883 25641
rect 7817 25574 7831 25626
rect 7765 25559 7883 25574
rect 7817 25507 7831 25559
rect 7765 25492 7883 25507
rect 7817 25440 7831 25492
rect 7765 25425 7883 25440
rect 7817 25373 7831 25425
rect 7765 25367 7883 25373
rect 8653 25707 8667 25759
rect 9019 34720 9137 34726
rect 9071 34668 9085 34720
rect 9019 34654 9137 34668
rect 9071 34602 9085 34654
rect 9019 34588 9137 34602
rect 9071 34536 9085 34588
rect 9019 34534 9025 34536
rect 9059 34534 9097 34536
rect 9131 34534 9137 34536
rect 9019 34522 9137 34534
rect 9071 34470 9085 34522
rect 9019 34461 9025 34470
rect 9059 34461 9097 34470
rect 9131 34461 9137 34470
rect 9019 34456 9137 34461
rect 9071 34422 9085 34456
rect 9019 34390 9025 34404
rect 9131 34390 9137 34404
rect 9019 34323 9025 34338
rect 9131 34323 9137 34338
rect 9019 34256 9025 34271
rect 9131 34256 9137 34271
rect 9019 33380 9025 34204
rect 9131 33380 9137 34204
rect 9019 32720 9137 33380
rect 9071 32668 9085 32720
rect 9019 32654 9137 32668
rect 9071 32602 9085 32654
rect 9019 32588 9137 32602
rect 9071 32536 9085 32588
rect 9019 32534 9025 32536
rect 9059 32534 9097 32536
rect 9131 32534 9137 32536
rect 9019 32522 9137 32534
rect 9071 32470 9085 32522
rect 9019 32461 9025 32470
rect 9059 32461 9097 32470
rect 9131 32461 9137 32470
rect 9019 32456 9137 32461
rect 9071 32422 9085 32456
rect 9019 32390 9025 32404
rect 9131 32390 9137 32404
rect 9019 32323 9025 32338
rect 9131 32323 9137 32338
rect 9019 32256 9025 32271
rect 9131 32256 9137 32271
rect 9019 31380 9025 32204
rect 9131 31380 9137 32204
rect 9019 30720 9137 31380
rect 9071 30668 9085 30720
rect 9019 30654 9137 30668
rect 9071 30602 9085 30654
rect 9019 30588 9137 30602
rect 9071 30536 9085 30588
rect 9019 30534 9025 30536
rect 9059 30534 9097 30536
rect 9131 30534 9137 30536
rect 9019 30522 9137 30534
rect 9071 30470 9085 30522
rect 9019 30461 9025 30470
rect 9059 30461 9097 30470
rect 9131 30461 9137 30470
rect 9019 30456 9137 30461
rect 9071 30422 9085 30456
rect 9019 30390 9025 30404
rect 9131 30390 9137 30404
rect 9019 30323 9025 30338
rect 9131 30323 9137 30338
rect 9019 30256 9025 30271
rect 9131 30256 9137 30271
rect 9019 29380 9025 30204
rect 9131 29380 9137 30204
rect 9019 28720 9137 29380
rect 9071 28668 9085 28720
rect 9019 28654 9137 28668
rect 9071 28602 9085 28654
rect 9019 28588 9137 28602
rect 9071 28536 9085 28588
rect 9019 28534 9025 28536
rect 9059 28534 9097 28536
rect 9131 28534 9137 28536
rect 9019 28522 9137 28534
rect 9071 28470 9085 28522
rect 9019 28461 9025 28470
rect 9059 28461 9097 28470
rect 9131 28461 9137 28470
rect 9019 28456 9137 28461
rect 9071 28422 9085 28456
rect 9019 28390 9025 28404
rect 9131 28390 9137 28404
rect 9019 28323 9025 28338
rect 9131 28323 9137 28338
rect 9019 28256 9025 28271
rect 9131 28256 9137 28271
rect 9019 27380 9025 28204
rect 9131 27380 9137 28204
rect 9019 26751 9137 27380
rect 9019 26720 9025 26751
rect 9059 26720 9097 26751
rect 9131 26720 9137 26751
rect 9071 26668 9085 26720
rect 9019 26654 9025 26668
rect 9059 26654 9097 26668
rect 9131 26654 9137 26668
rect 9071 26602 9085 26654
rect 9019 26601 9137 26602
rect 9019 26588 9025 26601
rect 9059 26588 9097 26601
rect 9131 26588 9137 26601
rect 9071 26536 9085 26588
rect 9019 26526 9137 26536
rect 9019 26522 9025 26526
rect 9059 26522 9097 26526
rect 9131 26522 9137 26526
rect 9071 26470 9085 26522
rect 9019 26456 9137 26470
rect 9071 26404 9085 26456
rect 9019 26389 9137 26404
rect 9071 26337 9085 26389
rect 9019 26322 9137 26337
rect 9071 26270 9085 26322
rect 9019 26267 9025 26270
rect 9059 26267 9097 26270
rect 9131 26267 9137 26270
rect 9019 26255 9137 26267
rect 9071 26203 9085 26255
rect 9019 26192 9025 26203
rect 9059 26192 9097 26203
rect 9131 26192 9137 26203
rect 9019 26151 9137 26192
rect 9019 26117 9025 26151
rect 9059 26117 9097 26151
rect 9131 26117 9137 26151
rect 9019 26076 9137 26117
rect 9019 26042 9025 26076
rect 9059 26042 9097 26076
rect 9131 26042 9137 26076
rect 9019 26002 9137 26042
rect 9019 25968 9025 26002
rect 9059 25968 9097 26002
rect 9131 25968 9137 26002
rect 9019 25928 9137 25968
rect 9019 25894 9025 25928
rect 9059 25894 9097 25928
rect 9131 25894 9137 25928
rect 9019 25854 9137 25894
rect 9019 25820 9025 25854
rect 9059 25820 9097 25854
rect 9131 25820 9137 25854
rect 9019 25780 9137 25820
rect 9019 25746 9025 25780
rect 9059 25746 9097 25780
rect 9131 25746 9137 25780
rect 9019 25732 9137 25746
rect 9437 34714 9555 34891
tri 9555 34821 9625 34891 nw
tri 10203 34821 10273 34891 ne
rect 9437 34680 9443 34714
rect 9477 34680 9515 34714
rect 9549 34680 9555 34714
rect 9437 34641 9555 34680
rect 9437 34607 9443 34641
rect 9477 34607 9515 34641
rect 9549 34607 9555 34641
rect 9437 34568 9555 34607
rect 9437 34534 9443 34568
rect 9477 34534 9515 34568
rect 9549 34534 9555 34568
rect 9437 34495 9555 34534
rect 9437 34461 9443 34495
rect 9477 34461 9515 34495
rect 9549 34461 9555 34495
rect 9437 34422 9555 34461
rect 9437 33892 9443 34422
rect 9549 33892 9555 34422
rect 9437 33826 9443 33840
rect 9549 33826 9555 33840
rect 9437 33760 9443 33774
rect 9549 33760 9555 33774
rect 9437 33694 9443 33708
rect 9549 33694 9555 33708
rect 9437 33627 9443 33642
rect 9549 33627 9555 33642
rect 9437 33560 9443 33575
rect 9549 33560 9555 33575
rect 9437 33493 9443 33508
rect 9549 33493 9555 33508
rect 9437 33426 9443 33441
rect 9549 33426 9555 33441
rect 9489 33374 9503 33380
rect 9437 32714 9555 33374
rect 9437 32680 9443 32714
rect 9477 32680 9515 32714
rect 9549 32680 9555 32714
rect 9437 32641 9555 32680
rect 9437 32607 9443 32641
rect 9477 32607 9515 32641
rect 9549 32607 9555 32641
rect 9437 32568 9555 32607
rect 9437 32534 9443 32568
rect 9477 32534 9515 32568
rect 9549 32534 9555 32568
rect 9437 32495 9555 32534
rect 9437 32461 9443 32495
rect 9477 32461 9515 32495
rect 9549 32461 9555 32495
rect 9437 32422 9555 32461
rect 9437 31892 9443 32422
rect 9549 31892 9555 32422
rect 9437 31826 9443 31840
rect 9549 31826 9555 31840
rect 9437 31760 9443 31774
rect 9549 31760 9555 31774
rect 9437 31694 9443 31708
rect 9549 31694 9555 31708
rect 9437 31627 9443 31642
rect 9549 31627 9555 31642
rect 9437 31560 9443 31575
rect 9549 31560 9555 31575
rect 9437 31493 9443 31508
rect 9549 31493 9555 31508
rect 9437 31426 9443 31441
rect 9549 31426 9555 31441
rect 9489 31374 9503 31380
rect 9437 30714 9555 31374
rect 9437 30680 9443 30714
rect 9477 30680 9515 30714
rect 9549 30680 9555 30714
rect 9437 30641 9555 30680
rect 9437 30607 9443 30641
rect 9477 30607 9515 30641
rect 9549 30607 9555 30641
rect 9437 30568 9555 30607
rect 9437 30534 9443 30568
rect 9477 30534 9515 30568
rect 9549 30534 9555 30568
rect 9437 30495 9555 30534
rect 9437 30461 9443 30495
rect 9477 30461 9515 30495
rect 9549 30461 9555 30495
rect 9437 30422 9555 30461
rect 9437 29892 9443 30422
rect 9549 29892 9555 30422
rect 9437 29826 9443 29840
rect 9549 29826 9555 29840
rect 9437 29760 9443 29774
rect 9549 29760 9555 29774
rect 9437 29694 9443 29708
rect 9549 29694 9555 29708
rect 9437 29627 9443 29642
rect 9549 29627 9555 29642
rect 9437 29560 9443 29575
rect 9549 29560 9555 29575
rect 9437 29493 9443 29508
rect 9549 29493 9555 29508
rect 9437 29426 9443 29441
rect 9549 29426 9555 29441
rect 9489 29374 9503 29380
rect 9437 28714 9555 29374
rect 9437 28680 9443 28714
rect 9477 28680 9515 28714
rect 9549 28680 9555 28714
rect 9437 28641 9555 28680
rect 9437 28607 9443 28641
rect 9477 28607 9515 28641
rect 9549 28607 9555 28641
rect 9437 28568 9555 28607
rect 9437 28534 9443 28568
rect 9477 28534 9515 28568
rect 9549 28534 9555 28568
rect 9437 28495 9555 28534
rect 9437 28461 9443 28495
rect 9477 28461 9515 28495
rect 9549 28461 9555 28495
rect 9437 28422 9555 28461
rect 9437 27892 9443 28422
rect 9549 27892 9555 28422
rect 9437 27826 9443 27840
rect 9549 27826 9555 27840
rect 9437 27760 9443 27774
rect 9549 27760 9555 27774
rect 9437 27694 9443 27708
rect 9549 27694 9555 27708
rect 9437 27627 9443 27642
rect 9549 27627 9555 27642
rect 9437 27560 9443 27575
rect 9549 27560 9555 27575
rect 9437 27493 9443 27508
rect 9549 27493 9555 27508
rect 9437 27426 9443 27441
rect 9549 27426 9555 27441
rect 9489 27374 9503 27380
rect 9437 26785 9555 27374
rect 9437 26751 9443 26785
rect 9477 26751 9515 26785
rect 9549 26751 9555 26785
rect 9437 26707 9555 26751
rect 9437 26673 9443 26707
rect 9477 26673 9515 26707
rect 9549 26673 9555 26707
rect 9437 26629 9555 26673
rect 9437 26595 9443 26629
rect 9477 26595 9515 26629
rect 9549 26595 9555 26629
rect 9437 26551 9555 26595
rect 9437 26517 9443 26551
rect 9477 26517 9515 26551
rect 9549 26517 9555 26551
rect 9437 26473 9555 26517
rect 9437 26439 9443 26473
rect 9477 26439 9515 26473
rect 9549 26439 9555 26473
rect 9437 26396 9555 26439
rect 9437 26362 9443 26396
rect 9477 26362 9515 26396
rect 9549 26362 9555 26396
rect 9437 26319 9555 26362
rect 9437 26285 9443 26319
rect 9477 26285 9515 26319
rect 9549 26285 9555 26319
rect 9437 26242 9555 26285
rect 9437 26208 9443 26242
rect 9477 26208 9515 26242
rect 9549 26208 9555 26242
rect 9437 26165 9555 26208
rect 9437 26131 9443 26165
rect 9477 26131 9515 26165
rect 9549 26131 9555 26165
rect 9437 26088 9555 26131
rect 9437 26054 9443 26088
rect 9477 26054 9515 26088
rect 9549 26054 9555 26088
rect 9437 26011 9555 26054
rect 9437 25977 9443 26011
rect 9477 25977 9515 26011
rect 9549 25977 9555 26011
rect 9437 25934 9555 25977
rect 9437 25900 9443 25934
rect 9477 25900 9515 25934
rect 9549 25900 9555 25934
rect 9437 25891 9555 25900
rect 9489 25839 9503 25891
rect 9437 25825 9443 25839
rect 9477 25825 9515 25839
rect 9549 25825 9555 25839
rect 9489 25773 9503 25825
rect 9437 25759 9443 25773
rect 9477 25759 9515 25773
rect 9549 25759 9555 25773
rect 8601 25693 8719 25707
rect 8653 25641 8667 25693
rect 8601 25626 8719 25641
rect 8653 25574 8667 25626
rect 8601 25559 8719 25574
rect 8653 25507 8667 25559
rect 8601 25492 8719 25507
rect 8653 25440 8667 25492
rect 8601 25425 8719 25440
rect 8653 25373 8667 25425
rect 8601 25367 8719 25373
rect 9489 25707 9503 25759
rect 9855 34720 9973 34726
rect 9907 34668 9921 34720
rect 9855 34654 9973 34668
rect 9907 34602 9921 34654
rect 9855 34588 9973 34602
rect 9907 34536 9921 34588
rect 9855 34534 9861 34536
rect 9895 34534 9933 34536
rect 9967 34534 9973 34536
rect 9855 34522 9973 34534
rect 9907 34470 9921 34522
rect 9855 34461 9861 34470
rect 9895 34461 9933 34470
rect 9967 34461 9973 34470
rect 9855 34456 9973 34461
rect 9907 34422 9921 34456
rect 9855 34390 9861 34404
rect 9967 34390 9973 34404
rect 9855 34323 9861 34338
rect 9967 34323 9973 34338
rect 9855 34256 9861 34271
rect 9967 34256 9973 34271
rect 9855 33380 9861 34204
rect 9967 33380 9973 34204
rect 9855 32720 9973 33380
rect 9907 32668 9921 32720
rect 9855 32654 9973 32668
rect 9907 32602 9921 32654
rect 9855 32588 9973 32602
rect 9907 32536 9921 32588
rect 9855 32534 9861 32536
rect 9895 32534 9933 32536
rect 9967 32534 9973 32536
rect 9855 32522 9973 32534
rect 9907 32470 9921 32522
rect 9855 32461 9861 32470
rect 9895 32461 9933 32470
rect 9967 32461 9973 32470
rect 9855 32456 9973 32461
rect 9907 32422 9921 32456
rect 9855 32390 9861 32404
rect 9967 32390 9973 32404
rect 9855 32323 9861 32338
rect 9967 32323 9973 32338
rect 9855 32256 9861 32271
rect 9967 32256 9973 32271
rect 9855 31380 9861 32204
rect 9967 31380 9973 32204
rect 9855 30720 9973 31380
rect 9907 30668 9921 30720
rect 9855 30654 9973 30668
rect 9907 30602 9921 30654
rect 9855 30588 9973 30602
rect 9907 30536 9921 30588
rect 9855 30534 9861 30536
rect 9895 30534 9933 30536
rect 9967 30534 9973 30536
rect 9855 30522 9973 30534
rect 9907 30470 9921 30522
rect 9855 30461 9861 30470
rect 9895 30461 9933 30470
rect 9967 30461 9973 30470
rect 9855 30456 9973 30461
rect 9907 30422 9921 30456
rect 9855 30390 9861 30404
rect 9967 30390 9973 30404
rect 9855 30323 9861 30338
rect 9967 30323 9973 30338
rect 9855 30256 9861 30271
rect 9967 30256 9973 30271
rect 9855 29380 9861 30204
rect 9967 29380 9973 30204
rect 9855 28720 9973 29380
rect 9907 28668 9921 28720
rect 9855 28654 9973 28668
rect 9907 28602 9921 28654
rect 9855 28588 9973 28602
rect 9907 28536 9921 28588
rect 9855 28534 9861 28536
rect 9895 28534 9933 28536
rect 9967 28534 9973 28536
rect 9855 28522 9973 28534
rect 9907 28470 9921 28522
rect 9855 28461 9861 28470
rect 9895 28461 9933 28470
rect 9967 28461 9973 28470
rect 9855 28456 9973 28461
rect 9907 28422 9921 28456
rect 9855 28390 9861 28404
rect 9967 28390 9973 28404
rect 9855 28323 9861 28338
rect 9967 28323 9973 28338
rect 9855 28256 9861 28271
rect 9967 28256 9973 28271
rect 9855 27380 9861 28204
rect 9967 27380 9973 28204
rect 9855 26751 9973 27380
rect 9855 26720 9861 26751
rect 9895 26720 9933 26751
rect 9967 26720 9973 26751
rect 9907 26668 9921 26720
rect 9855 26654 9861 26668
rect 9895 26654 9933 26668
rect 9967 26654 9973 26668
rect 9907 26602 9921 26654
rect 9855 26601 9973 26602
rect 9855 26588 9861 26601
rect 9895 26588 9933 26601
rect 9967 26588 9973 26601
rect 9907 26536 9921 26588
rect 9855 26526 9973 26536
rect 9855 26522 9861 26526
rect 9895 26522 9933 26526
rect 9967 26522 9973 26526
rect 9907 26470 9921 26522
rect 9855 26456 9973 26470
rect 9907 26404 9921 26456
rect 9855 26389 9973 26404
rect 9907 26337 9921 26389
rect 9855 26322 9973 26337
rect 9907 26270 9921 26322
rect 9855 26267 9861 26270
rect 9895 26267 9933 26270
rect 9967 26267 9973 26270
rect 9855 26255 9973 26267
rect 9907 26203 9921 26255
rect 9855 26192 9861 26203
rect 9895 26192 9933 26203
rect 9967 26192 9973 26203
rect 9855 26151 9973 26192
rect 9855 26117 9861 26151
rect 9895 26117 9933 26151
rect 9967 26117 9973 26151
rect 9855 26076 9973 26117
rect 9855 26042 9861 26076
rect 9895 26042 9933 26076
rect 9967 26042 9973 26076
rect 9855 26002 9973 26042
rect 9855 25968 9861 26002
rect 9895 25968 9933 26002
rect 9967 25968 9973 26002
rect 9855 25928 9973 25968
rect 9855 25894 9861 25928
rect 9895 25894 9933 25928
rect 9967 25894 9973 25928
rect 9855 25854 9973 25894
rect 9855 25820 9861 25854
rect 9895 25820 9933 25854
rect 9967 25820 9973 25854
rect 9855 25780 9973 25820
rect 9855 25746 9861 25780
rect 9895 25746 9933 25780
rect 9967 25746 9973 25780
rect 9855 25732 9973 25746
rect 10273 34714 10391 34891
tri 10391 34821 10461 34891 nw
tri 11039 34821 11109 34891 ne
rect 10273 34680 10279 34714
rect 10313 34680 10351 34714
rect 10385 34680 10391 34714
rect 10273 34641 10391 34680
rect 10273 34607 10279 34641
rect 10313 34607 10351 34641
rect 10385 34607 10391 34641
rect 10273 34568 10391 34607
rect 10273 34534 10279 34568
rect 10313 34534 10351 34568
rect 10385 34534 10391 34568
rect 10273 34495 10391 34534
rect 10273 34461 10279 34495
rect 10313 34461 10351 34495
rect 10385 34461 10391 34495
rect 10273 34422 10391 34461
rect 10273 33892 10279 34422
rect 10385 33892 10391 34422
rect 10273 33826 10279 33840
rect 10385 33826 10391 33840
rect 10273 33760 10279 33774
rect 10385 33760 10391 33774
rect 10273 33694 10279 33708
rect 10385 33694 10391 33708
rect 10273 33627 10279 33642
rect 10385 33627 10391 33642
rect 10273 33560 10279 33575
rect 10385 33560 10391 33575
rect 10273 33493 10279 33508
rect 10385 33493 10391 33508
rect 10273 33426 10279 33441
rect 10385 33426 10391 33441
rect 10325 33374 10339 33380
rect 10273 32714 10391 33374
rect 10273 32680 10279 32714
rect 10313 32680 10351 32714
rect 10385 32680 10391 32714
rect 10273 32641 10391 32680
rect 10273 32607 10279 32641
rect 10313 32607 10351 32641
rect 10385 32607 10391 32641
rect 10273 32568 10391 32607
rect 10273 32534 10279 32568
rect 10313 32534 10351 32568
rect 10385 32534 10391 32568
rect 10273 32495 10391 32534
rect 10273 32461 10279 32495
rect 10313 32461 10351 32495
rect 10385 32461 10391 32495
rect 10273 32422 10391 32461
rect 10273 31892 10279 32422
rect 10385 31892 10391 32422
rect 10273 31826 10279 31840
rect 10385 31826 10391 31840
rect 10273 31760 10279 31774
rect 10385 31760 10391 31774
rect 10273 31694 10279 31708
rect 10385 31694 10391 31708
rect 10273 31627 10279 31642
rect 10385 31627 10391 31642
rect 10273 31560 10279 31575
rect 10385 31560 10391 31575
rect 10273 31493 10279 31508
rect 10385 31493 10391 31508
rect 10273 31426 10279 31441
rect 10385 31426 10391 31441
rect 10325 31374 10339 31380
rect 10273 30714 10391 31374
rect 10273 30680 10279 30714
rect 10313 30680 10351 30714
rect 10385 30680 10391 30714
rect 10273 30641 10391 30680
rect 10273 30607 10279 30641
rect 10313 30607 10351 30641
rect 10385 30607 10391 30641
rect 10273 30568 10391 30607
rect 10273 30534 10279 30568
rect 10313 30534 10351 30568
rect 10385 30534 10391 30568
rect 10273 30495 10391 30534
rect 10273 30461 10279 30495
rect 10313 30461 10351 30495
rect 10385 30461 10391 30495
rect 10273 30422 10391 30461
rect 10273 29892 10279 30422
rect 10385 29892 10391 30422
rect 10273 29826 10279 29840
rect 10385 29826 10391 29840
rect 10273 29760 10279 29774
rect 10385 29760 10391 29774
rect 10273 29694 10279 29708
rect 10385 29694 10391 29708
rect 10273 29627 10279 29642
rect 10385 29627 10391 29642
rect 10273 29560 10279 29575
rect 10385 29560 10391 29575
rect 10273 29493 10279 29508
rect 10385 29493 10391 29508
rect 10273 29426 10279 29441
rect 10385 29426 10391 29441
rect 10325 29374 10339 29380
rect 10273 28714 10391 29374
rect 10273 28680 10279 28714
rect 10313 28680 10351 28714
rect 10385 28680 10391 28714
rect 10273 28641 10391 28680
rect 10273 28607 10279 28641
rect 10313 28607 10351 28641
rect 10385 28607 10391 28641
rect 10273 28568 10391 28607
rect 10273 28534 10279 28568
rect 10313 28534 10351 28568
rect 10385 28534 10391 28568
rect 10273 28495 10391 28534
rect 10273 28461 10279 28495
rect 10313 28461 10351 28495
rect 10385 28461 10391 28495
rect 10273 28422 10391 28461
rect 10273 27892 10279 28422
rect 10385 27892 10391 28422
rect 10273 27826 10279 27840
rect 10385 27826 10391 27840
rect 10273 27760 10279 27774
rect 10385 27760 10391 27774
rect 10273 27694 10279 27708
rect 10385 27694 10391 27708
rect 10273 27627 10279 27642
rect 10385 27627 10391 27642
rect 10273 27560 10279 27575
rect 10385 27560 10391 27575
rect 10273 27493 10279 27508
rect 10385 27493 10391 27508
rect 10273 27426 10279 27441
rect 10385 27426 10391 27441
rect 10325 27374 10339 27380
rect 10273 26785 10391 27374
rect 10273 26751 10279 26785
rect 10313 26751 10351 26785
rect 10385 26751 10391 26785
rect 10273 26707 10391 26751
rect 10273 26673 10279 26707
rect 10313 26673 10351 26707
rect 10385 26673 10391 26707
rect 10273 26629 10391 26673
rect 10273 26595 10279 26629
rect 10313 26595 10351 26629
rect 10385 26595 10391 26629
rect 10273 26551 10391 26595
rect 10273 26517 10279 26551
rect 10313 26517 10351 26551
rect 10385 26517 10391 26551
rect 10273 26473 10391 26517
rect 10273 26439 10279 26473
rect 10313 26439 10351 26473
rect 10385 26439 10391 26473
rect 10273 26396 10391 26439
rect 10273 26362 10279 26396
rect 10313 26362 10351 26396
rect 10385 26362 10391 26396
rect 10273 26319 10391 26362
rect 10273 26285 10279 26319
rect 10313 26285 10351 26319
rect 10385 26285 10391 26319
rect 10273 26242 10391 26285
rect 10273 26208 10279 26242
rect 10313 26208 10351 26242
rect 10385 26208 10391 26242
rect 10273 26165 10391 26208
rect 10273 26131 10279 26165
rect 10313 26131 10351 26165
rect 10385 26131 10391 26165
rect 10273 26088 10391 26131
rect 10273 26054 10279 26088
rect 10313 26054 10351 26088
rect 10385 26054 10391 26088
rect 10273 26011 10391 26054
rect 10273 25977 10279 26011
rect 10313 25977 10351 26011
rect 10385 25977 10391 26011
rect 10273 25934 10391 25977
rect 10273 25900 10279 25934
rect 10313 25900 10351 25934
rect 10385 25900 10391 25934
rect 10273 25891 10391 25900
rect 10325 25839 10339 25891
rect 10273 25825 10279 25839
rect 10313 25825 10351 25839
rect 10385 25825 10391 25839
rect 10325 25773 10339 25825
rect 10273 25759 10279 25773
rect 10313 25759 10351 25773
rect 10385 25759 10391 25773
rect 9437 25693 9555 25707
rect 9489 25641 9503 25693
rect 9437 25626 9555 25641
rect 9489 25574 9503 25626
rect 9437 25559 9555 25574
rect 9489 25507 9503 25559
rect 9437 25492 9555 25507
rect 9489 25440 9503 25492
rect 9437 25425 9555 25440
rect 9489 25373 9503 25425
rect 9437 25367 9555 25373
rect 10325 25707 10339 25759
rect 10691 34720 10809 34726
rect 10743 34668 10757 34720
rect 10691 34654 10809 34668
rect 10743 34602 10757 34654
rect 10691 34588 10809 34602
rect 10743 34536 10757 34588
rect 10691 34534 10697 34536
rect 10731 34534 10769 34536
rect 10803 34534 10809 34536
rect 10691 34522 10809 34534
rect 10743 34470 10757 34522
rect 10691 34461 10697 34470
rect 10731 34461 10769 34470
rect 10803 34461 10809 34470
rect 10691 34456 10809 34461
rect 10743 34422 10757 34456
rect 10691 34390 10697 34404
rect 10803 34390 10809 34404
rect 10691 34323 10697 34338
rect 10803 34323 10809 34338
rect 10691 34256 10697 34271
rect 10803 34256 10809 34271
rect 10691 33380 10697 34204
rect 10803 33380 10809 34204
rect 10691 32720 10809 33380
rect 10743 32668 10757 32720
rect 10691 32654 10809 32668
rect 10743 32602 10757 32654
rect 10691 32588 10809 32602
rect 10743 32536 10757 32588
rect 10691 32534 10697 32536
rect 10731 32534 10769 32536
rect 10803 32534 10809 32536
rect 10691 32522 10809 32534
rect 10743 32470 10757 32522
rect 10691 32461 10697 32470
rect 10731 32461 10769 32470
rect 10803 32461 10809 32470
rect 10691 32456 10809 32461
rect 10743 32422 10757 32456
rect 10691 32390 10697 32404
rect 10803 32390 10809 32404
rect 10691 32323 10697 32338
rect 10803 32323 10809 32338
rect 10691 32256 10697 32271
rect 10803 32256 10809 32271
rect 10691 31380 10697 32204
rect 10803 31380 10809 32204
rect 10691 30720 10809 31380
rect 10743 30668 10757 30720
rect 10691 30654 10809 30668
rect 10743 30602 10757 30654
rect 10691 30588 10809 30602
rect 10743 30536 10757 30588
rect 10691 30534 10697 30536
rect 10731 30534 10769 30536
rect 10803 30534 10809 30536
rect 10691 30522 10809 30534
rect 10743 30470 10757 30522
rect 10691 30461 10697 30470
rect 10731 30461 10769 30470
rect 10803 30461 10809 30470
rect 10691 30456 10809 30461
rect 10743 30422 10757 30456
rect 10691 30390 10697 30404
rect 10803 30390 10809 30404
rect 10691 30323 10697 30338
rect 10803 30323 10809 30338
rect 10691 30256 10697 30271
rect 10803 30256 10809 30271
rect 10691 29380 10697 30204
rect 10803 29380 10809 30204
rect 10691 28720 10809 29380
rect 10743 28668 10757 28720
rect 10691 28654 10809 28668
rect 10743 28602 10757 28654
rect 10691 28588 10809 28602
rect 10743 28536 10757 28588
rect 10691 28534 10697 28536
rect 10731 28534 10769 28536
rect 10803 28534 10809 28536
rect 10691 28522 10809 28534
rect 10743 28470 10757 28522
rect 10691 28461 10697 28470
rect 10731 28461 10769 28470
rect 10803 28461 10809 28470
rect 10691 28456 10809 28461
rect 10743 28422 10757 28456
rect 10691 28390 10697 28404
rect 10803 28390 10809 28404
rect 10691 28323 10697 28338
rect 10803 28323 10809 28338
rect 10691 28256 10697 28271
rect 10803 28256 10809 28271
rect 10691 27380 10697 28204
rect 10803 27380 10809 28204
rect 10691 26751 10809 27380
rect 10691 26720 10697 26751
rect 10731 26720 10769 26751
rect 10803 26720 10809 26751
rect 10743 26668 10757 26720
rect 10691 26654 10697 26668
rect 10731 26654 10769 26668
rect 10803 26654 10809 26668
rect 10743 26602 10757 26654
rect 10691 26601 10809 26602
rect 10691 26588 10697 26601
rect 10731 26588 10769 26601
rect 10803 26588 10809 26601
rect 10743 26536 10757 26588
rect 10691 26526 10809 26536
rect 10691 26522 10697 26526
rect 10731 26522 10769 26526
rect 10803 26522 10809 26526
rect 10743 26470 10757 26522
rect 10691 26456 10809 26470
rect 10743 26404 10757 26456
rect 10691 26389 10809 26404
rect 10743 26337 10757 26389
rect 10691 26322 10809 26337
rect 10743 26270 10757 26322
rect 10691 26267 10697 26270
rect 10731 26267 10769 26270
rect 10803 26267 10809 26270
rect 10691 26255 10809 26267
rect 10743 26203 10757 26255
rect 10691 26192 10697 26203
rect 10731 26192 10769 26203
rect 10803 26192 10809 26203
rect 10691 26151 10809 26192
rect 10691 26117 10697 26151
rect 10731 26117 10769 26151
rect 10803 26117 10809 26151
rect 10691 26076 10809 26117
rect 10691 26042 10697 26076
rect 10731 26042 10769 26076
rect 10803 26042 10809 26076
rect 10691 26002 10809 26042
rect 10691 25968 10697 26002
rect 10731 25968 10769 26002
rect 10803 25968 10809 26002
rect 10691 25928 10809 25968
rect 10691 25894 10697 25928
rect 10731 25894 10769 25928
rect 10803 25894 10809 25928
rect 10691 25854 10809 25894
rect 10691 25820 10697 25854
rect 10731 25820 10769 25854
rect 10803 25820 10809 25854
rect 10691 25780 10809 25820
rect 10691 25746 10697 25780
rect 10731 25746 10769 25780
rect 10803 25746 10809 25780
rect 10691 25732 10809 25746
rect 11109 34714 11227 34891
tri 11227 34821 11297 34891 nw
tri 11875 34821 11945 34891 ne
rect 11109 34680 11115 34714
rect 11149 34680 11187 34714
rect 11221 34680 11227 34714
rect 11109 34641 11227 34680
rect 11109 34607 11115 34641
rect 11149 34607 11187 34641
rect 11221 34607 11227 34641
rect 11109 34568 11227 34607
rect 11109 34534 11115 34568
rect 11149 34534 11187 34568
rect 11221 34534 11227 34568
rect 11109 34495 11227 34534
rect 11109 34461 11115 34495
rect 11149 34461 11187 34495
rect 11221 34461 11227 34495
rect 11109 34422 11227 34461
rect 11109 33892 11115 34422
rect 11221 33892 11227 34422
rect 11109 33826 11115 33840
rect 11221 33826 11227 33840
rect 11109 33760 11115 33774
rect 11221 33760 11227 33774
rect 11109 33694 11115 33708
rect 11221 33694 11227 33708
rect 11109 33627 11115 33642
rect 11221 33627 11227 33642
rect 11109 33560 11115 33575
rect 11221 33560 11227 33575
rect 11109 33493 11115 33508
rect 11221 33493 11227 33508
rect 11109 33426 11115 33441
rect 11221 33426 11227 33441
rect 11161 33374 11175 33380
rect 11109 32714 11227 33374
rect 11109 32680 11115 32714
rect 11149 32680 11187 32714
rect 11221 32680 11227 32714
rect 11109 32641 11227 32680
rect 11109 32607 11115 32641
rect 11149 32607 11187 32641
rect 11221 32607 11227 32641
rect 11109 32568 11227 32607
rect 11109 32534 11115 32568
rect 11149 32534 11187 32568
rect 11221 32534 11227 32568
rect 11109 32495 11227 32534
rect 11109 32461 11115 32495
rect 11149 32461 11187 32495
rect 11221 32461 11227 32495
rect 11109 32422 11227 32461
rect 11109 31892 11115 32422
rect 11221 31892 11227 32422
rect 11109 31826 11115 31840
rect 11221 31826 11227 31840
rect 11109 31760 11115 31774
rect 11221 31760 11227 31774
rect 11109 31694 11115 31708
rect 11221 31694 11227 31708
rect 11109 31627 11115 31642
rect 11221 31627 11227 31642
rect 11109 31560 11115 31575
rect 11221 31560 11227 31575
rect 11109 31493 11115 31508
rect 11221 31493 11227 31508
rect 11109 31426 11115 31441
rect 11221 31426 11227 31441
rect 11161 31374 11175 31380
rect 11109 30714 11227 31374
rect 11109 30680 11115 30714
rect 11149 30680 11187 30714
rect 11221 30680 11227 30714
rect 11109 30641 11227 30680
rect 11109 30607 11115 30641
rect 11149 30607 11187 30641
rect 11221 30607 11227 30641
rect 11109 30568 11227 30607
rect 11109 30534 11115 30568
rect 11149 30534 11187 30568
rect 11221 30534 11227 30568
rect 11109 30495 11227 30534
rect 11109 30461 11115 30495
rect 11149 30461 11187 30495
rect 11221 30461 11227 30495
rect 11109 30422 11227 30461
rect 11109 29892 11115 30422
rect 11221 29892 11227 30422
rect 11109 29826 11115 29840
rect 11221 29826 11227 29840
rect 11109 29760 11115 29774
rect 11221 29760 11227 29774
rect 11109 29694 11115 29708
rect 11221 29694 11227 29708
rect 11109 29627 11115 29642
rect 11221 29627 11227 29642
rect 11109 29560 11115 29575
rect 11221 29560 11227 29575
rect 11109 29493 11115 29508
rect 11221 29493 11227 29508
rect 11109 29426 11115 29441
rect 11221 29426 11227 29441
rect 11161 29374 11175 29380
rect 11109 28714 11227 29374
rect 11109 28680 11115 28714
rect 11149 28680 11187 28714
rect 11221 28680 11227 28714
rect 11109 28641 11227 28680
rect 11109 28607 11115 28641
rect 11149 28607 11187 28641
rect 11221 28607 11227 28641
rect 11109 28568 11227 28607
rect 11109 28534 11115 28568
rect 11149 28534 11187 28568
rect 11221 28534 11227 28568
rect 11109 28495 11227 28534
rect 11109 28461 11115 28495
rect 11149 28461 11187 28495
rect 11221 28461 11227 28495
rect 11109 28422 11227 28461
rect 11109 27892 11115 28422
rect 11221 27892 11227 28422
rect 11109 27826 11115 27840
rect 11221 27826 11227 27840
rect 11109 27760 11115 27774
rect 11221 27760 11227 27774
rect 11109 27694 11115 27708
rect 11221 27694 11227 27708
rect 11109 27627 11115 27642
rect 11221 27627 11227 27642
rect 11109 27560 11115 27575
rect 11221 27560 11227 27575
rect 11109 27493 11115 27508
rect 11221 27493 11227 27508
rect 11109 27426 11115 27441
rect 11221 27426 11227 27441
rect 11161 27374 11175 27380
rect 11109 26785 11227 27374
rect 11109 26751 11115 26785
rect 11149 26751 11187 26785
rect 11221 26751 11227 26785
rect 11109 26707 11227 26751
rect 11109 26673 11115 26707
rect 11149 26673 11187 26707
rect 11221 26673 11227 26707
rect 11109 26629 11227 26673
rect 11109 26595 11115 26629
rect 11149 26595 11187 26629
rect 11221 26595 11227 26629
rect 11109 26551 11227 26595
rect 11109 26517 11115 26551
rect 11149 26517 11187 26551
rect 11221 26517 11227 26551
rect 11109 26473 11227 26517
rect 11109 26439 11115 26473
rect 11149 26439 11187 26473
rect 11221 26439 11227 26473
rect 11109 26396 11227 26439
rect 11109 26362 11115 26396
rect 11149 26362 11187 26396
rect 11221 26362 11227 26396
rect 11109 26319 11227 26362
rect 11109 26285 11115 26319
rect 11149 26285 11187 26319
rect 11221 26285 11227 26319
rect 11109 26242 11227 26285
rect 11109 26208 11115 26242
rect 11149 26208 11187 26242
rect 11221 26208 11227 26242
rect 11109 26165 11227 26208
rect 11109 26131 11115 26165
rect 11149 26131 11187 26165
rect 11221 26131 11227 26165
rect 11109 26088 11227 26131
rect 11109 26054 11115 26088
rect 11149 26054 11187 26088
rect 11221 26054 11227 26088
rect 11109 26011 11227 26054
rect 11109 25977 11115 26011
rect 11149 25977 11187 26011
rect 11221 25977 11227 26011
rect 11109 25934 11227 25977
rect 11109 25900 11115 25934
rect 11149 25900 11187 25934
rect 11221 25900 11227 25934
rect 11109 25891 11227 25900
rect 11161 25839 11175 25891
rect 11109 25825 11115 25839
rect 11149 25825 11187 25839
rect 11221 25825 11227 25839
rect 11161 25773 11175 25825
rect 11109 25759 11115 25773
rect 11149 25759 11187 25773
rect 11221 25759 11227 25773
rect 10273 25693 10391 25707
rect 10325 25641 10339 25693
rect 10273 25626 10391 25641
rect 10325 25574 10339 25626
rect 10273 25559 10391 25574
rect 10325 25507 10339 25559
rect 10273 25492 10391 25507
rect 10325 25440 10339 25492
rect 10273 25425 10391 25440
rect 10325 25373 10339 25425
rect 10273 25367 10391 25373
rect 11161 25707 11175 25759
rect 11527 34720 11645 34726
rect 11579 34668 11593 34720
rect 11527 34654 11645 34668
rect 11579 34602 11593 34654
rect 11527 34588 11645 34602
rect 11579 34536 11593 34588
rect 11527 34534 11533 34536
rect 11567 34534 11605 34536
rect 11639 34534 11645 34536
rect 11527 34522 11645 34534
rect 11579 34470 11593 34522
rect 11527 34461 11533 34470
rect 11567 34461 11605 34470
rect 11639 34461 11645 34470
rect 11527 34456 11645 34461
rect 11579 34422 11593 34456
rect 11527 34390 11533 34404
rect 11639 34390 11645 34404
rect 11527 34323 11533 34338
rect 11639 34323 11645 34338
rect 11527 34256 11533 34271
rect 11639 34256 11645 34271
rect 11527 33380 11533 34204
rect 11639 33380 11645 34204
rect 11527 32720 11645 33380
rect 11579 32668 11593 32720
rect 11527 32654 11645 32668
rect 11579 32602 11593 32654
rect 11527 32588 11645 32602
rect 11579 32536 11593 32588
rect 11527 32534 11533 32536
rect 11567 32534 11605 32536
rect 11639 32534 11645 32536
rect 11527 32522 11645 32534
rect 11579 32470 11593 32522
rect 11527 32461 11533 32470
rect 11567 32461 11605 32470
rect 11639 32461 11645 32470
rect 11527 32456 11645 32461
rect 11579 32422 11593 32456
rect 11527 32390 11533 32404
rect 11639 32390 11645 32404
rect 11527 32323 11533 32338
rect 11639 32323 11645 32338
rect 11527 32256 11533 32271
rect 11639 32256 11645 32271
rect 11527 31380 11533 32204
rect 11639 31380 11645 32204
rect 11527 30720 11645 31380
rect 11579 30668 11593 30720
rect 11527 30654 11645 30668
rect 11579 30602 11593 30654
rect 11527 30588 11645 30602
rect 11579 30536 11593 30588
rect 11527 30534 11533 30536
rect 11567 30534 11605 30536
rect 11639 30534 11645 30536
rect 11527 30522 11645 30534
rect 11579 30470 11593 30522
rect 11527 30461 11533 30470
rect 11567 30461 11605 30470
rect 11639 30461 11645 30470
rect 11527 30456 11645 30461
rect 11579 30422 11593 30456
rect 11527 30390 11533 30404
rect 11639 30390 11645 30404
rect 11527 30323 11533 30338
rect 11639 30323 11645 30338
rect 11527 30256 11533 30271
rect 11639 30256 11645 30271
rect 11527 29380 11533 30204
rect 11639 29380 11645 30204
rect 11527 28720 11645 29380
rect 11579 28668 11593 28720
rect 11527 28654 11645 28668
rect 11579 28602 11593 28654
rect 11527 28588 11645 28602
rect 11579 28536 11593 28588
rect 11527 28534 11533 28536
rect 11567 28534 11605 28536
rect 11639 28534 11645 28536
rect 11527 28522 11645 28534
rect 11579 28470 11593 28522
rect 11527 28461 11533 28470
rect 11567 28461 11605 28470
rect 11639 28461 11645 28470
rect 11527 28456 11645 28461
rect 11579 28422 11593 28456
rect 11527 28390 11533 28404
rect 11639 28390 11645 28404
rect 11527 28323 11533 28338
rect 11639 28323 11645 28338
rect 11527 28256 11533 28271
rect 11639 28256 11645 28271
rect 11527 27380 11533 28204
rect 11639 27380 11645 28204
rect 11527 26751 11645 27380
rect 11527 26720 11533 26751
rect 11567 26720 11605 26751
rect 11639 26720 11645 26751
rect 11579 26668 11593 26720
rect 11527 26654 11533 26668
rect 11567 26654 11605 26668
rect 11639 26654 11645 26668
rect 11579 26602 11593 26654
rect 11527 26601 11645 26602
rect 11527 26588 11533 26601
rect 11567 26588 11605 26601
rect 11639 26588 11645 26601
rect 11579 26536 11593 26588
rect 11527 26526 11645 26536
rect 11527 26522 11533 26526
rect 11567 26522 11605 26526
rect 11639 26522 11645 26526
rect 11579 26470 11593 26522
rect 11527 26456 11645 26470
rect 11579 26404 11593 26456
rect 11527 26389 11645 26404
rect 11579 26337 11593 26389
rect 11527 26322 11645 26337
rect 11579 26270 11593 26322
rect 11527 26267 11533 26270
rect 11567 26267 11605 26270
rect 11639 26267 11645 26270
rect 11527 26255 11645 26267
rect 11579 26203 11593 26255
rect 11527 26192 11533 26203
rect 11567 26192 11605 26203
rect 11639 26192 11645 26203
rect 11527 26151 11645 26192
rect 11527 26117 11533 26151
rect 11567 26117 11605 26151
rect 11639 26117 11645 26151
rect 11527 26076 11645 26117
rect 11527 26042 11533 26076
rect 11567 26042 11605 26076
rect 11639 26042 11645 26076
rect 11527 26002 11645 26042
rect 11527 25968 11533 26002
rect 11567 25968 11605 26002
rect 11639 25968 11645 26002
rect 11527 25928 11645 25968
rect 11527 25894 11533 25928
rect 11567 25894 11605 25928
rect 11639 25894 11645 25928
rect 11527 25854 11645 25894
rect 11527 25820 11533 25854
rect 11567 25820 11605 25854
rect 11639 25820 11645 25854
rect 11527 25780 11645 25820
rect 11527 25746 11533 25780
rect 11567 25746 11605 25780
rect 11639 25746 11645 25780
rect 11527 25732 11645 25746
rect 11945 34714 12063 34891
tri 12063 34821 12133 34891 nw
tri 12711 34821 12781 34891 ne
rect 11945 34680 11951 34714
rect 11985 34680 12023 34714
rect 12057 34680 12063 34714
rect 11945 34641 12063 34680
rect 11945 34607 11951 34641
rect 11985 34607 12023 34641
rect 12057 34607 12063 34641
rect 11945 34568 12063 34607
rect 11945 34534 11951 34568
rect 11985 34534 12023 34568
rect 12057 34534 12063 34568
rect 11945 34495 12063 34534
rect 11945 34461 11951 34495
rect 11985 34461 12023 34495
rect 12057 34461 12063 34495
rect 11945 34422 12063 34461
rect 11945 33892 11951 34422
rect 12057 33892 12063 34422
rect 11945 33826 11951 33840
rect 12057 33826 12063 33840
rect 11945 33760 11951 33774
rect 12057 33760 12063 33774
rect 11945 33694 11951 33708
rect 12057 33694 12063 33708
rect 11945 33627 11951 33642
rect 12057 33627 12063 33642
rect 11945 33560 11951 33575
rect 12057 33560 12063 33575
rect 11945 33493 11951 33508
rect 12057 33493 12063 33508
rect 11945 33426 11951 33441
rect 12057 33426 12063 33441
rect 11997 33374 12011 33380
rect 11945 32714 12063 33374
rect 11945 32680 11951 32714
rect 11985 32680 12023 32714
rect 12057 32680 12063 32714
rect 11945 32641 12063 32680
rect 11945 32607 11951 32641
rect 11985 32607 12023 32641
rect 12057 32607 12063 32641
rect 11945 32568 12063 32607
rect 11945 32534 11951 32568
rect 11985 32534 12023 32568
rect 12057 32534 12063 32568
rect 11945 32495 12063 32534
rect 11945 32461 11951 32495
rect 11985 32461 12023 32495
rect 12057 32461 12063 32495
rect 11945 32422 12063 32461
rect 11945 31892 11951 32422
rect 12057 31892 12063 32422
rect 11945 31826 11951 31840
rect 12057 31826 12063 31840
rect 11945 31760 11951 31774
rect 12057 31760 12063 31774
rect 11945 31694 11951 31708
rect 12057 31694 12063 31708
rect 11945 31627 11951 31642
rect 12057 31627 12063 31642
rect 11945 31560 11951 31575
rect 12057 31560 12063 31575
rect 11945 31493 11951 31508
rect 12057 31493 12063 31508
rect 11945 31426 11951 31441
rect 12057 31426 12063 31441
rect 11997 31374 12011 31380
rect 11945 30714 12063 31374
rect 11945 30680 11951 30714
rect 11985 30680 12023 30714
rect 12057 30680 12063 30714
rect 11945 30641 12063 30680
rect 11945 30607 11951 30641
rect 11985 30607 12023 30641
rect 12057 30607 12063 30641
rect 11945 30568 12063 30607
rect 11945 30534 11951 30568
rect 11985 30534 12023 30568
rect 12057 30534 12063 30568
rect 11945 30495 12063 30534
rect 11945 30461 11951 30495
rect 11985 30461 12023 30495
rect 12057 30461 12063 30495
rect 11945 30422 12063 30461
rect 11945 29892 11951 30422
rect 12057 29892 12063 30422
rect 11945 29826 11951 29840
rect 12057 29826 12063 29840
rect 11945 29760 11951 29774
rect 12057 29760 12063 29774
rect 11945 29694 11951 29708
rect 12057 29694 12063 29708
rect 11945 29627 11951 29642
rect 12057 29627 12063 29642
rect 11945 29560 11951 29575
rect 12057 29560 12063 29575
rect 11945 29493 11951 29508
rect 12057 29493 12063 29508
rect 11945 29426 11951 29441
rect 12057 29426 12063 29441
rect 11997 29374 12011 29380
rect 11945 28714 12063 29374
rect 11945 28680 11951 28714
rect 11985 28680 12023 28714
rect 12057 28680 12063 28714
rect 11945 28641 12063 28680
rect 11945 28607 11951 28641
rect 11985 28607 12023 28641
rect 12057 28607 12063 28641
rect 11945 28568 12063 28607
rect 11945 28534 11951 28568
rect 11985 28534 12023 28568
rect 12057 28534 12063 28568
rect 11945 28495 12063 28534
rect 11945 28461 11951 28495
rect 11985 28461 12023 28495
rect 12057 28461 12063 28495
rect 11945 28422 12063 28461
rect 11945 27892 11951 28422
rect 12057 27892 12063 28422
rect 11945 27826 11951 27840
rect 12057 27826 12063 27840
rect 11945 27760 11951 27774
rect 12057 27760 12063 27774
rect 11945 27694 11951 27708
rect 12057 27694 12063 27708
rect 11945 27627 11951 27642
rect 12057 27627 12063 27642
rect 11945 27560 11951 27575
rect 12057 27560 12063 27575
rect 11945 27493 11951 27508
rect 12057 27493 12063 27508
rect 11945 27426 11951 27441
rect 12057 27426 12063 27441
rect 11997 27374 12011 27380
rect 11945 26785 12063 27374
rect 11945 26751 11951 26785
rect 11985 26751 12023 26785
rect 12057 26751 12063 26785
rect 11945 26707 12063 26751
rect 11945 26673 11951 26707
rect 11985 26673 12023 26707
rect 12057 26673 12063 26707
rect 11945 26629 12063 26673
rect 11945 26595 11951 26629
rect 11985 26595 12023 26629
rect 12057 26595 12063 26629
rect 11945 26551 12063 26595
rect 11945 26517 11951 26551
rect 11985 26517 12023 26551
rect 12057 26517 12063 26551
rect 11945 26473 12063 26517
rect 11945 26439 11951 26473
rect 11985 26439 12023 26473
rect 12057 26439 12063 26473
rect 11945 26396 12063 26439
rect 11945 26362 11951 26396
rect 11985 26362 12023 26396
rect 12057 26362 12063 26396
rect 11945 26319 12063 26362
rect 11945 26285 11951 26319
rect 11985 26285 12023 26319
rect 12057 26285 12063 26319
rect 11945 26242 12063 26285
rect 11945 26208 11951 26242
rect 11985 26208 12023 26242
rect 12057 26208 12063 26242
rect 11945 26165 12063 26208
rect 11945 26131 11951 26165
rect 11985 26131 12023 26165
rect 12057 26131 12063 26165
rect 11945 26088 12063 26131
rect 11945 26054 11951 26088
rect 11985 26054 12023 26088
rect 12057 26054 12063 26088
rect 11945 26011 12063 26054
rect 11945 25977 11951 26011
rect 11985 25977 12023 26011
rect 12057 25977 12063 26011
rect 11945 25934 12063 25977
rect 11945 25900 11951 25934
rect 11985 25900 12023 25934
rect 12057 25900 12063 25934
rect 11945 25891 12063 25900
rect 11997 25839 12011 25891
rect 11945 25825 11951 25839
rect 11985 25825 12023 25839
rect 12057 25825 12063 25839
rect 11997 25773 12011 25825
rect 11945 25759 11951 25773
rect 11985 25759 12023 25773
rect 12057 25759 12063 25773
rect 11109 25693 11227 25707
rect 11161 25641 11175 25693
rect 11109 25626 11227 25641
rect 11161 25574 11175 25626
rect 11109 25559 11227 25574
rect 11161 25507 11175 25559
rect 11109 25492 11227 25507
rect 11161 25440 11175 25492
rect 11109 25425 11227 25440
rect 11161 25373 11175 25425
rect 11109 25367 11227 25373
rect 11997 25707 12011 25759
rect 12363 34720 12481 34726
rect 12415 34668 12429 34720
rect 12363 34654 12481 34668
rect 12415 34602 12429 34654
rect 12363 34588 12481 34602
rect 12415 34536 12429 34588
rect 12363 34534 12369 34536
rect 12403 34534 12441 34536
rect 12475 34534 12481 34536
rect 12363 34522 12481 34534
rect 12415 34470 12429 34522
rect 12363 34461 12369 34470
rect 12403 34461 12441 34470
rect 12475 34461 12481 34470
rect 12363 34456 12481 34461
rect 12415 34422 12429 34456
rect 12363 34390 12369 34404
rect 12475 34390 12481 34404
rect 12363 34323 12369 34338
rect 12475 34323 12481 34338
rect 12363 34256 12369 34271
rect 12475 34256 12481 34271
rect 12363 33380 12369 34204
rect 12475 33380 12481 34204
rect 12363 32720 12481 33380
rect 12415 32668 12429 32720
rect 12363 32654 12481 32668
rect 12415 32602 12429 32654
rect 12363 32588 12481 32602
rect 12415 32536 12429 32588
rect 12363 32534 12369 32536
rect 12403 32534 12441 32536
rect 12475 32534 12481 32536
rect 12363 32522 12481 32534
rect 12415 32470 12429 32522
rect 12363 32461 12369 32470
rect 12403 32461 12441 32470
rect 12475 32461 12481 32470
rect 12363 32456 12481 32461
rect 12415 32422 12429 32456
rect 12363 32390 12369 32404
rect 12475 32390 12481 32404
rect 12363 32323 12369 32338
rect 12475 32323 12481 32338
rect 12363 32256 12369 32271
rect 12475 32256 12481 32271
rect 12363 31380 12369 32204
rect 12475 31380 12481 32204
rect 12363 30720 12481 31380
rect 12415 30668 12429 30720
rect 12363 30654 12481 30668
rect 12415 30602 12429 30654
rect 12363 30588 12481 30602
rect 12415 30536 12429 30588
rect 12363 30534 12369 30536
rect 12403 30534 12441 30536
rect 12475 30534 12481 30536
rect 12363 30522 12481 30534
rect 12415 30470 12429 30522
rect 12363 30461 12369 30470
rect 12403 30461 12441 30470
rect 12475 30461 12481 30470
rect 12363 30456 12481 30461
rect 12415 30422 12429 30456
rect 12363 30390 12369 30404
rect 12475 30390 12481 30404
rect 12363 30323 12369 30338
rect 12475 30323 12481 30338
rect 12363 30256 12369 30271
rect 12475 30256 12481 30271
rect 12363 29380 12369 30204
rect 12475 29380 12481 30204
rect 12363 28720 12481 29380
rect 12415 28668 12429 28720
rect 12363 28654 12481 28668
rect 12415 28602 12429 28654
rect 12363 28588 12481 28602
rect 12415 28536 12429 28588
rect 12363 28534 12369 28536
rect 12403 28534 12441 28536
rect 12475 28534 12481 28536
rect 12363 28522 12481 28534
rect 12415 28470 12429 28522
rect 12363 28461 12369 28470
rect 12403 28461 12441 28470
rect 12475 28461 12481 28470
rect 12363 28456 12481 28461
rect 12415 28422 12429 28456
rect 12363 28390 12369 28404
rect 12475 28390 12481 28404
rect 12363 28323 12369 28338
rect 12475 28323 12481 28338
rect 12363 28256 12369 28271
rect 12475 28256 12481 28271
rect 12363 27380 12369 28204
rect 12475 27380 12481 28204
rect 12363 26751 12481 27380
rect 12363 26720 12369 26751
rect 12403 26720 12441 26751
rect 12475 26720 12481 26751
rect 12415 26668 12429 26720
rect 12363 26654 12369 26668
rect 12403 26654 12441 26668
rect 12475 26654 12481 26668
rect 12415 26602 12429 26654
rect 12363 26601 12481 26602
rect 12363 26588 12369 26601
rect 12403 26588 12441 26601
rect 12475 26588 12481 26601
rect 12415 26536 12429 26588
rect 12363 26526 12481 26536
rect 12363 26522 12369 26526
rect 12403 26522 12441 26526
rect 12475 26522 12481 26526
rect 12415 26470 12429 26522
rect 12363 26456 12481 26470
rect 12415 26404 12429 26456
rect 12363 26389 12481 26404
rect 12415 26337 12429 26389
rect 12363 26322 12481 26337
rect 12415 26270 12429 26322
rect 12363 26267 12369 26270
rect 12403 26267 12441 26270
rect 12475 26267 12481 26270
rect 12363 26255 12481 26267
rect 12415 26203 12429 26255
rect 12363 26192 12369 26203
rect 12403 26192 12441 26203
rect 12475 26192 12481 26203
rect 12363 26151 12481 26192
rect 12363 26117 12369 26151
rect 12403 26117 12441 26151
rect 12475 26117 12481 26151
rect 12363 26076 12481 26117
rect 12363 26042 12369 26076
rect 12403 26042 12441 26076
rect 12475 26042 12481 26076
rect 12363 26002 12481 26042
rect 12363 25968 12369 26002
rect 12403 25968 12441 26002
rect 12475 25968 12481 26002
rect 12363 25928 12481 25968
rect 12363 25894 12369 25928
rect 12403 25894 12441 25928
rect 12475 25894 12481 25928
rect 12363 25854 12481 25894
rect 12363 25820 12369 25854
rect 12403 25820 12441 25854
rect 12475 25820 12481 25854
rect 12363 25780 12481 25820
rect 12363 25746 12369 25780
rect 12403 25746 12441 25780
rect 12475 25746 12481 25780
rect 12363 25732 12481 25746
rect 12781 34714 12899 34891
tri 12899 34821 12969 34891 nw
rect 12781 34680 12787 34714
rect 12821 34680 12859 34714
rect 12893 34680 12899 34714
rect 12781 34641 12899 34680
rect 12781 34607 12787 34641
rect 12821 34607 12859 34641
rect 12893 34607 12899 34641
rect 12781 34568 12899 34607
rect 12781 34534 12787 34568
rect 12821 34534 12859 34568
rect 12893 34534 12899 34568
rect 12781 34495 12899 34534
rect 12781 34461 12787 34495
rect 12821 34461 12859 34495
rect 12893 34461 12899 34495
rect 12781 34422 12899 34461
rect 12781 33892 12787 34422
rect 12893 33892 12899 34422
rect 12781 33826 12787 33840
rect 12893 33826 12899 33840
rect 12781 33760 12787 33774
rect 12893 33760 12899 33774
rect 12781 33694 12787 33708
rect 12893 33694 12899 33708
rect 12781 33627 12787 33642
rect 12893 33627 12899 33642
rect 12781 33560 12787 33575
rect 12893 33560 12899 33575
rect 12781 33493 12787 33508
rect 12893 33493 12899 33508
rect 12781 33426 12787 33441
rect 12893 33426 12899 33441
rect 12833 33374 12847 33380
rect 12781 32714 12899 33374
rect 12781 32680 12787 32714
rect 12821 32680 12859 32714
rect 12893 32680 12899 32714
rect 12781 32641 12899 32680
rect 12781 32607 12787 32641
rect 12821 32607 12859 32641
rect 12893 32607 12899 32641
rect 12781 32568 12899 32607
rect 12781 32534 12787 32568
rect 12821 32534 12859 32568
rect 12893 32534 12899 32568
rect 12781 32495 12899 32534
rect 12781 32461 12787 32495
rect 12821 32461 12859 32495
rect 12893 32461 12899 32495
rect 12781 32422 12899 32461
rect 12781 31892 12787 32422
rect 12893 31892 12899 32422
rect 12781 31826 12787 31840
rect 12893 31826 12899 31840
rect 12781 31760 12787 31774
rect 12893 31760 12899 31774
rect 12781 31694 12787 31708
rect 12893 31694 12899 31708
rect 12781 31627 12787 31642
rect 12893 31627 12899 31642
rect 12781 31560 12787 31575
rect 12893 31560 12899 31575
rect 12781 31493 12787 31508
rect 12893 31493 12899 31508
rect 12781 31426 12787 31441
rect 12893 31426 12899 31441
rect 12833 31374 12847 31380
rect 12781 30714 12899 31374
rect 12781 30680 12787 30714
rect 12821 30680 12859 30714
rect 12893 30680 12899 30714
rect 12781 30641 12899 30680
rect 12781 30607 12787 30641
rect 12821 30607 12859 30641
rect 12893 30607 12899 30641
rect 12781 30568 12899 30607
rect 12781 30534 12787 30568
rect 12821 30534 12859 30568
rect 12893 30534 12899 30568
rect 12781 30495 12899 30534
rect 12781 30461 12787 30495
rect 12821 30461 12859 30495
rect 12893 30461 12899 30495
rect 12781 30422 12899 30461
rect 12781 29892 12787 30422
rect 12893 29892 12899 30422
rect 12781 29826 12787 29840
rect 12893 29826 12899 29840
rect 12781 29760 12787 29774
rect 12893 29760 12899 29774
rect 12781 29694 12787 29708
rect 12893 29694 12899 29708
rect 12781 29627 12787 29642
rect 12893 29627 12899 29642
rect 12781 29560 12787 29575
rect 12893 29560 12899 29575
rect 12781 29493 12787 29508
rect 12893 29493 12899 29508
rect 12781 29426 12787 29441
rect 12893 29426 12899 29441
rect 12833 29374 12847 29380
rect 12781 28714 12899 29374
rect 12781 28680 12787 28714
rect 12821 28680 12859 28714
rect 12893 28680 12899 28714
rect 12781 28641 12899 28680
rect 12781 28607 12787 28641
rect 12821 28607 12859 28641
rect 12893 28607 12899 28641
rect 12781 28568 12899 28607
rect 12781 28534 12787 28568
rect 12821 28534 12859 28568
rect 12893 28534 12899 28568
rect 12781 28495 12899 28534
rect 12781 28461 12787 28495
rect 12821 28461 12859 28495
rect 12893 28461 12899 28495
rect 12781 28422 12899 28461
rect 12781 27892 12787 28422
rect 12893 27892 12899 28422
rect 12781 27826 12787 27840
rect 12893 27826 12899 27840
rect 12781 27760 12787 27774
rect 12893 27760 12899 27774
rect 12781 27694 12787 27708
rect 12893 27694 12899 27708
rect 12781 27627 12787 27642
rect 12893 27627 12899 27642
rect 12781 27560 12787 27575
rect 12893 27560 12899 27575
rect 12781 27493 12787 27508
rect 12893 27493 12899 27508
rect 12781 27426 12787 27441
rect 12893 27426 12899 27441
rect 12833 27374 12847 27380
rect 12781 26785 12899 27374
rect 12781 26751 12787 26785
rect 12821 26751 12859 26785
rect 12893 26751 12899 26785
rect 12781 26707 12899 26751
rect 12781 26673 12787 26707
rect 12821 26673 12859 26707
rect 12893 26673 12899 26707
rect 12781 26629 12899 26673
rect 12781 26595 12787 26629
rect 12821 26595 12859 26629
rect 12893 26595 12899 26629
rect 12781 26551 12899 26595
rect 12781 26517 12787 26551
rect 12821 26517 12859 26551
rect 12893 26517 12899 26551
rect 12781 26473 12899 26517
rect 12781 26439 12787 26473
rect 12821 26439 12859 26473
rect 12893 26439 12899 26473
rect 12781 26396 12899 26439
rect 12781 26362 12787 26396
rect 12821 26362 12859 26396
rect 12893 26362 12899 26396
rect 12781 26319 12899 26362
rect 12781 26285 12787 26319
rect 12821 26285 12859 26319
rect 12893 26285 12899 26319
rect 12781 26242 12899 26285
rect 12781 26208 12787 26242
rect 12821 26208 12859 26242
rect 12893 26208 12899 26242
rect 12781 26165 12899 26208
rect 12781 26131 12787 26165
rect 12821 26131 12859 26165
rect 12893 26131 12899 26165
rect 12781 26088 12899 26131
rect 12781 26054 12787 26088
rect 12821 26054 12859 26088
rect 12893 26054 12899 26088
rect 12781 26011 12899 26054
rect 12781 25977 12787 26011
rect 12821 25977 12859 26011
rect 12893 25977 12899 26011
rect 12781 25934 12899 25977
rect 12781 25900 12787 25934
rect 12821 25900 12859 25934
rect 12893 25900 12899 25934
rect 12781 25891 12899 25900
rect 12833 25839 12847 25891
rect 12781 25825 12787 25839
rect 12821 25825 12859 25839
rect 12893 25825 12899 25839
rect 12833 25773 12847 25825
rect 12781 25759 12787 25773
rect 12821 25759 12859 25773
rect 12893 25759 12899 25773
rect 11945 25693 12063 25707
rect 11997 25641 12011 25693
rect 11945 25626 12063 25641
rect 11997 25574 12011 25626
rect 11945 25559 12063 25574
rect 11997 25507 12011 25559
rect 11945 25492 12063 25507
rect 11997 25440 12011 25492
rect 11945 25425 12063 25440
rect 11997 25373 12011 25425
rect 11945 25367 12063 25373
rect 12833 25707 12847 25759
rect 12781 25693 12899 25707
rect 12833 25641 12847 25693
rect 12781 25626 12899 25641
rect 12833 25574 12847 25626
rect 12781 25559 12899 25574
rect 12833 25507 12847 25559
rect 12781 25492 12899 25507
rect 12833 25440 12847 25492
rect 12781 25425 12899 25440
rect 12833 25373 12847 25425
rect 12781 25367 12899 25373
rect 13199 34720 13521 35380
rect 13199 34668 13200 34720
rect 13252 34668 13270 34720
rect 13322 34668 13340 34720
rect 13392 34668 13410 34720
rect 13462 34668 13480 34720
rect 13199 34654 13521 34668
rect 13199 34602 13200 34654
rect 13252 34602 13270 34654
rect 13322 34602 13340 34654
rect 13392 34602 13410 34654
rect 13462 34602 13480 34654
rect 13199 34588 13521 34602
rect 13199 34536 13200 34588
rect 13252 34536 13270 34588
rect 13322 34536 13340 34588
rect 13392 34536 13410 34588
rect 13462 34536 13480 34588
rect 13199 34534 13205 34536
rect 13239 34534 13277 34536
rect 13311 34534 13521 34536
rect 13199 34522 13521 34534
rect 13199 34470 13200 34522
rect 13252 34470 13270 34522
rect 13322 34470 13340 34522
rect 13392 34470 13410 34522
rect 13462 34470 13480 34522
rect 13199 34461 13205 34470
rect 13239 34461 13277 34470
rect 13311 34461 13521 34470
rect 13199 34456 13521 34461
rect 13199 34404 13200 34456
rect 13252 34422 13270 34456
rect 13322 34404 13340 34456
rect 13392 34404 13410 34456
rect 13462 34404 13480 34456
rect 13199 34390 13205 34404
rect 13311 34390 13521 34404
rect 13199 34338 13200 34390
rect 13322 34338 13340 34390
rect 13392 34338 13410 34390
rect 13462 34338 13480 34390
rect 13199 34323 13205 34338
rect 13311 34323 13521 34338
rect 13199 34271 13200 34323
rect 13322 34271 13340 34323
rect 13392 34271 13410 34323
rect 13462 34271 13480 34323
rect 13199 34256 13205 34271
rect 13311 34256 13521 34271
rect 13199 34204 13200 34256
rect 13322 34204 13340 34256
rect 13392 34204 13410 34256
rect 13462 34204 13480 34256
rect 13199 33380 13205 34204
rect 13311 33380 13521 34204
rect 13199 32720 13521 33380
rect 13199 32668 13200 32720
rect 13252 32668 13270 32720
rect 13322 32668 13340 32720
rect 13392 32668 13410 32720
rect 13462 32668 13480 32720
rect 13199 32654 13521 32668
rect 13199 32602 13200 32654
rect 13252 32602 13270 32654
rect 13322 32602 13340 32654
rect 13392 32602 13410 32654
rect 13462 32602 13480 32654
rect 13199 32588 13521 32602
rect 13199 32536 13200 32588
rect 13252 32536 13270 32588
rect 13322 32536 13340 32588
rect 13392 32536 13410 32588
rect 13462 32536 13480 32588
rect 13199 32534 13205 32536
rect 13239 32534 13277 32536
rect 13311 32534 13521 32536
rect 13199 32522 13521 32534
rect 13199 32470 13200 32522
rect 13252 32470 13270 32522
rect 13322 32470 13340 32522
rect 13392 32470 13410 32522
rect 13462 32470 13480 32522
rect 13199 32461 13205 32470
rect 13239 32461 13277 32470
rect 13311 32461 13521 32470
rect 13199 32456 13521 32461
rect 13199 32404 13200 32456
rect 13252 32422 13270 32456
rect 13322 32404 13340 32456
rect 13392 32404 13410 32456
rect 13462 32404 13480 32456
rect 13199 32390 13205 32404
rect 13311 32390 13521 32404
rect 13199 32338 13200 32390
rect 13322 32338 13340 32390
rect 13392 32338 13410 32390
rect 13462 32338 13480 32390
rect 13199 32323 13205 32338
rect 13311 32323 13521 32338
rect 13199 32271 13200 32323
rect 13322 32271 13340 32323
rect 13392 32271 13410 32323
rect 13462 32271 13480 32323
rect 13199 32256 13205 32271
rect 13311 32256 13521 32271
rect 13199 32204 13200 32256
rect 13322 32204 13340 32256
rect 13392 32204 13410 32256
rect 13462 32204 13480 32256
rect 13199 31380 13205 32204
rect 13311 31380 13521 32204
rect 13199 30720 13521 31380
rect 13199 30668 13200 30720
rect 13252 30668 13270 30720
rect 13322 30668 13340 30720
rect 13392 30668 13410 30720
rect 13462 30668 13480 30720
rect 13199 30654 13521 30668
rect 13199 30602 13200 30654
rect 13252 30602 13270 30654
rect 13322 30602 13340 30654
rect 13392 30602 13410 30654
rect 13462 30602 13480 30654
rect 13199 30588 13521 30602
rect 13199 30536 13200 30588
rect 13252 30536 13270 30588
rect 13322 30536 13340 30588
rect 13392 30536 13410 30588
rect 13462 30536 13480 30588
rect 13199 30534 13205 30536
rect 13239 30534 13277 30536
rect 13311 30534 13521 30536
rect 13199 30522 13521 30534
rect 13199 30470 13200 30522
rect 13252 30470 13270 30522
rect 13322 30470 13340 30522
rect 13392 30470 13410 30522
rect 13462 30470 13480 30522
rect 13199 30461 13205 30470
rect 13239 30461 13277 30470
rect 13311 30461 13521 30470
rect 13199 30456 13521 30461
rect 13199 30404 13200 30456
rect 13252 30422 13270 30456
rect 13322 30404 13340 30456
rect 13392 30404 13410 30456
rect 13462 30404 13480 30456
rect 13199 30390 13205 30404
rect 13311 30390 13521 30404
rect 13199 30338 13200 30390
rect 13322 30338 13340 30390
rect 13392 30338 13410 30390
rect 13462 30338 13480 30390
rect 13199 30323 13205 30338
rect 13311 30323 13521 30338
rect 13199 30271 13200 30323
rect 13322 30271 13340 30323
rect 13392 30271 13410 30323
rect 13462 30271 13480 30323
rect 13199 30256 13205 30271
rect 13311 30256 13521 30271
rect 13199 30204 13200 30256
rect 13322 30204 13340 30256
rect 13392 30204 13410 30256
rect 13462 30204 13480 30256
rect 13199 29380 13205 30204
rect 13311 29380 13521 30204
rect 13199 28720 13521 29380
rect 13199 28668 13200 28720
rect 13252 28668 13270 28720
rect 13322 28668 13340 28720
rect 13392 28668 13410 28720
rect 13462 28668 13480 28720
rect 13199 28654 13521 28668
rect 13199 28602 13200 28654
rect 13252 28602 13270 28654
rect 13322 28602 13340 28654
rect 13392 28602 13410 28654
rect 13462 28602 13480 28654
rect 13199 28588 13521 28602
rect 13199 28536 13200 28588
rect 13252 28536 13270 28588
rect 13322 28536 13340 28588
rect 13392 28536 13410 28588
rect 13462 28536 13480 28588
rect 13199 28534 13205 28536
rect 13239 28534 13277 28536
rect 13311 28534 13521 28536
rect 13199 28522 13521 28534
rect 13199 28470 13200 28522
rect 13252 28470 13270 28522
rect 13322 28470 13340 28522
rect 13392 28470 13410 28522
rect 13462 28470 13480 28522
rect 13199 28461 13205 28470
rect 13239 28461 13277 28470
rect 13311 28461 13521 28470
rect 13199 28456 13521 28461
rect 13199 28404 13200 28456
rect 13252 28422 13270 28456
rect 13322 28404 13340 28456
rect 13392 28404 13410 28456
rect 13462 28404 13480 28456
rect 13199 28390 13205 28404
rect 13311 28390 13521 28404
rect 13199 28338 13200 28390
rect 13322 28338 13340 28390
rect 13392 28338 13410 28390
rect 13462 28338 13480 28390
rect 13199 28323 13205 28338
rect 13311 28323 13521 28338
rect 13199 28271 13200 28323
rect 13322 28271 13340 28323
rect 13392 28271 13410 28323
rect 13462 28271 13480 28323
rect 13199 28256 13205 28271
rect 13311 28256 13521 28271
rect 13199 28204 13200 28256
rect 13322 28204 13340 28256
rect 13392 28204 13410 28256
rect 13462 28204 13480 28256
rect 13199 27380 13205 28204
rect 13311 27380 13521 28204
rect 13199 26751 13521 27380
rect 13199 26720 13205 26751
rect 13239 26720 13277 26751
rect 13311 26720 13521 26751
rect 13199 26668 13200 26720
rect 13252 26668 13270 26720
rect 13322 26668 13340 26720
rect 13392 26668 13410 26720
rect 13462 26668 13480 26720
rect 13199 26654 13205 26668
rect 13239 26654 13277 26668
rect 13311 26654 13521 26668
rect 13199 26602 13200 26654
rect 13252 26602 13270 26654
rect 13322 26602 13340 26654
rect 13392 26602 13410 26654
rect 13462 26602 13480 26654
rect 13199 26601 13521 26602
rect 13199 26588 13205 26601
rect 13239 26588 13277 26601
rect 13311 26588 13521 26601
rect 13199 26536 13200 26588
rect 13252 26536 13270 26588
rect 13322 26536 13340 26588
rect 13392 26536 13410 26588
rect 13462 26536 13480 26588
rect 13199 26526 13521 26536
rect 13199 26522 13205 26526
rect 13239 26522 13277 26526
rect 13311 26522 13521 26526
rect 13199 26470 13200 26522
rect 13252 26470 13270 26522
rect 13322 26470 13340 26522
rect 13392 26470 13410 26522
rect 13462 26470 13480 26522
rect 13199 26456 13521 26470
rect 13199 26404 13200 26456
rect 13252 26404 13270 26456
rect 13322 26404 13340 26456
rect 13392 26404 13410 26456
rect 13462 26404 13480 26456
rect 13199 26389 13521 26404
rect 13199 26337 13200 26389
rect 13252 26337 13270 26389
rect 13322 26337 13340 26389
rect 13392 26337 13410 26389
rect 13462 26337 13480 26389
rect 13199 26322 13521 26337
rect 13199 26270 13200 26322
rect 13252 26270 13270 26322
rect 13322 26270 13340 26322
rect 13392 26270 13410 26322
rect 13462 26270 13480 26322
rect 13199 26267 13205 26270
rect 13239 26267 13277 26270
rect 13311 26267 13521 26270
rect 13199 26255 13521 26267
rect 13199 26203 13200 26255
rect 13252 26203 13270 26255
rect 13322 26203 13340 26255
rect 13392 26203 13410 26255
rect 13462 26203 13480 26255
rect 13199 26192 13205 26203
rect 13239 26192 13277 26203
rect 13311 26192 13521 26203
rect 13199 26151 13521 26192
rect 13199 26117 13205 26151
rect 13239 26117 13277 26151
rect 13311 26117 13521 26151
rect 13199 26076 13521 26117
rect 13199 26042 13205 26076
rect 13239 26042 13277 26076
rect 13311 26042 13521 26076
rect 13199 26002 13521 26042
rect 13199 25968 13205 26002
rect 13239 25968 13277 26002
rect 13311 25968 13521 26002
rect 13199 25928 13521 25968
rect 13199 25894 13205 25928
rect 13239 25894 13277 25928
rect 13311 25894 13521 25928
rect 13199 25854 13521 25894
rect 13199 25820 13205 25854
rect 13239 25820 13277 25854
rect 13311 25820 13521 25854
rect 13199 25780 13521 25820
rect 13199 25746 13205 25780
rect 13239 25746 13277 25780
rect 13311 25746 13521 25780
tri 4532 25071 4678 25217 sw
tri 13129 25071 13199 25141 se
rect 13199 25071 13521 25746
rect 4332 25059 4767 25071
rect 4332 25025 4727 25059
rect 4761 25025 4767 25059
rect 4332 24986 4767 25025
rect 4332 24952 4727 24986
rect 4761 24952 4767 24986
tri 13042 24984 13129 25071 se
rect 13129 24984 13521 25071
rect 4332 24914 4767 24952
rect 4332 24880 4727 24914
rect 4761 24880 4767 24914
rect 4332 24842 4767 24880
rect 4332 24808 4727 24842
rect 4761 24808 4767 24842
rect 4332 24770 4767 24808
rect 4332 24736 4727 24770
rect 4761 24736 4767 24770
rect 4332 24698 4767 24736
rect 4332 24664 4727 24698
rect 4761 24664 4767 24698
rect 4332 24626 4767 24664
rect 4332 24592 4727 24626
rect 4761 24592 4767 24626
rect 4332 24554 4767 24592
rect 4332 24520 4727 24554
rect 4761 24520 4767 24554
rect 4332 24482 4767 24520
rect 4332 24448 4727 24482
rect 4761 24448 4767 24482
rect 4332 24410 4767 24448
rect 4332 24376 4727 24410
rect 4761 24376 4767 24410
rect 4332 24338 4767 24376
rect 4332 24304 4727 24338
rect 4761 24304 4767 24338
rect 4332 24266 4767 24304
rect 4332 24232 4727 24266
rect 4761 24232 4767 24266
rect 4332 24194 4767 24232
rect 4332 24160 4727 24194
rect 4761 24160 4767 24194
rect 4332 24122 4767 24160
rect 4332 24088 4727 24122
rect 4761 24088 4767 24122
rect 4332 24050 4767 24088
rect 4332 24016 4727 24050
rect 4761 24016 4767 24050
rect 4332 23110 4767 24016
rect 5067 24972 13521 24984
rect 5067 24938 5073 24972
rect 5107 24938 6719 24972
rect 6753 24938 8374 24972
rect 8408 24938 10030 24972
rect 10064 24938 11686 24972
rect 11720 24938 13342 24972
rect 13376 24938 13521 24972
rect 5067 24895 13521 24938
rect 5067 24861 5073 24895
rect 5107 24861 6719 24895
rect 6753 24861 8374 24895
rect 8408 24861 10030 24895
rect 10064 24861 11686 24895
rect 11720 24861 13342 24895
rect 13376 24861 13521 24895
rect 5067 24818 13521 24861
rect 5067 24784 5073 24818
rect 5107 24784 6719 24818
rect 6753 24784 8374 24818
rect 8408 24784 10030 24818
rect 10064 24784 11686 24818
rect 11720 24784 13342 24818
rect 13376 24784 13521 24818
rect 5067 24741 13521 24784
rect 5067 24707 5073 24741
rect 5107 24707 6719 24741
rect 6753 24707 8374 24741
rect 8408 24707 10030 24741
rect 10064 24707 11686 24741
rect 11720 24707 13342 24741
rect 13376 24707 13521 24741
rect 5067 24664 13521 24707
rect 5067 24630 5073 24664
rect 5107 24630 6719 24664
rect 6753 24630 8374 24664
rect 8408 24630 10030 24664
rect 10064 24630 11686 24664
rect 11720 24630 13342 24664
rect 13376 24630 13521 24664
rect 5067 24587 13521 24630
rect 5067 24553 5073 24587
rect 5107 24553 6719 24587
rect 6753 24553 8374 24587
rect 8408 24553 10030 24587
rect 10064 24553 11686 24587
rect 11720 24553 13342 24587
rect 13376 24553 13521 24587
rect 5067 24510 13521 24553
rect 5067 24476 5073 24510
rect 5107 24476 6719 24510
rect 6753 24476 8374 24510
rect 8408 24476 10030 24510
rect 10064 24476 11686 24510
rect 11720 24476 13342 24510
rect 13376 24476 13521 24510
rect 5067 24433 13521 24476
rect 5067 24399 5073 24433
rect 5107 24399 6719 24433
rect 6753 24399 8374 24433
rect 8408 24399 10030 24433
rect 10064 24399 11686 24433
rect 11720 24399 13342 24433
rect 13376 24399 13521 24433
rect 5067 24356 13521 24399
rect 5067 24322 5073 24356
rect 5107 24322 6719 24356
rect 6753 24322 8374 24356
rect 8408 24322 10030 24356
rect 10064 24322 11686 24356
rect 11720 24322 13342 24356
rect 13376 24322 13521 24356
rect 5067 24279 13521 24322
rect 5067 24245 5073 24279
rect 5107 24245 6719 24279
rect 6753 24245 8374 24279
rect 8408 24245 10030 24279
rect 10064 24245 11686 24279
rect 11720 24245 13342 24279
rect 13376 24245 13521 24279
rect 5067 24202 13521 24245
rect 5067 24168 5073 24202
rect 5107 24168 6719 24202
rect 6753 24168 8374 24202
rect 8408 24168 10030 24202
rect 10064 24168 11686 24202
rect 11720 24168 13342 24202
rect 13376 24168 13521 24202
rect 5067 24126 13521 24168
rect 5067 24092 5073 24126
rect 5107 24092 6719 24126
rect 6753 24092 8374 24126
rect 8408 24092 10030 24126
rect 10064 24092 11686 24126
rect 11720 24092 13342 24126
rect 13376 24092 13521 24126
rect 5067 24050 13521 24092
rect 5067 24016 5073 24050
rect 5107 24016 6719 24050
rect 6753 24016 8374 24050
rect 8408 24016 10030 24050
rect 10064 24016 11686 24050
rect 11720 24016 13342 24050
rect 13376 24016 13521 24050
rect 5067 24004 13521 24016
tri 13358 23847 13515 24004 ne
rect 5069 23651 5075 23703
rect 5127 23651 5151 23703
rect 5203 23651 5226 23703
rect 5278 23697 5301 23703
rect 5353 23697 5376 23703
rect 5428 23697 5451 23703
rect 5503 23697 13343 23703
rect 5278 23663 5300 23697
rect 5353 23663 5373 23697
rect 5428 23663 5446 23697
rect 5503 23663 5519 23697
rect 5553 23663 5592 23697
rect 5626 23663 5665 23697
rect 5699 23663 5737 23697
rect 5771 23663 5809 23697
rect 5843 23663 5881 23697
rect 5915 23663 5953 23697
rect 5987 23663 6025 23697
rect 6059 23663 6097 23697
rect 6131 23663 6169 23697
rect 6203 23663 6241 23697
rect 6275 23663 6313 23697
rect 6347 23663 6385 23697
rect 6419 23663 6457 23697
rect 6491 23663 6529 23697
rect 6563 23663 6601 23697
rect 6635 23663 6673 23697
rect 6707 23663 6745 23697
rect 6779 23663 6817 23697
rect 6851 23663 6889 23697
rect 6923 23663 6961 23697
rect 6995 23663 7033 23697
rect 7067 23663 7105 23697
rect 7139 23663 7177 23697
rect 7211 23663 7249 23697
rect 7283 23663 7321 23697
rect 7355 23663 7393 23697
rect 7427 23663 7465 23697
rect 7499 23663 7537 23697
rect 7571 23663 7609 23697
rect 7643 23663 7681 23697
rect 7715 23663 7753 23697
rect 7787 23663 7825 23697
rect 7859 23663 7897 23697
rect 7931 23663 7969 23697
rect 8003 23663 8041 23697
rect 8075 23663 8113 23697
rect 8147 23663 8185 23697
rect 8219 23663 8257 23697
rect 8291 23663 8329 23697
rect 8363 23663 8401 23697
rect 8435 23663 8473 23697
rect 8507 23663 8545 23697
rect 8579 23663 8617 23697
rect 8651 23663 8689 23697
rect 8723 23663 8761 23697
rect 8795 23663 8833 23697
rect 8867 23663 8905 23697
rect 8939 23663 8977 23697
rect 9011 23663 9049 23697
rect 9083 23663 9121 23697
rect 9155 23663 9193 23697
rect 9227 23663 9265 23697
rect 9299 23663 9337 23697
rect 9371 23663 9409 23697
rect 9443 23663 9481 23697
rect 9515 23663 9553 23697
rect 9587 23663 9625 23697
rect 9659 23663 9697 23697
rect 9731 23663 9769 23697
rect 9803 23663 9841 23697
rect 9875 23663 9913 23697
rect 9947 23663 9985 23697
rect 10019 23663 10057 23697
rect 10091 23663 10129 23697
rect 10163 23663 10201 23697
rect 10235 23663 10273 23697
rect 10307 23663 10345 23697
rect 10379 23663 10417 23697
rect 10451 23663 10489 23697
rect 10523 23663 10561 23697
rect 10595 23663 10633 23697
rect 10667 23663 10705 23697
rect 10739 23663 10777 23697
rect 10811 23663 10849 23697
rect 10883 23663 10921 23697
rect 10955 23663 10993 23697
rect 11027 23663 11065 23697
rect 11099 23663 11137 23697
rect 11171 23663 11209 23697
rect 11243 23663 11281 23697
rect 11315 23663 11353 23697
rect 11387 23663 11425 23697
rect 11459 23663 11497 23697
rect 11531 23663 11569 23697
rect 11603 23663 11641 23697
rect 11675 23663 11713 23697
rect 11747 23663 11785 23697
rect 11819 23663 11857 23697
rect 11891 23663 11929 23697
rect 11963 23663 12001 23697
rect 12035 23663 12073 23697
rect 12107 23663 12145 23697
rect 12179 23663 12217 23697
rect 12251 23663 12289 23697
rect 12323 23663 12361 23697
rect 12395 23663 12433 23697
rect 12467 23663 12505 23697
rect 12539 23663 12577 23697
rect 12611 23663 12649 23697
rect 12683 23663 12721 23697
rect 12755 23663 12793 23697
rect 12827 23663 12865 23697
rect 12899 23663 12937 23697
rect 12971 23663 13009 23697
rect 13043 23663 13081 23697
rect 13115 23663 13153 23697
rect 13187 23663 13225 23697
rect 13259 23663 13297 23697
rect 13331 23663 13343 23697
rect 5278 23651 5301 23663
rect 5353 23651 5376 23663
rect 5428 23651 5451 23663
rect 5503 23651 13343 23663
rect 5069 23627 13343 23651
rect 5069 23575 5075 23627
rect 5127 23575 5151 23627
rect 5203 23575 5226 23627
rect 5278 23575 5301 23627
rect 5353 23575 5376 23627
rect 5428 23575 5451 23627
rect 5503 23575 13343 23627
rect 5069 23551 13343 23575
rect 5069 23499 5075 23551
rect 5127 23499 5151 23551
rect 5203 23499 5226 23551
rect 5278 23499 5301 23551
rect 5353 23499 5376 23551
rect 5428 23499 5451 23551
rect 5503 23499 13343 23551
rect 5069 23475 13343 23499
rect 5069 23423 5075 23475
rect 5127 23423 5151 23475
rect 5203 23423 5226 23475
rect 5278 23462 5301 23475
rect 5353 23462 5376 23475
rect 5428 23462 5451 23475
rect 5503 23462 13343 23475
rect 5278 23428 5300 23462
rect 5353 23428 5373 23462
rect 5428 23428 5446 23462
rect 5503 23428 5519 23462
rect 5553 23428 5592 23462
rect 5626 23428 5665 23462
rect 5699 23428 5737 23462
rect 5771 23428 5809 23462
rect 5843 23428 5881 23462
rect 5915 23428 5953 23462
rect 5987 23428 6025 23462
rect 6059 23428 6097 23462
rect 6131 23428 6169 23462
rect 6203 23428 6241 23462
rect 6275 23428 6313 23462
rect 6347 23428 6385 23462
rect 6419 23428 6457 23462
rect 6491 23428 6529 23462
rect 6563 23428 6601 23462
rect 6635 23428 6673 23462
rect 6707 23428 6745 23462
rect 6779 23428 6817 23462
rect 6851 23428 6889 23462
rect 6923 23428 6961 23462
rect 6995 23428 7033 23462
rect 7067 23428 7105 23462
rect 7139 23428 7177 23462
rect 7211 23428 7249 23462
rect 7283 23428 7321 23462
rect 7355 23428 7393 23462
rect 7427 23428 7465 23462
rect 7499 23428 7537 23462
rect 7571 23428 7609 23462
rect 7643 23428 7681 23462
rect 7715 23428 7753 23462
rect 7787 23428 7825 23462
rect 7859 23428 7897 23462
rect 7931 23428 7969 23462
rect 8003 23428 8041 23462
rect 8075 23428 8113 23462
rect 8147 23428 8185 23462
rect 8219 23428 8257 23462
rect 8291 23428 8329 23462
rect 8363 23428 8401 23462
rect 8435 23428 8473 23462
rect 8507 23428 8545 23462
rect 8579 23428 8617 23462
rect 8651 23428 8689 23462
rect 8723 23428 8761 23462
rect 8795 23428 8833 23462
rect 8867 23428 8905 23462
rect 8939 23428 8977 23462
rect 9011 23428 9049 23462
rect 9083 23428 9121 23462
rect 9155 23428 9193 23462
rect 9227 23428 9265 23462
rect 9299 23428 9337 23462
rect 9371 23428 9409 23462
rect 9443 23428 9481 23462
rect 9515 23428 9553 23462
rect 9587 23428 9625 23462
rect 9659 23428 9697 23462
rect 9731 23428 9769 23462
rect 9803 23428 9841 23462
rect 9875 23428 9913 23462
rect 9947 23428 9985 23462
rect 10019 23428 10057 23462
rect 10091 23428 10129 23462
rect 10163 23428 10201 23462
rect 10235 23428 10273 23462
rect 10307 23428 10345 23462
rect 10379 23428 10417 23462
rect 10451 23428 10489 23462
rect 10523 23428 10561 23462
rect 10595 23428 10633 23462
rect 10667 23428 10705 23462
rect 10739 23428 10777 23462
rect 10811 23428 10849 23462
rect 10883 23428 10921 23462
rect 10955 23428 10993 23462
rect 11027 23428 11065 23462
rect 11099 23428 11137 23462
rect 11171 23428 11209 23462
rect 11243 23428 11281 23462
rect 11315 23428 11353 23462
rect 11387 23428 11425 23462
rect 11459 23428 11497 23462
rect 11531 23428 11569 23462
rect 11603 23428 11641 23462
rect 11675 23428 11713 23462
rect 11747 23428 11785 23462
rect 11819 23428 11857 23462
rect 11891 23428 11929 23462
rect 11963 23428 12001 23462
rect 12035 23428 12073 23462
rect 12107 23428 12145 23462
rect 12179 23428 12217 23462
rect 12251 23428 12289 23462
rect 12323 23428 12361 23462
rect 12395 23428 12433 23462
rect 12467 23428 12505 23462
rect 12539 23428 12577 23462
rect 12611 23428 12649 23462
rect 12683 23428 12721 23462
rect 12755 23428 12793 23462
rect 12827 23428 12865 23462
rect 12899 23428 12937 23462
rect 12971 23428 13009 23462
rect 13043 23428 13081 23462
rect 13115 23428 13153 23462
rect 13187 23428 13225 23462
rect 13259 23428 13297 23462
rect 13331 23428 13343 23462
rect 5278 23423 5301 23428
rect 5353 23423 5376 23428
rect 5428 23423 5451 23428
rect 5503 23423 13343 23428
rect 5069 23422 13343 23423
rect 4332 23076 4727 23110
rect 4761 23076 4767 23110
tri 13358 23078 13515 23235 se
rect 13515 23078 13521 24004
rect 4332 23037 4767 23076
rect 4332 23003 4727 23037
rect 4761 23003 4767 23037
rect 4332 22964 4767 23003
rect 4332 22930 4727 22964
rect 4761 22930 4767 22964
rect 4332 22891 4767 22930
rect 4332 22857 4727 22891
rect 4761 22857 4767 22891
rect 4332 22818 4767 22857
rect 4332 22784 4727 22818
rect 4761 22784 4767 22818
rect 4332 22745 4767 22784
rect 4332 22711 4727 22745
rect 4761 22711 4767 22745
rect 4332 22672 4767 22711
rect 4332 22638 4727 22672
rect 4761 22638 4767 22672
rect 4332 22599 4767 22638
rect 4332 22565 4727 22599
rect 4761 22565 4767 22599
rect 4332 22526 4767 22565
rect 4332 22492 4727 22526
rect 4761 22492 4767 22526
rect 4332 22453 4767 22492
rect 4332 22419 4727 22453
rect 4761 22419 4767 22453
rect 4332 22380 4767 22419
rect 4332 22346 4727 22380
rect 4761 22346 4767 22380
rect 4332 22306 4767 22346
rect 4332 22272 4727 22306
rect 4761 22272 4767 22306
rect 4332 22232 4767 22272
rect 4332 22198 4727 22232
rect 4761 22198 4767 22232
rect 4332 22158 4767 22198
rect 4332 22124 4727 22158
rect 4761 22124 4767 22158
rect 4332 22084 4767 22124
rect 4332 22050 4727 22084
rect 4761 22050 4767 22084
rect 5067 23066 13521 23078
rect 5067 23032 5073 23066
rect 5107 23054 13521 23066
rect 5107 23032 6718 23054
rect 5067 23020 6718 23032
rect 6752 23020 8374 23054
rect 8408 23020 10030 23054
rect 10064 23020 11686 23054
rect 11720 23020 13342 23054
rect 13376 23020 13521 23054
rect 5067 22993 13521 23020
rect 5067 22959 5073 22993
rect 5107 22976 13521 22993
rect 5107 22959 6718 22976
rect 5067 22942 6718 22959
rect 6752 22942 8374 22976
rect 8408 22942 10030 22976
rect 10064 22942 11686 22976
rect 11720 22942 13342 22976
rect 13376 22942 13521 22976
rect 5067 22920 13521 22942
rect 5067 22886 5073 22920
rect 5107 22898 13521 22920
rect 5107 22886 6718 22898
rect 5067 22864 6718 22886
rect 6752 22864 8374 22898
rect 8408 22864 10030 22898
rect 10064 22864 11686 22898
rect 11720 22864 13342 22898
rect 13376 22864 13521 22898
rect 5067 22847 13521 22864
rect 5067 22813 5073 22847
rect 5107 22820 13521 22847
rect 5107 22813 6718 22820
rect 5067 22786 6718 22813
rect 6752 22786 8374 22820
rect 8408 22786 10030 22820
rect 10064 22786 11686 22820
rect 11720 22786 13342 22820
rect 13376 22786 13521 22820
rect 5067 22774 13521 22786
rect 5067 22740 5073 22774
rect 5107 22742 13521 22774
rect 5107 22740 6718 22742
rect 5067 22708 6718 22740
rect 6752 22708 8374 22742
rect 8408 22708 10030 22742
rect 10064 22708 11686 22742
rect 11720 22708 13342 22742
rect 13376 22708 13521 22742
rect 5067 22701 13521 22708
rect 5067 22667 5073 22701
rect 5107 22667 13521 22701
rect 5067 22664 13521 22667
rect 5067 22630 6718 22664
rect 6752 22630 8374 22664
rect 8408 22630 10030 22664
rect 10064 22630 11686 22664
rect 11720 22630 13342 22664
rect 13376 22630 13521 22664
rect 5067 22628 13521 22630
rect 5067 22594 5073 22628
rect 5107 22594 13521 22628
rect 5067 22586 13521 22594
rect 5067 22556 6718 22586
rect 5067 22522 5073 22556
rect 5107 22552 6718 22556
rect 6752 22552 8374 22586
rect 8408 22552 10030 22586
rect 10064 22552 11686 22586
rect 11720 22552 13342 22586
rect 13376 22552 13521 22586
rect 5107 22522 13521 22552
rect 5067 22509 13521 22522
rect 5067 22484 6718 22509
rect 5067 22450 5073 22484
rect 5107 22475 6718 22484
rect 6752 22475 8374 22509
rect 8408 22475 10030 22509
rect 10064 22475 11686 22509
rect 11720 22475 13342 22509
rect 13376 22475 13521 22509
rect 5107 22450 13521 22475
rect 5067 22432 13521 22450
rect 5067 22412 6718 22432
rect 5067 22378 5073 22412
rect 5107 22398 6718 22412
rect 6752 22398 8374 22432
rect 8408 22398 10030 22432
rect 10064 22398 11686 22432
rect 11720 22398 13342 22432
rect 13376 22398 13521 22432
rect 5107 22378 13521 22398
rect 5067 22355 13521 22378
rect 5067 22340 6718 22355
rect 5067 22306 5073 22340
rect 5107 22321 6718 22340
rect 6752 22321 8374 22355
rect 8408 22321 10030 22355
rect 10064 22321 11686 22355
rect 11720 22321 13342 22355
rect 13376 22321 13521 22355
rect 5107 22306 13521 22321
rect 5067 22278 13521 22306
rect 5067 22268 6718 22278
rect 5067 22234 5073 22268
rect 5107 22244 6718 22268
rect 6752 22244 8374 22278
rect 8408 22244 10030 22278
rect 10064 22244 11686 22278
rect 11720 22244 13342 22278
rect 13376 22244 13521 22278
rect 5107 22234 13521 22244
rect 5067 22217 13521 22234
rect 13699 22217 13705 39099
rect 5067 22201 13705 22217
rect 5067 22196 6718 22201
rect 5067 22162 5073 22196
rect 5107 22167 6718 22196
rect 6752 22167 8374 22201
rect 8408 22167 10030 22201
rect 10064 22167 11686 22201
rect 11720 22167 13342 22201
rect 13376 22178 13705 22201
rect 13376 22167 13521 22178
rect 5107 22162 13521 22167
rect 5067 22144 13521 22162
rect 13555 22144 13593 22178
rect 13627 22144 13665 22178
rect 13699 22144 13705 22178
rect 5067 22124 13705 22144
rect 5067 22090 5073 22124
rect 5107 22090 6718 22124
rect 6752 22090 8374 22124
rect 8408 22090 10030 22124
rect 10064 22090 11686 22124
rect 11720 22090 13342 22124
rect 13376 22105 13705 22124
rect 13376 22090 13521 22105
rect 5067 22078 13521 22090
tri 13358 22071 13365 22078 ne
rect 13365 22071 13521 22078
rect 13555 22071 13593 22105
rect 13627 22071 13665 22105
rect 13699 22071 13705 22105
tri 13365 22055 13381 22071 ne
rect 13381 22055 13705 22071
rect 4332 22010 4767 22050
tri 13381 22032 13404 22055 ne
rect 13404 22032 13705 22055
rect 4332 21976 4727 22010
rect 4761 21976 4767 22010
tri 13404 21998 13438 22032 ne
rect 13438 21998 13521 22032
rect 13555 21998 13593 22032
rect 13627 21998 13665 22032
rect 13699 21998 13705 22032
tri 13438 21982 13454 21998 ne
rect 13454 21982 13705 21998
rect 4332 21635 4767 21976
tri 13454 21959 13477 21982 ne
rect 13477 21959 13705 21982
tri 13477 21925 13511 21959 ne
rect 13511 21925 13521 21959
rect 13555 21925 13593 21959
rect 13627 21925 13665 21959
rect 13699 21925 13705 21959
tri 13511 21921 13515 21925 ne
rect 13515 21886 13705 21925
rect 13515 21852 13521 21886
rect 13555 21852 13593 21886
rect 13627 21852 13665 21886
rect 13699 21852 13705 21886
rect 13515 21813 13705 21852
rect 13515 21779 13521 21813
rect 13555 21779 13593 21813
rect 13627 21779 13665 21813
rect 13699 21779 13705 21813
rect 5067 21723 5073 21775
rect 5125 21723 5140 21775
rect 5192 21723 5206 21775
rect 5258 21763 5272 21775
rect 5324 21769 5330 21775
tri 5330 21769 5336 21775 sw
rect 5324 21763 13343 21769
rect 5259 21729 5272 21763
rect 5332 21729 5371 21763
rect 5405 21729 5444 21763
rect 5478 21729 5517 21763
rect 5551 21729 5590 21763
rect 5624 21729 5663 21763
rect 5697 21729 5736 21763
rect 5770 21729 5809 21763
rect 5843 21729 5881 21763
rect 5915 21729 5953 21763
rect 5987 21729 6025 21763
rect 6059 21729 6097 21763
rect 6131 21729 6169 21763
rect 6203 21729 6241 21763
rect 6275 21729 6313 21763
rect 6347 21729 6385 21763
rect 6419 21729 6457 21763
rect 6491 21729 6529 21763
rect 6563 21729 6601 21763
rect 6635 21729 6673 21763
rect 6707 21729 6745 21763
rect 6779 21729 6817 21763
rect 6851 21729 6889 21763
rect 6923 21729 6961 21763
rect 6995 21729 7033 21763
rect 7067 21729 7105 21763
rect 7139 21729 7177 21763
rect 7211 21729 7249 21763
rect 7283 21729 7321 21763
rect 7355 21729 7393 21763
rect 7427 21729 7465 21763
rect 7499 21729 7537 21763
rect 7571 21729 7609 21763
rect 7643 21729 7681 21763
rect 7715 21729 7753 21763
rect 7787 21729 7825 21763
rect 7859 21729 7897 21763
rect 7931 21729 7969 21763
rect 8003 21729 8041 21763
rect 8075 21729 8113 21763
rect 8147 21729 8185 21763
rect 8219 21729 8257 21763
rect 8291 21729 8329 21763
rect 8363 21729 8401 21763
rect 8435 21729 8473 21763
rect 8507 21729 8545 21763
rect 8579 21729 8617 21763
rect 8651 21729 8689 21763
rect 8723 21729 8761 21763
rect 8795 21729 8833 21763
rect 8867 21729 8905 21763
rect 8939 21729 8977 21763
rect 9011 21729 9049 21763
rect 9083 21729 9121 21763
rect 9155 21729 9193 21763
rect 9227 21729 9265 21763
rect 9299 21729 9337 21763
rect 9371 21729 9409 21763
rect 9443 21729 9481 21763
rect 9515 21729 9553 21763
rect 9587 21729 9625 21763
rect 9659 21729 9697 21763
rect 9731 21729 9769 21763
rect 9803 21729 9841 21763
rect 9875 21729 9913 21763
rect 9947 21729 9985 21763
rect 10019 21729 10057 21763
rect 10091 21729 10129 21763
rect 10163 21729 10201 21763
rect 10235 21729 10273 21763
rect 10307 21729 10345 21763
rect 10379 21729 10417 21763
rect 10451 21729 10489 21763
rect 10523 21729 10561 21763
rect 10595 21729 10633 21763
rect 10667 21729 10705 21763
rect 10739 21729 10777 21763
rect 10811 21729 10849 21763
rect 10883 21729 10921 21763
rect 10955 21729 10993 21763
rect 11027 21729 11065 21763
rect 11099 21729 11137 21763
rect 11171 21729 11209 21763
rect 11243 21729 11281 21763
rect 11315 21729 11353 21763
rect 11387 21729 11425 21763
rect 11459 21729 11497 21763
rect 11531 21729 11569 21763
rect 11603 21729 11641 21763
rect 11675 21729 11713 21763
rect 11747 21729 11785 21763
rect 11819 21729 11857 21763
rect 11891 21729 11929 21763
rect 11963 21729 12001 21763
rect 12035 21729 12073 21763
rect 12107 21729 12145 21763
rect 12179 21729 12217 21763
rect 12251 21729 12289 21763
rect 12323 21729 12361 21763
rect 12395 21729 12433 21763
rect 12467 21729 12505 21763
rect 12539 21729 12577 21763
rect 12611 21729 12649 21763
rect 12683 21729 12721 21763
rect 12755 21729 12793 21763
rect 12827 21729 12865 21763
rect 12899 21729 12937 21763
rect 12971 21729 13009 21763
rect 13043 21729 13081 21763
rect 13115 21729 13153 21763
rect 13187 21729 13225 21763
rect 13259 21729 13297 21763
rect 13331 21729 13343 21763
rect 5258 21723 5272 21729
rect 5324 21723 13343 21729
rect 13515 21740 13705 21779
rect 4332 21601 4727 21635
rect 4761 21601 4767 21635
rect 4332 21561 4767 21601
rect 4332 21527 4727 21561
rect 4761 21527 4767 21561
rect 4332 21487 4767 21527
rect 4332 21453 4727 21487
rect 4761 21453 4767 21487
rect 4332 21413 4767 21453
rect 13515 21706 13521 21740
rect 13555 21706 13593 21740
rect 13627 21706 13665 21740
rect 13699 21706 13705 21740
rect 13515 21667 13705 21706
rect 13515 21633 13521 21667
rect 13555 21633 13593 21667
rect 13627 21633 13665 21667
rect 13699 21633 13705 21667
rect 13515 21594 13705 21633
rect 13515 21560 13521 21594
rect 13555 21560 13593 21594
rect 13627 21560 13665 21594
rect 13699 21560 13705 21594
rect 13515 21521 13705 21560
rect 13515 21487 13521 21521
rect 13555 21487 13593 21521
rect 13627 21487 13665 21521
rect 13699 21487 13705 21521
rect 13515 21448 13705 21487
tri 13510 21414 13515 21419 se
rect 13515 21414 13521 21448
rect 13555 21414 13593 21448
rect 13627 21414 13665 21448
rect 13699 21414 13705 21448
rect 4332 21379 4727 21413
rect 4761 21379 4767 21413
rect 4332 21339 4767 21379
tri 13471 21375 13510 21414 se
rect 13510 21375 13705 21414
tri 13437 21341 13471 21375 se
rect 13471 21341 13521 21375
rect 13555 21341 13593 21375
rect 13627 21341 13665 21375
rect 13699 21341 13705 21375
rect 4332 21305 4727 21339
rect 4761 21305 4767 21339
tri 13425 21329 13437 21341 se
rect 13437 21329 13705 21341
rect 4332 21265 4767 21305
tri 13398 21302 13425 21329 se
rect 13425 21302 13705 21329
tri 13364 21268 13398 21302 se
rect 13398 21268 13521 21302
rect 13555 21268 13593 21302
rect 13627 21268 13665 21302
rect 13699 21268 13705 21302
rect 4332 21231 4727 21265
rect 4761 21231 4767 21265
tri 13359 21263 13364 21268 se
rect 13364 21263 13705 21268
rect 4332 21191 4767 21231
rect 4332 21157 4727 21191
rect 4761 21157 4767 21191
rect 4332 21117 4767 21157
rect 4332 21083 4727 21117
rect 4761 21083 4767 21117
rect 4332 21043 4767 21083
rect 4332 21009 4727 21043
rect 4761 21009 4767 21043
rect 4332 20969 4767 21009
rect 4332 20935 4727 20969
rect 4761 20935 4767 20969
rect 4332 20895 4767 20935
rect 4332 20861 4727 20895
rect 4761 20861 4767 20895
rect 4332 20822 4767 20861
rect 4332 20788 4727 20822
rect 4761 20788 4767 20822
rect 4332 20749 4767 20788
rect 4332 20715 4727 20749
rect 4761 20715 4767 20749
rect 4332 20676 4767 20715
rect 4332 20642 4727 20676
rect 4761 20642 4767 20676
rect 4332 20603 4767 20642
rect 4332 20569 4727 20603
rect 4761 20569 4767 20603
rect 4332 20530 4767 20569
rect 4332 20496 4727 20530
rect 4761 20496 4767 20530
rect 4332 20457 4767 20496
rect 4332 20423 4727 20457
rect 4761 20423 4767 20457
tri 418 20421 420 20423 se
rect 420 20421 3860 20423
tri 3860 20421 3862 20423 nw
tri 390 20393 418 20421 se
rect 418 20393 3832 20421
tri 3832 20393 3860 20421 nw
tri 389 20392 390 20393 se
rect 390 20392 3831 20393
tri 3831 20392 3832 20393 nw
tri 4331 20392 4332 20393 se
rect 4332 20392 4767 20423
tri 382 20385 389 20392 se
rect 389 20385 3824 20392
tri 3824 20385 3831 20392 nw
tri 4324 20385 4331 20392 se
rect 4331 20385 4767 20392
rect 382 20384 3823 20385
tri 3823 20384 3824 20385 nw
tri 4323 20384 4324 20385 se
rect 4324 20384 4767 20385
rect 382 20350 3789 20384
tri 3789 20350 3823 20384 nw
tri 4289 20350 4323 20384 se
rect 4323 20350 4727 20384
rect 4761 20350 4767 20384
rect 382 20349 3788 20350
tri 3788 20349 3789 20350 nw
tri 4288 20349 4289 20350 se
rect 4289 20349 4767 20350
rect 382 20339 3778 20349
tri 3778 20339 3788 20349 nw
tri 4278 20339 4288 20349 se
rect 4288 20339 4767 20349
rect 382 20319 524 20339
tri 524 20319 544 20339 nw
tri 4258 20319 4278 20339 se
rect 4278 20319 4767 20339
rect 382 20311 516 20319
tri 516 20311 524 20319 nw
tri 4250 20311 4258 20319 se
rect 4258 20311 4767 20319
rect 382 4606 500 20311
tri 500 20295 516 20311 nw
tri 4234 20295 4250 20311 se
rect 4250 20295 4727 20311
tri 4216 20277 4234 20295 se
rect 4234 20277 4727 20295
rect 4761 20277 4767 20311
tri 4204 20265 4216 20277 se
rect 4216 20265 4767 20277
rect 5067 21251 13705 21263
rect 5067 21217 5073 21251
rect 5107 21217 6718 21251
rect 6752 21217 8374 21251
rect 8408 21217 10030 21251
rect 10064 21217 11686 21251
rect 11720 21217 13342 21251
rect 13376 21229 13705 21251
rect 13376 21217 13521 21229
rect 5067 21195 13521 21217
rect 13555 21195 13593 21229
rect 13627 21195 13665 21229
rect 13699 21195 13705 21229
rect 5067 21178 13705 21195
rect 5067 21144 5073 21178
rect 5107 21144 6718 21178
rect 6752 21144 8374 21178
rect 8408 21144 10030 21178
rect 10064 21144 11686 21178
rect 11720 21144 13342 21178
rect 13376 21156 13705 21178
rect 13376 21144 13521 21156
rect 5067 21122 13521 21144
rect 13555 21122 13593 21156
rect 13627 21122 13665 21156
rect 13699 21122 13705 21156
rect 5067 21105 13705 21122
rect 5067 21071 5073 21105
rect 5107 21071 6718 21105
rect 6752 21071 8374 21105
rect 8408 21071 10030 21105
rect 10064 21071 11686 21105
rect 11720 21071 13342 21105
rect 13376 21083 13705 21105
rect 13376 21071 13521 21083
rect 5067 21049 13521 21071
rect 13555 21049 13593 21083
rect 13627 21049 13665 21083
rect 13699 21049 13705 21083
rect 5067 21032 13705 21049
rect 5067 20998 5073 21032
rect 5107 20998 6718 21032
rect 6752 20998 8374 21032
rect 8408 20998 10030 21032
rect 10064 20998 11686 21032
rect 11720 20998 13342 21032
rect 13376 21010 13705 21032
rect 13376 20998 13521 21010
rect 5067 20976 13521 20998
rect 13555 20976 13593 21010
rect 13627 20976 13665 21010
rect 13699 20976 13705 21010
rect 5067 20959 13705 20976
rect 5067 20925 5073 20959
rect 5107 20925 6718 20959
rect 6752 20925 8374 20959
rect 8408 20925 10030 20959
rect 10064 20925 11686 20959
rect 11720 20925 13342 20959
rect 13376 20937 13705 20959
rect 13376 20925 13521 20937
rect 5067 20903 13521 20925
rect 13555 20903 13593 20937
rect 13627 20903 13665 20937
rect 13699 20903 13705 20937
rect 5067 20887 13705 20903
rect 5067 20853 5073 20887
rect 5107 20853 6718 20887
rect 6752 20853 8374 20887
rect 8408 20853 10030 20887
rect 10064 20853 11686 20887
rect 11720 20853 13342 20887
rect 13376 20864 13705 20887
rect 13376 20853 13521 20864
rect 5067 20830 13521 20853
rect 13555 20830 13593 20864
rect 13627 20830 13665 20864
rect 13699 20830 13705 20864
rect 5067 20815 13705 20830
rect 5067 20781 5073 20815
rect 5107 20781 6718 20815
rect 6752 20781 8374 20815
rect 8408 20781 10030 20815
rect 10064 20781 11686 20815
rect 11720 20781 13342 20815
rect 13376 20791 13705 20815
rect 13376 20781 13521 20791
rect 5067 20757 13521 20781
rect 13555 20757 13593 20791
rect 13627 20757 13665 20791
rect 13699 20757 13705 20791
rect 5067 20743 13705 20757
rect 5067 20709 5073 20743
rect 5107 20709 6718 20743
rect 6752 20709 8374 20743
rect 8408 20709 10030 20743
rect 10064 20709 11686 20743
rect 11720 20709 13342 20743
rect 13376 20718 13705 20743
rect 13376 20709 13521 20718
rect 5067 20684 13521 20709
rect 13555 20684 13593 20718
rect 13627 20684 13665 20718
rect 13699 20684 13705 20718
rect 5067 20671 13705 20684
rect 5067 20637 5073 20671
rect 5107 20637 6718 20671
rect 6752 20637 8374 20671
rect 8408 20637 10030 20671
rect 10064 20637 11686 20671
rect 11720 20637 13342 20671
rect 13376 20645 13705 20671
rect 13376 20637 13521 20645
rect 5067 20611 13521 20637
rect 13555 20611 13593 20645
rect 13627 20611 13665 20645
rect 13699 20611 13705 20645
rect 5067 20599 13705 20611
rect 5067 20565 5073 20599
rect 5107 20565 6718 20599
rect 6752 20565 8374 20599
rect 8408 20565 10030 20599
rect 10064 20565 11686 20599
rect 11720 20565 13342 20599
rect 13376 20572 13705 20599
rect 13376 20565 13521 20572
rect 5067 20538 13521 20565
rect 13555 20538 13593 20572
rect 13627 20538 13665 20572
rect 13699 20538 13705 20572
rect 5067 20527 13705 20538
rect 5067 20493 5073 20527
rect 5107 20493 6718 20527
rect 6752 20493 8374 20527
rect 8408 20493 10030 20527
rect 10064 20493 11686 20527
rect 11720 20493 13342 20527
rect 13376 20499 13705 20527
rect 13376 20493 13521 20499
rect 5067 20465 13521 20493
rect 13555 20465 13593 20499
rect 13627 20465 13665 20499
rect 13699 20465 13705 20499
rect 5067 20455 13705 20465
rect 5067 20421 5073 20455
rect 5107 20421 6718 20455
rect 6752 20421 8374 20455
rect 8408 20421 10030 20455
rect 10064 20421 11686 20455
rect 11720 20421 13342 20455
rect 13376 20426 13705 20455
rect 13376 20421 13521 20426
rect 5067 20392 13521 20421
rect 13555 20392 13593 20426
rect 13627 20392 13665 20426
rect 13699 20392 13705 20426
rect 5067 20383 13705 20392
rect 5067 20349 5073 20383
rect 5107 20349 6718 20383
rect 6752 20349 8374 20383
rect 8408 20349 10030 20383
rect 10064 20349 11686 20383
rect 11720 20349 13342 20383
rect 13376 20353 13705 20383
rect 13376 20349 13521 20353
rect 5067 20319 13521 20349
rect 13555 20319 13593 20353
rect 13627 20319 13665 20353
rect 13699 20319 13705 20353
rect 5067 20311 13705 20319
rect 5067 20277 5073 20311
rect 5107 20277 6718 20311
rect 6752 20277 8374 20311
rect 8408 20277 10030 20311
rect 10064 20277 11686 20311
rect 11720 20277 13342 20311
rect 13376 20280 13705 20311
rect 13376 20277 13521 20280
rect 5067 20265 13521 20277
tri 4185 20246 4204 20265 se
rect 4204 20246 4767 20265
tri 13411 20246 13430 20265 ne
rect 13430 20246 13521 20265
rect 13555 20246 13593 20280
rect 13627 20246 13665 20280
rect 13699 20246 13705 20280
tri 4146 20207 4185 20246 se
rect 4185 20210 4767 20246
rect 4185 20207 4764 20210
tri 4764 20207 4767 20210 nw
tri 13430 20207 13469 20246 ne
rect 13469 20207 13705 20246
tri 4112 20173 4146 20207 se
rect 4146 20173 4730 20207
tri 4730 20173 4764 20207 nw
tri 13469 20173 13503 20207 ne
rect 13503 20173 13521 20207
rect 13555 20173 13593 20207
rect 13627 20173 13665 20207
rect 13699 20173 13705 20207
tri 4100 20161 4112 20173 se
rect 4112 20161 4718 20173
tri 4718 20161 4730 20173 nw
tri 13503 20161 13515 20173 ne
rect 13515 20161 13705 20173
rect 13832 26620 13838 39364
rect 13944 26620 13950 39470
rect 13832 26581 13950 26620
rect 13832 26547 13838 26581
rect 13872 26547 13910 26581
rect 13944 26547 13950 26581
rect 13832 26508 13950 26547
rect 13832 26474 13838 26508
rect 13872 26474 13910 26508
rect 13944 26474 13950 26508
rect 13832 26435 13950 26474
rect 13832 26401 13838 26435
rect 13872 26401 13910 26435
rect 13944 26401 13950 26435
rect 13832 26362 13950 26401
rect 13832 26328 13838 26362
rect 13872 26328 13910 26362
rect 13944 26328 13950 26362
rect 13832 26289 13950 26328
rect 13832 26255 13838 26289
rect 13872 26255 13910 26289
rect 13944 26255 13950 26289
rect 13832 26216 13950 26255
rect 13832 26182 13838 26216
rect 13872 26182 13910 26216
rect 13944 26182 13950 26216
rect 13832 26143 13950 26182
rect 13832 26109 13838 26143
rect 13872 26109 13910 26143
rect 13944 26109 13950 26143
rect 13832 26070 13950 26109
rect 13832 26036 13838 26070
rect 13872 26036 13910 26070
rect 13944 26036 13950 26070
rect 13832 25997 13950 26036
rect 13832 25963 13838 25997
rect 13872 25963 13910 25997
rect 13944 25963 13950 25997
rect 13832 25924 13950 25963
rect 13832 25890 13838 25924
rect 13872 25890 13910 25924
rect 13944 25890 13950 25924
rect 13832 25851 13950 25890
rect 13832 25817 13838 25851
rect 13872 25817 13910 25851
rect 13944 25817 13950 25851
rect 13832 25778 13950 25817
rect 13832 25744 13838 25778
rect 13872 25744 13910 25778
rect 13944 25744 13950 25778
rect 13832 25705 13950 25744
rect 13832 25671 13838 25705
rect 13872 25671 13910 25705
rect 13944 25671 13950 25705
rect 13832 25632 13950 25671
rect 13832 25598 13838 25632
rect 13872 25598 13910 25632
rect 13944 25598 13950 25632
rect 13832 25559 13950 25598
rect 13832 25525 13838 25559
rect 13872 25525 13910 25559
rect 13944 25525 13950 25559
rect 13832 25486 13950 25525
rect 13832 25452 13838 25486
rect 13872 25452 13910 25486
rect 13944 25452 13950 25486
rect 13832 25413 13950 25452
rect 13832 25379 13838 25413
rect 13872 25379 13910 25413
rect 13944 25379 13950 25413
rect 13832 25340 13950 25379
rect 13832 25306 13838 25340
rect 13872 25306 13910 25340
rect 13944 25306 13950 25340
rect 13832 25267 13950 25306
rect 13832 25233 13838 25267
rect 13872 25233 13910 25267
rect 13944 25233 13950 25267
rect 13832 25194 13950 25233
rect 13832 25160 13838 25194
rect 13872 25160 13910 25194
rect 13944 25160 13950 25194
rect 13832 25121 13950 25160
rect 13832 25087 13838 25121
rect 13872 25087 13910 25121
rect 13944 25087 13950 25121
rect 13832 25048 13950 25087
rect 13832 25014 13838 25048
rect 13872 25014 13910 25048
rect 13944 25014 13950 25048
rect 13832 24975 13950 25014
rect 13832 24941 13838 24975
rect 13872 24941 13910 24975
rect 13944 24941 13950 24975
rect 13832 24902 13950 24941
rect 13832 24868 13838 24902
rect 13872 24868 13910 24902
rect 13944 24868 13950 24902
rect 13832 24829 13950 24868
rect 13832 24795 13838 24829
rect 13872 24795 13910 24829
rect 13944 24795 13950 24829
rect 13832 24756 13950 24795
rect 13832 24722 13838 24756
rect 13872 24722 13910 24756
rect 13944 24722 13950 24756
rect 13832 24683 13950 24722
rect 13832 24649 13838 24683
rect 13872 24649 13910 24683
rect 13944 24649 13950 24683
rect 13832 24610 13950 24649
rect 13832 24576 13838 24610
rect 13872 24576 13910 24610
rect 13944 24576 13950 24610
rect 13832 24537 13950 24576
rect 13832 24503 13838 24537
rect 13872 24503 13910 24537
rect 13944 24503 13950 24537
rect 13832 24464 13950 24503
rect 13832 24430 13838 24464
rect 13872 24430 13910 24464
rect 13944 24430 13950 24464
rect 13832 24391 13950 24430
rect 13832 24357 13838 24391
rect 13872 24357 13910 24391
rect 13944 24357 13950 24391
rect 13832 24318 13950 24357
rect 13832 24284 13838 24318
rect 13872 24284 13910 24318
rect 13944 24284 13950 24318
rect 13832 24245 13950 24284
rect 13832 24211 13838 24245
rect 13872 24211 13910 24245
rect 13944 24211 13950 24245
rect 13832 24172 13950 24211
rect 13832 24138 13838 24172
rect 13872 24138 13910 24172
rect 13944 24138 13950 24172
rect 13832 24099 13950 24138
rect 13832 24065 13838 24099
rect 13872 24065 13910 24099
rect 13944 24065 13950 24099
rect 13832 24026 13950 24065
rect 13832 23992 13838 24026
rect 13872 23992 13910 24026
rect 13944 23992 13950 24026
rect 13832 23953 13950 23992
rect 13832 23919 13838 23953
rect 13872 23919 13910 23953
rect 13944 23919 13950 23953
rect 13832 23880 13950 23919
rect 13832 23846 13838 23880
rect 13872 23846 13910 23880
rect 13944 23846 13950 23880
rect 13832 23807 13950 23846
rect 13832 23773 13838 23807
rect 13872 23773 13910 23807
rect 13944 23773 13950 23807
rect 13832 23734 13950 23773
rect 13832 23700 13838 23734
rect 13872 23700 13910 23734
rect 13944 23700 13950 23734
rect 13832 23661 13950 23700
rect 13832 23627 13838 23661
rect 13872 23627 13910 23661
rect 13944 23627 13950 23661
rect 13832 23588 13950 23627
rect 13832 23554 13838 23588
rect 13872 23554 13910 23588
rect 13944 23554 13950 23588
rect 13832 23515 13950 23554
rect 13832 23481 13838 23515
rect 13872 23481 13910 23515
rect 13944 23481 13950 23515
rect 13832 23442 13950 23481
rect 13832 23408 13838 23442
rect 13872 23408 13910 23442
rect 13944 23408 13950 23442
rect 13832 23369 13950 23408
rect 13832 23335 13838 23369
rect 13872 23335 13910 23369
rect 13944 23335 13950 23369
rect 13832 23296 13950 23335
rect 13832 23262 13838 23296
rect 13872 23262 13910 23296
rect 13944 23262 13950 23296
rect 13832 23223 13950 23262
rect 13832 23189 13838 23223
rect 13872 23189 13910 23223
rect 13944 23189 13950 23223
rect 13832 23150 13950 23189
rect 13832 23116 13838 23150
rect 13872 23116 13910 23150
rect 13944 23116 13950 23150
rect 13832 23077 13950 23116
rect 13832 23043 13838 23077
rect 13872 23043 13910 23077
rect 13944 23043 13950 23077
rect 13832 23004 13950 23043
rect 13832 22970 13838 23004
rect 13872 22970 13910 23004
rect 13944 22970 13950 23004
rect 13832 22931 13950 22970
rect 13832 22897 13838 22931
rect 13872 22897 13910 22931
rect 13944 22897 13950 22931
rect 13832 22858 13950 22897
rect 13832 22824 13838 22858
rect 13872 22824 13910 22858
rect 13944 22824 13950 22858
rect 13832 22785 13950 22824
rect 13832 22751 13838 22785
rect 13872 22751 13910 22785
rect 13944 22751 13950 22785
rect 13832 22712 13950 22751
rect 13832 22678 13838 22712
rect 13872 22678 13910 22712
rect 13944 22678 13950 22712
rect 13832 22639 13950 22678
rect 13832 22605 13838 22639
rect 13872 22605 13910 22639
rect 13944 22605 13950 22639
rect 13832 22566 13950 22605
rect 13832 22532 13838 22566
rect 13872 22532 13910 22566
rect 13944 22532 13950 22566
rect 13832 22493 13950 22532
rect 13832 22459 13838 22493
rect 13872 22459 13910 22493
rect 13944 22459 13950 22493
rect 13832 22420 13950 22459
rect 13832 22386 13838 22420
rect 13872 22386 13910 22420
rect 13944 22386 13950 22420
rect 13832 22347 13950 22386
rect 13832 22313 13838 22347
rect 13872 22313 13910 22347
rect 13944 22313 13950 22347
rect 13832 22274 13950 22313
rect 13832 22240 13838 22274
rect 13872 22240 13910 22274
rect 13944 22240 13950 22274
rect 13832 22201 13950 22240
rect 13832 22167 13838 22201
rect 13872 22167 13910 22201
rect 13944 22167 13950 22201
rect 13832 22128 13950 22167
rect 13832 22094 13838 22128
rect 13872 22094 13910 22128
rect 13944 22094 13950 22128
rect 13832 22055 13950 22094
rect 13832 22021 13838 22055
rect 13872 22021 13910 22055
rect 13944 22021 13950 22055
rect 13832 21982 13950 22021
rect 13832 21948 13838 21982
rect 13872 21948 13910 21982
rect 13944 21948 13950 21982
rect 13832 21909 13950 21948
rect 13832 21875 13838 21909
rect 13872 21875 13910 21909
rect 13944 21875 13950 21909
rect 13832 21836 13950 21875
rect 13832 21802 13838 21836
rect 13872 21802 13910 21836
rect 13944 21802 13950 21836
rect 13832 21763 13950 21802
rect 13832 21729 13838 21763
rect 13872 21729 13910 21763
rect 13944 21729 13950 21763
rect 13832 21690 13950 21729
rect 13832 21656 13838 21690
rect 13872 21656 13910 21690
rect 13944 21656 13950 21690
rect 13832 21617 13950 21656
rect 13832 21583 13838 21617
rect 13872 21583 13910 21617
rect 13944 21583 13950 21617
rect 13832 21544 13950 21583
rect 13832 21510 13838 21544
rect 13872 21510 13910 21544
rect 13944 21510 13950 21544
rect 13832 21471 13950 21510
rect 13832 21437 13838 21471
rect 13872 21437 13910 21471
rect 13944 21437 13950 21471
rect 13832 21329 13950 21437
tri 3849 19910 4100 20161 se
rect 4100 19910 4453 20161
rect 1831 19898 1949 19910
rect 1831 19864 1837 19898
rect 1871 19864 1909 19898
rect 1943 19864 1949 19898
tri 3835 19896 3849 19910 se
rect 3849 19896 4453 19910
tri 4453 19896 4718 20161 nw
rect 1831 19821 1949 19864
rect 1831 19787 1837 19821
rect 1871 19787 1909 19821
rect 1943 19787 1949 19821
rect 1831 19744 1949 19787
rect 1831 19710 1837 19744
rect 1871 19710 1909 19744
rect 1943 19710 1949 19744
rect 1831 19667 1949 19710
rect 1831 19633 1837 19667
rect 1871 19633 1909 19667
rect 1943 19633 1949 19667
rect 1831 19580 1949 19633
tri 3832 19893 3835 19896 se
rect 3835 19893 4450 19896
tri 4450 19893 4453 19896 nw
rect 3832 19754 4311 19893
tri 4311 19754 4450 19893 nw
rect 3832 19745 4302 19754
tri 4302 19745 4311 19754 nw
rect 3832 19742 4299 19745
tri 4299 19742 4302 19745 nw
tri 1949 19580 1964 19595 sw
rect 1831 19578 1964 19580
tri 1964 19578 1966 19580 sw
rect 1831 19547 1966 19578
tri 1831 19544 1834 19547 ne
rect 1834 19544 1966 19547
tri 1966 19544 2000 19578 sw
tri 1834 19540 1838 19544 ne
rect 1838 19540 2000 19544
tri 2000 19540 2004 19544 sw
tri 1838 19506 1872 19540 ne
rect 1872 19506 2004 19540
tri 2004 19506 2038 19540 sw
tri 1872 19505 1873 19506 ne
rect 1873 19505 2038 19506
tri 2038 19505 2039 19506 sw
tri 1873 19489 1889 19505 ne
rect 1889 19489 2039 19505
tri 2039 19489 2055 19505 sw
tri 1889 19477 1901 19489 ne
rect 1901 19477 2055 19489
tri 1901 19443 1935 19477 ne
rect 1935 19443 1943 19477
rect 1977 19443 2015 19477
rect 2049 19443 2055 19477
tri 1935 19441 1937 19443 ne
rect 1937 19403 2055 19443
rect 1937 19369 1943 19403
rect 1977 19369 2015 19403
rect 2049 19369 2055 19403
rect 1937 19329 2055 19369
rect 1937 19295 1943 19329
rect 1977 19295 2015 19329
rect 2049 19295 2055 19329
rect 1937 19255 2055 19295
rect 1937 19221 1943 19255
rect 1977 19221 2015 19255
rect 2049 19221 2055 19255
rect 1937 19181 2055 19221
rect 1937 19147 1943 19181
rect 1977 19147 2015 19181
rect 2049 19147 2055 19181
rect 1937 19107 2055 19147
rect 1937 19073 1943 19107
rect 1977 19073 2015 19107
rect 2049 19073 2055 19107
rect 1937 19033 2055 19073
rect 1937 18999 1943 19033
rect 1977 18999 2015 19033
rect 2049 18999 2055 19033
rect 1937 18959 2055 18999
rect 1937 18925 1943 18959
rect 1977 18925 2015 18959
rect 2049 18925 2055 18959
rect 1937 18884 2055 18925
rect 1937 18850 1943 18884
rect 1977 18850 2015 18884
rect 2049 18850 2055 18884
rect 1937 18809 2055 18850
rect 1937 18775 1943 18809
rect 1977 18775 2015 18809
rect 2049 18775 2055 18809
rect 1937 18734 2055 18775
rect 1937 18700 1943 18734
rect 1977 18700 2015 18734
rect 2049 18700 2055 18734
rect 1937 18659 2055 18700
rect 1937 18625 1943 18659
rect 1977 18625 2015 18659
rect 2049 18625 2055 18659
rect 1937 18584 2055 18625
rect 1937 18550 1943 18584
rect 1977 18550 2015 18584
rect 2049 18550 2055 18584
rect 1937 18509 2055 18550
rect 1937 18475 1943 18509
rect 1977 18475 2015 18509
rect 2049 18475 2055 18509
rect 1937 18434 2055 18475
rect 1937 18400 1943 18434
rect 1977 18400 2015 18434
rect 2049 18400 2055 18434
rect 1937 18359 2055 18400
rect 1937 18325 1943 18359
rect 1977 18325 2015 18359
rect 2049 18325 2055 18359
rect 1937 18284 2055 18325
rect 1937 18250 1943 18284
rect 1977 18250 2015 18284
rect 2049 18250 2055 18284
rect 1937 18209 2055 18250
rect 1937 18175 1943 18209
rect 1977 18175 2015 18209
rect 2049 18175 2055 18209
rect 1937 18134 2055 18175
rect 1937 18100 1943 18134
rect 1977 18100 2015 18134
rect 2049 18100 2055 18134
rect 1937 18059 2055 18100
rect 1937 18025 1943 18059
rect 1977 18025 2015 18059
rect 2049 18025 2055 18059
rect 1937 17984 2055 18025
rect 1937 17950 1943 17984
rect 1977 17950 2015 17984
rect 2049 17950 2055 17984
rect 1937 17909 2055 17950
rect 1937 17875 1943 17909
rect 1977 17875 2015 17909
rect 2049 17875 2055 17909
rect 1937 17863 2055 17875
tri 3828 17605 3832 17609 se
rect 3832 17605 4268 19742
tri 4268 19711 4299 19742 nw
rect 4911 19702 4917 19754
rect 4969 19702 4981 19754
rect 5033 19748 5039 19754
tri 5039 19748 5045 19754 sw
rect 5033 19742 12975 19748
rect 5033 19708 5069 19742
rect 5103 19708 5142 19742
rect 5176 19708 5215 19742
rect 5249 19708 5288 19742
rect 5322 19708 5361 19742
rect 5395 19708 5434 19742
rect 5468 19708 5507 19742
rect 5541 19708 5580 19742
rect 5614 19708 5653 19742
rect 5687 19708 5726 19742
rect 5760 19708 5799 19742
rect 5833 19708 5872 19742
rect 5906 19708 5945 19742
rect 5979 19708 6017 19742
rect 6051 19708 6089 19742
rect 6123 19708 6161 19742
rect 6195 19708 6233 19742
rect 6267 19708 6305 19742
rect 6339 19708 6377 19742
rect 6411 19708 6449 19742
rect 6483 19708 6521 19742
rect 6555 19708 6593 19742
rect 6627 19708 6665 19742
rect 6699 19708 6737 19742
rect 6771 19708 6809 19742
rect 6843 19708 6881 19742
rect 6915 19708 6953 19742
rect 6987 19708 7025 19742
rect 7059 19708 7097 19742
rect 7131 19708 7169 19742
rect 7203 19708 7241 19742
rect 7275 19708 7313 19742
rect 7347 19708 7385 19742
rect 7419 19708 7457 19742
rect 7491 19708 7529 19742
rect 7563 19708 7601 19742
rect 7635 19708 7673 19742
rect 7707 19708 7745 19742
rect 7779 19708 7817 19742
rect 7851 19708 7889 19742
rect 7923 19708 7961 19742
rect 7995 19708 8033 19742
rect 8067 19708 8105 19742
rect 8139 19708 8177 19742
rect 8211 19708 8249 19742
rect 8283 19708 8321 19742
rect 8355 19708 8393 19742
rect 8427 19708 8465 19742
rect 8499 19708 8537 19742
rect 8571 19708 8609 19742
rect 8643 19708 8681 19742
rect 8715 19708 8753 19742
rect 8787 19708 8825 19742
rect 8859 19708 8897 19742
rect 8931 19708 8969 19742
rect 9003 19708 9041 19742
rect 9075 19708 9113 19742
rect 9147 19708 9185 19742
rect 9219 19708 9257 19742
rect 9291 19708 9329 19742
rect 9363 19708 9401 19742
rect 9435 19708 9473 19742
rect 9507 19708 9545 19742
rect 9579 19708 9617 19742
rect 9651 19708 9689 19742
rect 9723 19708 9761 19742
rect 9795 19708 9833 19742
rect 9867 19708 9905 19742
rect 9939 19708 9977 19742
rect 10011 19708 10049 19742
rect 10083 19708 10121 19742
rect 10155 19708 10193 19742
rect 10227 19708 10265 19742
rect 10299 19708 10337 19742
rect 10371 19708 10409 19742
rect 10443 19708 10481 19742
rect 10515 19708 10553 19742
rect 10587 19708 10625 19742
rect 10659 19708 10697 19742
rect 10731 19708 10769 19742
rect 10803 19708 10841 19742
rect 10875 19708 10913 19742
rect 10947 19708 10985 19742
rect 11019 19708 11057 19742
rect 11091 19708 11129 19742
rect 11163 19708 11201 19742
rect 11235 19708 11273 19742
rect 11307 19708 11345 19742
rect 11379 19708 11417 19742
rect 11451 19708 11489 19742
rect 11523 19708 11561 19742
rect 11595 19708 11633 19742
rect 11667 19708 11705 19742
rect 11739 19708 11777 19742
rect 11811 19708 11849 19742
rect 11883 19708 11921 19742
rect 11955 19708 11993 19742
rect 12027 19708 12065 19742
rect 12099 19708 12137 19742
rect 12171 19708 12209 19742
rect 12243 19708 12281 19742
rect 12315 19708 12353 19742
rect 12387 19708 12425 19742
rect 12459 19708 12497 19742
rect 12531 19708 12569 19742
rect 12603 19708 12641 19742
rect 12675 19708 12713 19742
rect 12747 19708 12785 19742
rect 12819 19708 12857 19742
rect 12891 19708 12929 19742
rect 12963 19708 12975 19742
rect 5033 19702 12975 19708
rect 13199 19745 13602 19896
rect 13199 19706 13490 19745
rect 13596 19706 13602 19745
rect 13199 19654 13200 19706
rect 13252 19654 13270 19706
rect 13322 19654 13340 19706
rect 13392 19654 13410 19706
rect 13462 19654 13480 19706
rect 13199 19642 13490 19654
rect 13596 19642 13602 19654
rect 4731 19614 4849 19626
tri 3794 17571 3828 17605 se
rect 3828 17571 4268 17605
tri 3771 17548 3794 17571 se
rect 3794 17548 4268 17571
tri 3768 17545 3771 17548 se
rect 3771 17545 4268 17548
tri 3754 17531 3768 17545 se
rect 3768 17531 4268 17545
tri 3735 17512 3754 17531 se
rect 3754 17512 4268 17531
rect 382 4572 423 4606
rect 457 4572 500 4606
rect 382 4529 500 4572
rect 382 4495 423 4529
rect 457 4495 500 4529
rect 382 4452 500 4495
rect 382 4418 423 4452
rect 457 4418 500 4452
rect 382 4375 500 4418
rect 382 4341 423 4375
rect 457 4341 500 4375
rect 382 4298 500 4341
rect 382 4264 423 4298
rect 457 4264 500 4298
rect 382 4220 500 4264
rect 382 4186 423 4220
rect 457 4186 500 4220
rect 382 4142 500 4186
rect 382 4108 423 4142
rect 457 4108 500 4142
rect 382 4096 500 4108
rect 560 17314 4268 17512
rect 4480 19578 4662 19590
rect 4480 19544 4486 19578
rect 4520 19544 4622 19578
rect 4656 19544 4662 19578
rect 4480 19505 4662 19544
rect 4480 19471 4486 19505
rect 4520 19471 4622 19505
rect 4656 19471 4662 19505
rect 4480 19432 4662 19471
rect 4480 19398 4486 19432
rect 4520 19398 4622 19432
rect 4656 19398 4662 19432
rect 4480 19359 4662 19398
rect 4480 19325 4486 19359
rect 4520 19325 4622 19359
rect 4656 19325 4662 19359
rect 4480 19286 4662 19325
rect 4480 19252 4486 19286
rect 4520 19252 4622 19286
rect 4656 19252 4662 19286
rect 4480 19213 4662 19252
rect 4480 19179 4486 19213
rect 4520 19179 4622 19213
rect 4656 19179 4662 19213
rect 4480 19140 4662 19179
rect 4480 19106 4486 19140
rect 4520 19106 4622 19140
rect 4656 19106 4662 19140
rect 4480 19067 4662 19106
rect 4480 19033 4486 19067
rect 4520 19033 4622 19067
rect 4656 19033 4662 19067
rect 4480 18994 4662 19033
rect 4480 18960 4486 18994
rect 4520 18960 4622 18994
rect 4656 18960 4662 18994
rect 4480 18921 4662 18960
rect 4480 18887 4486 18921
rect 4520 18887 4622 18921
rect 4656 18887 4662 18921
rect 4480 18848 4662 18887
rect 4480 18814 4486 18848
rect 4520 18814 4622 18848
rect 4656 18814 4662 18848
rect 4480 18775 4662 18814
rect 4480 18741 4486 18775
rect 4520 18741 4622 18775
rect 4656 18741 4662 18775
rect 4480 18702 4662 18741
rect 4480 18668 4486 18702
rect 4520 18668 4622 18702
rect 4656 18668 4662 18702
rect 4480 18629 4662 18668
rect 4480 18595 4486 18629
rect 4520 18595 4622 18629
rect 4656 18595 4662 18629
rect 4480 18556 4662 18595
rect 4480 18522 4486 18556
rect 4520 18522 4622 18556
rect 4656 18522 4662 18556
rect 4480 18483 4662 18522
rect 4480 18449 4486 18483
rect 4520 18449 4622 18483
rect 4656 18449 4662 18483
rect 4480 18410 4662 18449
rect 4480 18376 4486 18410
rect 4520 18376 4622 18410
rect 4656 18376 4662 18410
rect 4480 18337 4662 18376
rect 4480 18303 4486 18337
rect 4520 18303 4622 18337
rect 4656 18303 4662 18337
rect 4480 18264 4662 18303
rect 4480 18230 4486 18264
rect 4520 18230 4622 18264
rect 4656 18230 4662 18264
rect 4480 18191 4662 18230
rect 4480 18157 4486 18191
rect 4520 18157 4622 18191
rect 4656 18157 4662 18191
rect 4480 18118 4662 18157
rect 4480 18084 4486 18118
rect 4520 18084 4622 18118
rect 4656 18084 4662 18118
rect 4480 18045 4662 18084
rect 4480 18011 4486 18045
rect 4520 18011 4622 18045
rect 4656 18011 4662 18045
rect 4480 17972 4662 18011
rect 4480 17938 4486 17972
rect 4520 17938 4622 17972
rect 4656 17938 4662 17972
rect 4480 17899 4662 17938
rect 4480 17865 4486 17899
rect 4520 17865 4622 17899
rect 4656 17865 4662 17899
rect 4480 17826 4662 17865
rect 4480 17792 4486 17826
rect 4520 17792 4622 17826
rect 4656 17792 4662 17826
rect 4480 17753 4662 17792
rect 4480 17719 4486 17753
rect 4520 17719 4622 17753
rect 4656 17719 4662 17753
rect 4480 17679 4662 17719
rect 4480 17645 4486 17679
rect 4520 17645 4622 17679
rect 4656 17645 4662 17679
rect 4480 17605 4662 17645
rect 4480 17571 4486 17605
rect 4520 17571 4622 17605
rect 4656 17571 4662 17605
rect 4480 17531 4662 17571
rect 4480 17497 4486 17531
rect 4520 17497 4622 17531
rect 4656 17497 4662 17531
rect 4480 17457 4662 17497
rect 4480 17423 4486 17457
rect 4520 17423 4622 17457
rect 4656 17423 4662 17457
rect 4480 17383 4662 17423
rect 4480 17349 4486 17383
rect 4520 17349 4622 17383
rect 4656 17349 4662 17383
rect 560 17309 843 17314
tri 843 17309 848 17314 nw
rect 4480 17309 4662 17349
rect 560 17275 809 17309
tri 809 17275 843 17309 nw
rect 4480 17275 4486 17309
rect 4520 17275 4622 17309
rect 4656 17275 4662 17309
rect 560 17252 786 17275
tri 786 17252 809 17275 nw
rect 560 17249 783 17252
tri 783 17249 786 17252 nw
rect 560 17235 769 17249
tri 769 17235 783 17249 nw
rect 4480 17235 4662 17275
tri 481 3984 560 4063 se
rect 560 3984 760 17235
tri 760 17226 769 17235 nw
rect 4480 17201 4486 17235
rect 4520 17201 4622 17235
rect 4656 17201 4662 17235
rect 4480 17161 4662 17201
rect 4480 17127 4486 17161
rect 4520 17127 4622 17161
rect 4656 17127 4662 17161
rect 4480 17087 4662 17127
rect 4480 17053 4486 17087
rect 4520 17053 4622 17087
rect 4656 17053 4662 17087
rect 4480 17013 4662 17053
rect 4480 16979 4486 17013
rect 4520 16979 4622 17013
rect 4656 16979 4662 17013
rect 4480 16939 4662 16979
rect 814 16917 2372 16929
rect 814 16883 2184 16917
rect 2218 16883 2258 16917
rect 2292 16883 2332 16917
rect 2366 16883 2372 16917
rect 814 16798 2372 16883
rect 814 16764 2184 16798
rect 2218 16764 2258 16798
rect 2292 16764 2332 16798
rect 2366 16764 2372 16798
rect 814 16749 2372 16764
rect 3893 16917 4087 16929
rect 3893 16883 3899 16917
rect 3933 16883 3973 16917
rect 4007 16883 4047 16917
rect 4081 16883 4087 16917
rect 3893 16798 4087 16883
rect 3893 16764 3899 16798
rect 3933 16764 3973 16798
rect 4007 16764 4047 16798
rect 4081 16764 4087 16798
rect 814 16737 944 16749
tri 944 16737 956 16749 nw
rect 814 16717 924 16737
tri 924 16717 944 16737 nw
rect 814 4332 914 16717
tri 914 16707 924 16717 nw
tri 3881 16591 3893 16603 se
rect 3893 16591 4087 16764
tri 3866 16576 3881 16591 se
rect 3881 16576 4087 16591
tri 1057 16569 1064 16576 se
rect 1064 16569 4087 16576
tri 1033 16545 1057 16569 se
rect 1057 16545 4087 16569
tri 1023 16535 1033 16545 se
rect 1033 16535 4087 16545
tri 983 16495 1023 16535 se
rect 1023 16495 4087 16535
tri 952 16464 983 16495 se
rect 983 16464 4087 16495
rect 952 16382 4087 16464
rect 4480 16905 4486 16939
rect 4520 16905 4622 16939
rect 4656 16905 4662 16939
rect 4480 16865 4662 16905
rect 4480 16831 4486 16865
rect 4520 16831 4622 16865
rect 4656 16831 4662 16865
rect 4480 16791 4662 16831
rect 4480 16757 4486 16791
rect 4520 16757 4622 16791
rect 4656 16757 4662 16791
rect 4480 16717 4662 16757
rect 4480 16683 4486 16717
rect 4520 16683 4622 16717
rect 4656 16683 4662 16717
rect 4480 16657 4662 16683
rect 4480 16605 4481 16657
rect 4533 16605 4545 16657
rect 4597 16605 4609 16657
rect 4661 16605 4662 16657
rect 4480 16569 4662 16605
rect 4480 16545 4486 16569
rect 4520 16545 4622 16569
rect 4656 16545 4662 16569
rect 4731 19580 4737 19614
rect 4771 19580 4809 19614
rect 4843 19580 4849 19614
rect 4731 19540 4849 19580
rect 13199 19590 13200 19642
rect 13252 19590 13270 19642
rect 13322 19590 13340 19642
rect 13392 19590 13410 19642
rect 13462 19590 13480 19642
rect 13199 19578 13490 19590
rect 13596 19578 13602 19590
tri 13198 19540 13199 19541 se
rect 13199 19540 13200 19578
rect 4731 19506 4737 19540
rect 4771 19506 4809 19540
rect 4843 19506 4849 19540
rect 4731 19466 4849 19506
tri 13156 19498 13198 19540 se
rect 13198 19526 13200 19540
rect 13252 19526 13270 19578
rect 13322 19526 13340 19578
rect 13392 19526 13410 19578
rect 13462 19526 13480 19578
rect 13198 19514 13490 19526
rect 13596 19514 13602 19526
rect 13198 19498 13200 19514
rect 4731 19432 4737 19466
rect 4771 19432 4809 19466
rect 4843 19432 4849 19466
tri 13122 19464 13156 19498 se
rect 13156 19464 13200 19498
rect 4731 19392 4849 19432
tri 13080 19422 13122 19464 se
rect 13122 19462 13200 19464
rect 13252 19462 13270 19514
rect 13322 19462 13340 19514
rect 13392 19462 13410 19514
rect 13462 19462 13480 19514
rect 13122 19450 13490 19462
rect 13596 19450 13602 19462
rect 13122 19422 13200 19450
tri 13055 19397 13080 19422 se
rect 13080 19398 13200 19422
rect 13252 19398 13270 19450
rect 13322 19398 13340 19450
rect 13392 19398 13410 19450
rect 13462 19398 13480 19450
rect 13080 19397 13342 19398
rect 4731 19358 4737 19392
rect 4771 19358 4809 19392
rect 4843 19358 4849 19392
rect 4731 19318 4849 19358
rect 4731 19284 4737 19318
rect 4771 19284 4809 19318
rect 4843 19284 4849 19318
rect 4731 19244 4849 19284
rect 4731 19210 4737 19244
rect 4771 19210 4809 19244
rect 4843 19210 4849 19244
rect 4731 19170 4849 19210
rect 4731 19136 4737 19170
rect 4771 19136 4809 19170
rect 4843 19136 4849 19170
rect 4731 19096 4849 19136
rect 4731 19062 4737 19096
rect 4771 19062 4809 19096
rect 4843 19062 4849 19096
rect 4731 19022 4849 19062
rect 4731 18988 4737 19022
rect 4771 18988 4809 19022
rect 4843 18988 4849 19022
rect 4731 18948 4849 18988
rect 4731 18914 4737 18948
rect 4771 18914 4809 18948
rect 4843 18914 4849 18948
rect 4731 18874 4849 18914
rect 4731 18840 4737 18874
rect 4771 18840 4809 18874
rect 4843 18840 4849 18874
rect 4731 18801 4849 18840
rect 4731 18767 4737 18801
rect 4771 18767 4809 18801
rect 4843 18767 4849 18801
rect 4731 18728 4849 18767
rect 4731 18694 4737 18728
rect 4771 18694 4809 18728
rect 4843 18694 4849 18728
rect 4731 18655 4849 18694
rect 4731 18621 4737 18655
rect 4771 18621 4809 18655
rect 4843 18621 4849 18655
rect 4731 18582 4849 18621
rect 4731 18548 4737 18582
rect 4771 18548 4809 18582
rect 4843 18548 4849 18582
rect 4731 18509 4849 18548
rect 4731 18475 4737 18509
rect 4771 18475 4809 18509
rect 4843 18475 4849 18509
rect 4731 18436 4849 18475
rect 4731 18402 4737 18436
rect 4771 18402 4809 18436
rect 4843 18402 4849 18436
rect 4731 18363 4849 18402
rect 5056 19388 13342 19397
rect 13376 19388 13490 19398
rect 5056 19386 13490 19388
rect 13596 19386 13602 19398
rect 5056 19385 13200 19386
rect 5056 19351 5062 19385
rect 5096 19351 6718 19385
rect 6752 19351 8374 19385
rect 8408 19351 10030 19385
rect 10064 19351 11686 19385
rect 11720 19351 13200 19385
rect 5056 19334 13200 19351
rect 13252 19334 13270 19386
rect 13322 19334 13340 19386
rect 13392 19334 13410 19386
rect 13462 19334 13480 19386
rect 5056 19322 13342 19334
rect 13376 19322 13490 19334
rect 13596 19322 13602 19334
rect 5056 19310 13200 19322
rect 5056 19276 5062 19310
rect 5096 19276 6718 19310
rect 6752 19276 8374 19310
rect 8408 19276 10030 19310
rect 10064 19276 11686 19310
rect 11720 19276 13200 19310
rect 5056 19270 13200 19276
rect 13252 19270 13270 19322
rect 13322 19270 13340 19322
rect 13392 19270 13410 19322
rect 13462 19270 13480 19322
rect 5056 19258 13342 19270
rect 13376 19258 13490 19270
rect 13596 19258 13602 19270
rect 5056 19235 13200 19258
rect 5056 19201 5062 19235
rect 5096 19201 6718 19235
rect 6752 19201 8374 19235
rect 8408 19201 10030 19235
rect 10064 19201 11686 19235
rect 11720 19206 13200 19235
rect 13252 19206 13270 19258
rect 13322 19206 13340 19258
rect 13392 19206 13410 19258
rect 13462 19206 13480 19258
rect 11720 19201 13490 19206
rect 5056 19194 13490 19201
rect 13596 19194 13602 19206
rect 5056 19160 13200 19194
rect 5056 19126 5062 19160
rect 5096 19126 6718 19160
rect 6752 19126 8374 19160
rect 8408 19126 10030 19160
rect 10064 19126 11686 19160
rect 11720 19142 13200 19160
rect 13252 19142 13270 19194
rect 13322 19142 13340 19194
rect 13392 19142 13410 19194
rect 13462 19142 13480 19194
rect 11720 19130 13490 19142
rect 13596 19130 13602 19142
rect 11720 19126 13200 19130
rect 5056 19086 13200 19126
rect 5056 19052 5062 19086
rect 5096 19052 6718 19086
rect 6752 19052 8374 19086
rect 8408 19052 10030 19086
rect 10064 19052 11686 19086
rect 11720 19078 13200 19086
rect 13252 19078 13270 19130
rect 13322 19078 13340 19130
rect 13392 19078 13410 19130
rect 13462 19078 13480 19130
rect 11720 19066 13490 19078
rect 13596 19066 13602 19078
rect 11720 19052 13200 19066
rect 5056 19014 13200 19052
rect 13252 19014 13270 19066
rect 13322 19014 13340 19066
rect 13392 19014 13410 19066
rect 13462 19014 13480 19066
rect 5056 19012 13342 19014
rect 5056 18978 5062 19012
rect 5096 18978 6718 19012
rect 6752 18978 8374 19012
rect 8408 18978 10030 19012
rect 10064 18978 11686 19012
rect 11720 19008 13342 19012
rect 13376 19008 13490 19014
rect 11720 19002 13490 19008
rect 13596 19002 13602 19014
rect 11720 18978 13200 19002
rect 5056 18950 13200 18978
rect 13252 18950 13270 19002
rect 13322 18950 13340 19002
rect 13392 18950 13410 19002
rect 13462 18950 13480 19002
rect 5056 18938 13342 18950
rect 13376 18938 13490 18950
rect 13596 18938 13602 18950
rect 5056 18904 5062 18938
rect 5096 18904 6718 18938
rect 6752 18904 8374 18938
rect 8408 18904 10030 18938
rect 10064 18904 11686 18938
rect 11720 18904 13200 18938
rect 5056 18886 13200 18904
rect 13252 18886 13270 18938
rect 13322 18886 13340 18938
rect 13392 18886 13410 18938
rect 13462 18886 13480 18938
rect 5056 18874 13342 18886
rect 13376 18874 13490 18886
rect 13596 18874 13602 18886
rect 5056 18864 13200 18874
rect 5056 18830 5062 18864
rect 5096 18830 6718 18864
rect 6752 18830 8374 18864
rect 8408 18830 10030 18864
rect 10064 18830 11686 18864
rect 11720 18830 13200 18864
rect 5056 18822 13200 18830
rect 13252 18822 13270 18874
rect 13322 18822 13340 18874
rect 13392 18822 13410 18874
rect 13462 18822 13480 18874
rect 5056 18815 13490 18822
rect 5056 18810 13342 18815
rect 13376 18810 13490 18815
rect 13596 18810 13602 18822
rect 5056 18790 13200 18810
rect 5056 18756 5062 18790
rect 5096 18756 6718 18790
rect 6752 18756 8374 18790
rect 8408 18756 10030 18790
rect 10064 18756 11686 18790
rect 11720 18758 13200 18790
rect 13252 18758 13270 18810
rect 13322 18758 13340 18810
rect 13392 18758 13410 18810
rect 13462 18758 13480 18810
rect 11720 18756 13490 18758
rect 5056 18746 13490 18756
rect 13596 18746 13602 18758
rect 5056 18716 13200 18746
rect 5056 18682 5062 18716
rect 5096 18682 6718 18716
rect 6752 18682 8374 18716
rect 8408 18682 10030 18716
rect 10064 18682 11686 18716
rect 11720 18694 13200 18716
rect 13252 18694 13270 18746
rect 13322 18694 13340 18746
rect 13392 18694 13410 18746
rect 13462 18694 13480 18746
rect 11720 18682 13490 18694
rect 13596 18682 13602 18694
rect 5056 18642 13200 18682
rect 5056 18608 5062 18642
rect 5096 18608 6718 18642
rect 6752 18608 8374 18642
rect 8408 18608 10030 18642
rect 10064 18608 11686 18642
rect 11720 18630 13200 18642
rect 13252 18630 13270 18682
rect 13322 18630 13340 18682
rect 13392 18630 13410 18682
rect 13462 18630 13480 18682
rect 11720 18618 13490 18630
rect 13596 18618 13602 18630
rect 11720 18608 13200 18618
rect 5056 18568 13200 18608
rect 5056 18534 5062 18568
rect 5096 18534 6718 18568
rect 6752 18534 8374 18568
rect 8408 18534 10030 18568
rect 10064 18534 11686 18568
rect 11720 18566 13200 18568
rect 13252 18566 13270 18618
rect 13322 18566 13340 18618
rect 13392 18566 13410 18618
rect 13462 18566 13480 18618
rect 11720 18556 13342 18566
rect 13376 18556 13490 18566
rect 11720 18554 13490 18556
rect 13596 18554 13602 18566
rect 11720 18534 13200 18554
rect 5056 18502 13200 18534
rect 13252 18502 13270 18554
rect 13322 18502 13340 18554
rect 13392 18502 13410 18554
rect 13462 18502 13480 18554
rect 5056 18494 13342 18502
rect 5056 18460 5062 18494
rect 5096 18460 6718 18494
rect 6752 18460 8374 18494
rect 8408 18460 10030 18494
rect 10064 18460 11686 18494
rect 11720 18490 13342 18494
rect 13376 18490 13490 18502
rect 13596 18490 13602 18502
rect 11720 18460 13200 18490
rect 5056 18438 13200 18460
rect 13252 18438 13270 18490
rect 13322 18438 13340 18490
rect 13392 18438 13410 18490
rect 13462 18438 13480 18490
rect 5056 18426 13342 18438
rect 13376 18426 13490 18438
rect 13596 18426 13602 18438
rect 5056 18420 13200 18426
rect 5056 18386 5062 18420
rect 5096 18386 6718 18420
rect 6752 18386 8374 18420
rect 8408 18386 10030 18420
rect 10064 18386 11686 18420
rect 11720 18386 13200 18420
rect 5056 18374 13200 18386
rect 13252 18374 13270 18426
rect 13322 18374 13340 18426
rect 13392 18374 13410 18426
rect 13462 18374 13480 18426
tri 12970 18365 12979 18374 ne
rect 12979 18365 13490 18374
rect 4731 18329 4737 18363
rect 4771 18329 4809 18363
rect 4843 18329 4849 18363
tri 12979 18331 13013 18365 ne
rect 13013 18362 13342 18365
rect 13376 18362 13490 18365
rect 13596 18362 13602 18374
rect 13013 18331 13200 18362
rect 4731 18290 4849 18329
tri 13013 18290 13054 18331 ne
rect 13054 18310 13200 18331
rect 13252 18310 13270 18362
rect 13322 18310 13340 18362
rect 13392 18310 13410 18362
rect 13462 18310 13480 18362
rect 13054 18298 13490 18310
rect 13596 18298 13602 18310
rect 13054 18290 13200 18298
rect 4731 18256 4737 18290
rect 4771 18256 4809 18290
rect 4843 18256 4849 18290
tri 13054 18256 13088 18290 ne
rect 13088 18256 13200 18290
rect 4731 17915 4849 18256
tri 13088 18223 13121 18256 ne
rect 13121 18246 13200 18256
rect 13252 18246 13270 18298
rect 13322 18246 13340 18298
rect 13392 18246 13410 18298
rect 13462 18246 13480 18298
rect 13121 18234 13490 18246
rect 13596 18234 13602 18246
rect 13121 18182 13200 18234
rect 13252 18182 13270 18234
rect 13322 18182 13340 18234
rect 13392 18182 13410 18234
rect 13462 18182 13480 18234
rect 13121 18170 13490 18182
rect 13596 18170 13602 18182
rect 13121 18118 13200 18170
rect 13252 18118 13270 18170
rect 13322 18118 13340 18170
rect 13392 18118 13410 18170
rect 13462 18118 13480 18170
rect 13121 18106 13490 18118
rect 13596 18106 13602 18118
rect 4911 18003 4917 18055
rect 4969 18003 4981 18055
rect 5033 18049 5039 18055
tri 5039 18049 5045 18055 sw
rect 13121 18054 13200 18106
rect 13252 18054 13270 18106
rect 13322 18054 13340 18106
rect 13392 18054 13410 18106
rect 13462 18054 13480 18106
rect 5033 18043 12975 18049
rect 5033 18009 5069 18043
rect 5103 18009 5142 18043
rect 5176 18009 5215 18043
rect 5249 18009 5288 18043
rect 5322 18009 5361 18043
rect 5395 18009 5434 18043
rect 5468 18009 5507 18043
rect 5541 18009 5580 18043
rect 5614 18009 5653 18043
rect 5687 18009 5726 18043
rect 5760 18009 5799 18043
rect 5833 18009 5872 18043
rect 5906 18009 5945 18043
rect 5979 18009 6017 18043
rect 6051 18009 6089 18043
rect 6123 18009 6161 18043
rect 6195 18009 6233 18043
rect 6267 18009 6305 18043
rect 6339 18009 6377 18043
rect 6411 18009 6449 18043
rect 6483 18009 6521 18043
rect 6555 18009 6593 18043
rect 6627 18009 6665 18043
rect 6699 18009 6737 18043
rect 6771 18009 6809 18043
rect 6843 18009 6881 18043
rect 6915 18009 6953 18043
rect 6987 18009 7025 18043
rect 7059 18009 7097 18043
rect 7131 18009 7169 18043
rect 7203 18009 7241 18043
rect 7275 18009 7313 18043
rect 7347 18009 7385 18043
rect 7419 18009 7457 18043
rect 7491 18009 7529 18043
rect 7563 18009 7601 18043
rect 7635 18009 7673 18043
rect 7707 18009 7745 18043
rect 7779 18009 7817 18043
rect 7851 18009 7889 18043
rect 7923 18009 7961 18043
rect 7995 18009 8033 18043
rect 8067 18009 8105 18043
rect 8139 18009 8177 18043
rect 8211 18009 8249 18043
rect 8283 18009 8321 18043
rect 8355 18009 8393 18043
rect 8427 18009 8465 18043
rect 8499 18009 8537 18043
rect 8571 18009 8609 18043
rect 8643 18009 8681 18043
rect 8715 18009 8753 18043
rect 8787 18009 8825 18043
rect 8859 18009 8897 18043
rect 8931 18009 8969 18043
rect 9003 18009 9041 18043
rect 9075 18009 9113 18043
rect 9147 18009 9185 18043
rect 9219 18009 9257 18043
rect 9291 18009 9329 18043
rect 9363 18009 9401 18043
rect 9435 18009 9473 18043
rect 9507 18009 9545 18043
rect 9579 18009 9617 18043
rect 9651 18009 9689 18043
rect 9723 18009 9761 18043
rect 9795 18009 9833 18043
rect 9867 18009 9905 18043
rect 9939 18009 9977 18043
rect 10011 18009 10049 18043
rect 10083 18009 10121 18043
rect 10155 18009 10193 18043
rect 10227 18009 10265 18043
rect 10299 18009 10337 18043
rect 10371 18009 10409 18043
rect 10443 18009 10481 18043
rect 10515 18009 10553 18043
rect 10587 18009 10625 18043
rect 10659 18009 10697 18043
rect 10731 18009 10769 18043
rect 10803 18009 10841 18043
rect 10875 18009 10913 18043
rect 10947 18009 10985 18043
rect 11019 18009 11057 18043
rect 11091 18009 11129 18043
rect 11163 18009 11201 18043
rect 11235 18009 11273 18043
rect 11307 18009 11345 18043
rect 11379 18009 11417 18043
rect 11451 18009 11489 18043
rect 11523 18009 11561 18043
rect 11595 18009 11633 18043
rect 11667 18009 11705 18043
rect 11739 18009 11777 18043
rect 11811 18009 11849 18043
rect 11883 18009 11921 18043
rect 11955 18009 11993 18043
rect 12027 18009 12065 18043
rect 12099 18009 12137 18043
rect 12171 18009 12209 18043
rect 12243 18009 12281 18043
rect 12315 18009 12353 18043
rect 12387 18009 12425 18043
rect 12459 18009 12497 18043
rect 12531 18009 12569 18043
rect 12603 18009 12641 18043
rect 12675 18009 12713 18043
rect 12747 18009 12785 18043
rect 12819 18009 12857 18043
rect 12891 18009 12929 18043
rect 12963 18009 12975 18043
rect 5033 18003 12975 18009
rect 13121 18042 13490 18054
rect 13596 18042 13602 18054
rect 13121 17990 13200 18042
rect 13252 17990 13270 18042
rect 13322 17990 13340 18042
rect 13392 17990 13410 18042
rect 13462 17990 13480 18042
rect 13121 17978 13490 17990
rect 13596 17978 13602 17990
rect 4731 17881 4737 17915
rect 4771 17881 4809 17915
rect 4843 17881 4849 17915
rect 4731 17841 4849 17881
tri 13035 17875 13121 17961 se
rect 13121 17926 13200 17978
rect 13252 17926 13270 17978
rect 13322 17926 13340 17978
rect 13392 17926 13410 17978
rect 13462 17926 13480 17978
rect 13121 17914 13490 17926
rect 13596 17914 13602 17926
rect 13121 17875 13200 17914
tri 13001 17841 13035 17875 se
rect 13035 17862 13200 17875
rect 13252 17862 13270 17914
rect 13322 17862 13340 17914
rect 13392 17862 13410 17914
rect 13462 17862 13480 17914
rect 13035 17850 13342 17862
rect 13376 17850 13490 17862
rect 13596 17850 13602 17862
rect 13035 17841 13200 17850
rect 4731 17807 4737 17841
rect 4771 17807 4809 17841
rect 4843 17807 4849 17841
tri 12976 17816 13001 17841 se
rect 13001 17816 13200 17841
rect 4731 17767 4849 17807
rect 4731 17733 4737 17767
rect 4771 17733 4809 17767
rect 4843 17733 4849 17767
rect 4731 17693 4849 17733
rect 4731 17659 4737 17693
rect 4771 17659 4809 17693
rect 4843 17659 4849 17693
rect 4731 17619 4849 17659
rect 4731 17585 4737 17619
rect 4771 17585 4809 17619
rect 4843 17585 4849 17619
rect 4731 17545 4849 17585
rect 4731 17511 4737 17545
rect 4771 17511 4809 17545
rect 4843 17511 4849 17545
rect 4731 17471 4849 17511
rect 4731 17437 4737 17471
rect 4771 17437 4809 17471
rect 4843 17437 4849 17471
rect 4731 17397 4849 17437
rect 4731 17363 4737 17397
rect 4771 17363 4809 17397
rect 4843 17363 4849 17397
rect 4731 17323 4849 17363
rect 4731 17289 4737 17323
rect 4771 17289 4809 17323
rect 4843 17289 4849 17323
rect 4731 17249 4849 17289
rect 4731 17215 4737 17249
rect 4771 17215 4809 17249
rect 4843 17215 4849 17249
rect 4731 17175 4849 17215
rect 4731 17141 4737 17175
rect 4771 17141 4809 17175
rect 4843 17141 4849 17175
rect 4731 17102 4849 17141
rect 4731 17068 4737 17102
rect 4771 17068 4809 17102
rect 4843 17068 4849 17102
rect 4731 17029 4849 17068
rect 4731 16995 4737 17029
rect 4771 16995 4809 17029
rect 4843 16995 4849 17029
rect 4731 16956 4849 16995
rect 4731 16922 4737 16956
rect 4771 16922 4809 16956
rect 4843 16922 4849 16956
rect 4731 16883 4849 16922
rect 4731 16849 4737 16883
rect 4771 16849 4809 16883
rect 4843 16849 4849 16883
rect 4731 16810 4849 16849
rect 4731 16809 4737 16810
rect 4771 16809 4809 16810
rect 4843 16809 4849 16810
rect 4783 16757 4797 16809
rect 4731 16737 4849 16757
rect 4731 16706 4737 16737
rect 4771 16706 4809 16737
rect 4843 16706 4849 16737
rect 4783 16654 4797 16706
rect 4731 16630 4737 16654
rect 4771 16630 4809 16654
rect 4843 16630 4849 16654
rect 4731 16603 4849 16630
rect 4783 16551 4797 16603
rect 5056 17804 13200 17816
rect 5056 17770 5062 17804
rect 5096 17770 6718 17804
rect 6752 17770 8374 17804
rect 8408 17770 10030 17804
rect 10064 17770 11686 17804
rect 11720 17798 13200 17804
rect 13252 17798 13270 17850
rect 13322 17798 13340 17850
rect 13392 17798 13410 17850
rect 13462 17798 13480 17850
rect 11720 17786 13342 17798
rect 13376 17786 13490 17798
rect 13596 17786 13602 17798
rect 11720 17770 13200 17786
rect 5056 17734 13200 17770
rect 13252 17734 13270 17786
rect 13322 17734 13340 17786
rect 13392 17734 13410 17786
rect 13462 17734 13480 17786
rect 5056 17730 13490 17734
rect 5056 17696 5062 17730
rect 5096 17696 6718 17730
rect 6752 17696 8374 17730
rect 8408 17696 10030 17730
rect 10064 17696 11686 17730
rect 11720 17725 13490 17730
rect 11720 17722 13342 17725
rect 13376 17722 13490 17725
rect 13596 17722 13602 17734
rect 11720 17696 13200 17722
rect 5056 17670 13200 17696
rect 13252 17670 13270 17722
rect 13322 17670 13340 17722
rect 13392 17670 13410 17722
rect 13462 17670 13480 17722
rect 5056 17658 13490 17670
rect 13596 17658 13602 17670
rect 5056 17656 13200 17658
rect 5056 17622 5062 17656
rect 5096 17622 6718 17656
rect 6752 17622 8374 17656
rect 8408 17622 10030 17656
rect 10064 17622 11686 17656
rect 11720 17622 13200 17656
rect 5056 17606 13200 17622
rect 13252 17606 13270 17658
rect 13322 17606 13340 17658
rect 13392 17606 13410 17658
rect 13462 17606 13480 17658
rect 5056 17594 13490 17606
rect 13596 17594 13602 17606
rect 5056 17582 13200 17594
rect 5056 17548 5062 17582
rect 5096 17548 6718 17582
rect 6752 17548 8374 17582
rect 8408 17548 10030 17582
rect 10064 17548 11686 17582
rect 11720 17548 13200 17582
rect 5056 17542 13200 17548
rect 13252 17542 13270 17594
rect 13322 17542 13340 17594
rect 13392 17542 13410 17594
rect 13462 17542 13480 17594
rect 5056 17541 13342 17542
rect 13376 17541 13490 17542
rect 5056 17530 13490 17541
rect 13596 17530 13602 17542
rect 5056 17508 13200 17530
rect 5056 17474 5062 17508
rect 5096 17474 6718 17508
rect 6752 17474 8374 17508
rect 8408 17474 10030 17508
rect 10064 17474 11686 17508
rect 11720 17478 13200 17508
rect 13252 17478 13270 17530
rect 13322 17478 13340 17530
rect 13392 17478 13410 17530
rect 13462 17478 13480 17530
rect 11720 17474 13342 17478
rect 5056 17466 13342 17474
rect 13376 17466 13490 17478
rect 13596 17466 13602 17478
rect 5056 17434 13200 17466
rect 5056 17400 5062 17434
rect 5096 17400 6718 17434
rect 6752 17400 8374 17434
rect 8408 17400 10030 17434
rect 10064 17400 11686 17434
rect 11720 17414 13200 17434
rect 13252 17414 13270 17466
rect 13322 17414 13340 17466
rect 13392 17414 13410 17466
rect 13462 17414 13480 17466
rect 11720 17402 13342 17414
rect 13376 17402 13490 17414
rect 13596 17402 13602 17414
rect 11720 17400 13200 17402
rect 5056 17360 13200 17400
rect 5056 17326 5062 17360
rect 5096 17326 6718 17360
rect 6752 17326 8374 17360
rect 8408 17326 10030 17360
rect 10064 17326 11686 17360
rect 11720 17350 13200 17360
rect 13252 17350 13270 17402
rect 13322 17350 13340 17402
rect 13392 17350 13410 17402
rect 13462 17350 13480 17402
rect 11720 17338 13342 17350
rect 13376 17338 13490 17350
rect 13596 17338 13602 17350
rect 11720 17326 13200 17338
rect 5056 17286 13200 17326
rect 13252 17286 13270 17338
rect 13322 17286 13340 17338
rect 13392 17286 13410 17338
rect 13462 17286 13480 17338
rect 5056 17252 5062 17286
rect 5096 17252 6718 17286
rect 6752 17252 8374 17286
rect 8408 17252 10030 17286
rect 10064 17252 11686 17286
rect 11720 17275 13490 17286
rect 11720 17274 13342 17275
rect 13376 17274 13490 17275
rect 13596 17274 13602 17286
rect 11720 17252 13200 17274
rect 5056 17222 13200 17252
rect 13252 17222 13270 17274
rect 13322 17222 13340 17274
rect 13392 17222 13410 17274
rect 13462 17222 13480 17274
rect 5056 17212 13490 17222
rect 5056 17178 5062 17212
rect 5096 17178 6718 17212
rect 6752 17178 8374 17212
rect 8408 17178 10030 17212
rect 10064 17178 11686 17212
rect 11720 17210 13490 17212
rect 13596 17210 13602 17222
rect 11720 17178 13200 17210
rect 5056 17158 13200 17178
rect 13252 17158 13270 17210
rect 13322 17158 13340 17210
rect 13392 17158 13410 17210
rect 13462 17158 13480 17210
rect 5056 17146 13490 17158
rect 13596 17146 13602 17158
rect 5056 17138 13200 17146
rect 5056 17104 5062 17138
rect 5096 17104 6718 17138
rect 6752 17104 8374 17138
rect 8408 17104 10030 17138
rect 10064 17104 11686 17138
rect 11720 17104 13200 17138
rect 5056 17094 13200 17104
rect 13252 17094 13270 17146
rect 13322 17094 13340 17146
rect 13392 17094 13410 17146
rect 13462 17094 13480 17146
rect 5056 17089 13342 17094
rect 13376 17089 13490 17094
rect 5056 17082 13490 17089
rect 13596 17082 13602 17094
rect 5056 17064 13200 17082
rect 5056 17030 5062 17064
rect 5096 17030 6718 17064
rect 6752 17030 8374 17064
rect 8408 17030 10030 17064
rect 10064 17030 11686 17064
rect 11720 17030 13200 17064
rect 13252 17030 13270 17082
rect 13322 17030 13340 17082
rect 13392 17030 13410 17082
rect 13462 17030 13480 17082
rect 5056 17018 13342 17030
rect 13376 17018 13490 17030
rect 13596 17018 13602 17030
rect 5056 16990 13200 17018
rect 5056 16956 5062 16990
rect 5096 16956 6718 16990
rect 6752 16956 8374 16990
rect 8408 16956 10030 16990
rect 10064 16956 11686 16990
rect 11720 16966 13200 16990
rect 13252 16966 13270 17018
rect 13322 16966 13340 17018
rect 13392 16966 13410 17018
rect 13462 16966 13480 17018
rect 11720 16956 13342 16966
rect 5056 16954 13342 16956
rect 13376 16954 13490 16966
rect 13596 16954 13602 16966
rect 5056 16916 13200 16954
rect 5056 16882 5062 16916
rect 5096 16882 6718 16916
rect 6752 16882 8374 16916
rect 8408 16882 10030 16916
rect 10064 16882 11686 16916
rect 11720 16902 13200 16916
rect 13252 16902 13270 16954
rect 13322 16902 13340 16954
rect 13392 16902 13410 16954
rect 13462 16902 13480 16954
rect 11720 16895 13490 16902
rect 11720 16890 13342 16895
rect 13376 16890 13490 16895
rect 13596 16890 13602 16902
rect 11720 16882 13200 16890
rect 5056 16842 13200 16882
rect 5056 16808 5062 16842
rect 5096 16808 6718 16842
rect 6752 16808 8374 16842
rect 8408 16808 10030 16842
rect 10064 16808 11686 16842
rect 11720 16838 13200 16842
rect 13252 16838 13270 16890
rect 13322 16838 13340 16890
rect 13392 16838 13410 16890
rect 13462 16838 13480 16890
rect 11720 16826 13490 16838
rect 13596 16826 13602 16838
rect 11720 16808 13200 16826
rect 5056 16774 13200 16808
rect 13252 16774 13270 16826
rect 13322 16774 13340 16826
rect 13392 16774 13410 16826
rect 13462 16774 13480 16826
rect 5056 16767 13490 16774
rect 5056 16733 5062 16767
rect 5096 16733 6718 16767
rect 6752 16733 8374 16767
rect 8408 16733 10030 16767
rect 10064 16733 11686 16767
rect 11720 16762 13490 16767
rect 13596 16762 13602 16774
rect 11720 16733 13200 16762
rect 5056 16710 13200 16733
rect 13252 16710 13270 16762
rect 13322 16710 13340 16762
rect 13392 16710 13410 16762
rect 13462 16710 13480 16762
rect 5056 16709 13342 16710
rect 13376 16709 13490 16710
rect 5056 16698 13490 16709
rect 13596 16698 13602 16710
rect 5056 16692 13200 16698
rect 5056 16658 5062 16692
rect 5096 16658 6718 16692
rect 6752 16658 8374 16692
rect 8408 16658 10030 16692
rect 10064 16658 11686 16692
rect 11720 16658 13200 16692
rect 5056 16646 13200 16658
rect 13252 16646 13270 16698
rect 13322 16646 13340 16698
rect 13392 16646 13410 16698
rect 13462 16646 13480 16698
rect 5056 16634 13342 16646
rect 13376 16634 13490 16646
rect 13596 16634 13602 16646
rect 5056 16617 13200 16634
rect 5056 16583 5062 16617
rect 5096 16583 6718 16617
rect 6752 16583 8374 16617
rect 8408 16583 10030 16617
rect 10064 16583 11686 16617
rect 11720 16583 13200 16617
rect 5056 16582 13200 16583
rect 13252 16582 13270 16634
rect 13322 16582 13340 16634
rect 13392 16582 13410 16634
rect 13462 16582 13480 16634
rect 5056 16571 13342 16582
tri 12978 16557 12992 16571 ne
rect 12992 16570 13342 16571
rect 13376 16570 13490 16582
rect 13596 16570 13602 16582
rect 12992 16557 13200 16570
rect 4731 16545 4849 16551
tri 12992 16545 13004 16557 ne
rect 13004 16545 13200 16557
rect 4480 16493 4481 16545
rect 4533 16493 4545 16545
rect 4597 16493 4609 16545
rect 4661 16493 4662 16545
rect 4480 16461 4486 16493
rect 4520 16461 4622 16493
rect 4656 16461 4662 16493
rect 4480 16433 4662 16461
rect 952 4602 1248 16382
tri 1248 16353 1277 16382 nw
rect 4480 16381 4481 16433
rect 4533 16381 4545 16433
rect 4597 16381 4609 16433
rect 4661 16381 4662 16433
tri 13004 16428 13121 16545 ne
rect 13121 16518 13200 16545
rect 13252 16518 13270 16570
rect 13322 16518 13340 16570
rect 13392 16518 13410 16570
rect 13462 16518 13480 16570
rect 13121 16506 13490 16518
rect 13596 16506 13602 16518
rect 13121 16454 13200 16506
rect 13252 16454 13270 16506
rect 13322 16454 13340 16506
rect 13392 16454 13410 16506
rect 13462 16454 13480 16506
rect 13121 16442 13490 16454
rect 13596 16442 13602 16454
rect 4480 16375 4662 16381
rect 13121 16390 13200 16442
rect 13252 16390 13270 16442
rect 13322 16390 13340 16442
rect 13392 16390 13410 16442
rect 13462 16390 13480 16442
rect 13121 16378 13490 16390
rect 13596 16378 13602 16390
rect 13121 16326 13200 16378
rect 13252 16326 13270 16378
rect 13322 16326 13340 16378
rect 13392 16326 13410 16378
rect 13462 16326 13480 16378
rect 13121 16314 13490 16326
rect 13596 16314 13602 16326
rect 952 4568 995 4602
rect 1029 4568 1099 4602
rect 1133 4568 1202 4602
rect 1236 4568 1248 4602
rect 952 4492 1248 4568
rect 952 4485 995 4492
tri 952 4458 979 4485 ne
rect 979 4458 995 4485
rect 1029 4458 1099 4492
rect 1133 4458 1202 4492
rect 1236 4458 1248 4492
tri 979 4454 983 4458 ne
rect 983 4452 1248 4458
tri 985 4443 994 4452 ne
rect 994 4443 1248 4452
rect 1287 16271 13000 16280
rect 1287 16219 4917 16271
rect 4969 16219 4981 16271
rect 5033 16243 13000 16271
rect 5033 16219 5069 16243
rect 1287 16209 4923 16219
rect 4957 16209 4996 16219
rect 5030 16209 5069 16219
rect 5103 16209 5142 16243
rect 5176 16209 5215 16243
rect 5249 16209 5288 16243
rect 5322 16209 5361 16243
rect 5395 16209 5434 16243
rect 5468 16209 5507 16243
rect 5541 16209 5580 16243
rect 5614 16209 5653 16243
rect 5687 16209 5726 16243
rect 5760 16209 5799 16243
rect 5833 16209 5872 16243
rect 5906 16209 5945 16243
rect 5979 16209 6017 16243
rect 6051 16209 6089 16243
rect 6123 16209 6161 16243
rect 6195 16209 6233 16243
rect 6267 16209 6305 16243
rect 6339 16209 6377 16243
rect 6411 16209 6449 16243
rect 6483 16209 6521 16243
rect 6555 16209 6593 16243
rect 6627 16209 6665 16243
rect 6699 16209 6737 16243
rect 6771 16209 6809 16243
rect 6843 16209 6881 16243
rect 6915 16209 6953 16243
rect 6987 16209 7025 16243
rect 7059 16209 7097 16243
rect 7131 16209 7169 16243
rect 7203 16209 7241 16243
rect 7275 16209 7313 16243
rect 7347 16209 7385 16243
rect 7419 16209 7457 16243
rect 7491 16209 7529 16243
rect 7563 16209 7601 16243
rect 7635 16209 7673 16243
rect 7707 16209 7745 16243
rect 7779 16209 7817 16243
rect 7851 16209 7889 16243
rect 7923 16209 7961 16243
rect 7995 16209 8033 16243
rect 8067 16209 8105 16243
rect 8139 16209 8177 16243
rect 8211 16209 8249 16243
rect 8283 16209 8321 16243
rect 8355 16209 8393 16243
rect 8427 16209 8465 16243
rect 8499 16209 8537 16243
rect 8571 16209 8609 16243
rect 8643 16209 8681 16243
rect 8715 16209 8753 16243
rect 8787 16209 8825 16243
rect 8859 16209 8897 16243
rect 8931 16209 8969 16243
rect 9003 16209 9041 16243
rect 9075 16209 9113 16243
rect 9147 16209 9185 16243
rect 9219 16209 9257 16243
rect 9291 16209 9329 16243
rect 9363 16209 9401 16243
rect 9435 16209 9473 16243
rect 9507 16209 9545 16243
rect 9579 16209 9617 16243
rect 9651 16209 9689 16243
rect 9723 16209 9761 16243
rect 9795 16209 9833 16243
rect 9867 16209 9905 16243
rect 9939 16209 9977 16243
rect 10011 16209 10049 16243
rect 10083 16209 10121 16243
rect 10155 16209 10193 16243
rect 10227 16209 10265 16243
rect 10299 16209 10337 16243
rect 10371 16209 10409 16243
rect 10443 16209 10481 16243
rect 10515 16209 10553 16243
rect 10587 16209 10625 16243
rect 10659 16209 10697 16243
rect 10731 16209 10769 16243
rect 10803 16209 10841 16243
rect 10875 16209 10913 16243
rect 10947 16209 10985 16243
rect 11019 16209 11057 16243
rect 11091 16209 11129 16243
rect 11163 16209 11201 16243
rect 11235 16209 11273 16243
rect 11307 16209 11345 16243
rect 11379 16209 11417 16243
rect 11451 16209 11489 16243
rect 11523 16209 11561 16243
rect 11595 16209 11633 16243
rect 11667 16209 11705 16243
rect 11739 16209 11777 16243
rect 11811 16209 11849 16243
rect 11883 16209 11921 16243
rect 11955 16209 11993 16243
rect 12027 16209 12065 16243
rect 12099 16209 12137 16243
rect 12171 16209 12209 16243
rect 12243 16209 12281 16243
rect 12315 16209 12353 16243
rect 12387 16209 12425 16243
rect 12459 16209 12497 16243
rect 12531 16209 12569 16243
rect 12603 16209 12641 16243
rect 12675 16209 12713 16243
rect 12747 16209 12785 16243
rect 12819 16209 12857 16243
rect 12891 16209 12929 16243
rect 12963 16209 13000 16243
rect 13121 16262 13200 16314
rect 13252 16262 13270 16314
rect 13322 16262 13340 16314
rect 13392 16262 13410 16314
rect 13462 16262 13480 16314
rect 13121 16250 13490 16262
rect 13596 16250 13602 16262
rect 1287 16203 13000 16209
tri 13096 16203 13121 16228 se
rect 13121 16203 13200 16250
rect 1287 4416 1417 16203
tri 1417 16174 1446 16203 nw
tri 13067 16174 13096 16203 se
rect 13096 16198 13200 16203
rect 13252 16198 13270 16250
rect 13322 16198 13340 16250
rect 13392 16198 13410 16250
rect 13462 16198 13480 16250
rect 13096 16186 13490 16198
rect 13596 16186 13602 16198
rect 13096 16174 13200 16186
tri 13025 16132 13067 16174 se
rect 13067 16134 13200 16174
rect 13252 16134 13270 16186
rect 13322 16134 13340 16186
rect 13392 16134 13410 16186
rect 13462 16134 13480 16186
rect 13067 16132 13490 16134
rect 1938 16100 2056 16132
tri 13000 16107 13025 16132 se
rect 13025 16122 13490 16132
rect 13596 16122 13602 16134
rect 13025 16107 13200 16122
rect 1938 15922 1944 16100
rect 2050 15922 2056 16100
tri 12966 16073 13000 16107 se
rect 13000 16073 13200 16107
tri 12965 16072 12966 16073 se
rect 12966 16072 13200 16073
rect 1938 15883 2056 15922
rect 1938 15849 1944 15883
rect 1978 15849 2016 15883
rect 2050 15849 2056 15883
rect 1938 15810 2056 15849
rect 1938 15776 1944 15810
rect 1978 15776 2016 15810
rect 2050 15776 2056 15810
rect 1938 15737 2056 15776
rect 1938 15703 1944 15737
rect 1978 15703 2016 15737
rect 2050 15703 2056 15737
rect 1938 15664 2056 15703
rect 1938 15630 1944 15664
rect 1978 15630 2016 15664
rect 2050 15630 2056 15664
rect 1938 15591 2056 15630
rect 1938 15557 1944 15591
rect 1978 15557 2016 15591
rect 2050 15557 2056 15591
rect 1938 15518 2056 15557
rect 1938 15484 1944 15518
rect 1978 15484 2016 15518
rect 2050 15484 2056 15518
rect 1938 15445 2056 15484
rect 1938 15411 1944 15445
rect 1978 15411 2016 15445
rect 2050 15411 2056 15445
rect 1938 15372 2056 15411
rect 1938 15338 1944 15372
rect 1978 15338 2016 15372
rect 2050 15338 2056 15372
rect 1938 15306 2056 15338
rect 2274 16070 13200 16072
rect 13252 16070 13270 16122
rect 13322 16070 13340 16122
rect 13392 16070 13410 16122
rect 13462 16070 13480 16122
rect 2274 16066 13490 16070
rect 2274 16060 4481 16066
rect 2274 16040 2550 16060
rect 2274 16006 2280 16040
rect 2314 16006 2404 16040
rect 2438 16026 2550 16040
rect 2584 16026 3406 16060
rect 3440 16026 4481 16060
rect 2438 16014 4481 16026
rect 4533 16014 4545 16066
rect 4597 16014 4609 16066
rect 4661 16060 13490 16066
rect 4661 16026 5062 16060
rect 5096 16026 6718 16060
rect 6752 16026 8374 16060
rect 8408 16026 10030 16060
rect 10064 16026 11686 16060
rect 11720 16058 13490 16060
rect 13596 16058 13602 16070
rect 11720 16026 13200 16058
rect 4661 16014 13200 16026
rect 2438 16006 13200 16014
rect 13252 16006 13270 16058
rect 13322 16006 13340 16058
rect 13392 16006 13410 16058
rect 13462 16006 13480 16058
rect 2274 15996 13342 16006
rect 13376 15996 13490 16006
rect 2274 15994 13490 15996
rect 13596 15994 13602 16006
rect 2274 15987 13200 15994
rect 2274 15965 2550 15987
rect 2274 15931 2280 15965
rect 2314 15931 2404 15965
rect 2438 15953 2550 15965
rect 2584 15953 3406 15987
rect 3440 15953 5062 15987
rect 5096 15953 6718 15987
rect 6752 15953 8374 15987
rect 8408 15953 10030 15987
rect 10064 15953 11686 15987
rect 11720 15953 13200 15987
rect 2438 15942 13200 15953
rect 13252 15942 13270 15994
rect 13322 15942 13340 15994
rect 13392 15942 13410 15994
rect 13462 15942 13480 15994
rect 2438 15931 13342 15942
rect 2274 15930 13342 15931
rect 13376 15930 13490 15942
rect 13596 15930 13602 15942
rect 2274 15922 13200 15930
rect 2274 15914 4481 15922
rect 2274 15890 2550 15914
rect 2274 15856 2280 15890
rect 2314 15856 2404 15890
rect 2438 15880 2550 15890
rect 2584 15880 3406 15914
rect 3440 15880 4481 15914
rect 2438 15870 4481 15880
rect 4533 15870 4545 15922
rect 4597 15870 4609 15922
rect 4661 15914 13200 15922
rect 4661 15880 5062 15914
rect 5096 15880 6718 15914
rect 6752 15880 8374 15914
rect 8408 15880 10030 15914
rect 10064 15880 11686 15914
rect 11720 15880 13200 15914
rect 4661 15878 13200 15880
rect 13252 15878 13270 15930
rect 13322 15878 13340 15930
rect 13392 15878 13410 15930
rect 13462 15878 13480 15930
rect 4661 15876 13490 15878
rect 4661 15870 13342 15876
rect 2438 15866 13342 15870
rect 13376 15866 13490 15876
rect 13596 15866 13602 15878
rect 2438 15856 13200 15866
rect 2274 15841 13200 15856
rect 2274 15815 2550 15841
rect 2274 15781 2280 15815
rect 2314 15781 2404 15815
rect 2438 15807 2550 15815
rect 2584 15807 3406 15841
rect 3440 15807 5062 15841
rect 5096 15807 6718 15841
rect 6752 15807 8374 15841
rect 8408 15807 10030 15841
rect 10064 15807 11686 15841
rect 11720 15814 13200 15841
rect 13252 15814 13270 15866
rect 13322 15814 13340 15866
rect 13392 15814 13410 15866
rect 13462 15814 13480 15866
rect 11720 15807 13490 15814
rect 2438 15802 13490 15807
rect 13596 15802 13602 15814
rect 2438 15781 13200 15802
rect 2274 15778 13200 15781
rect 2274 15768 4481 15778
rect 2274 15740 2550 15768
rect 2274 15706 2280 15740
rect 2314 15706 2404 15740
rect 2438 15734 2550 15740
rect 2584 15734 3406 15768
rect 3440 15734 4481 15768
rect 2438 15726 4481 15734
rect 4533 15726 4545 15778
rect 4597 15726 4609 15778
rect 4661 15768 13200 15778
rect 4661 15734 5062 15768
rect 5096 15734 6718 15768
rect 6752 15734 8374 15768
rect 8408 15734 10030 15768
rect 10064 15734 11686 15768
rect 11720 15750 13200 15768
rect 13252 15750 13270 15802
rect 13322 15750 13340 15802
rect 13392 15750 13410 15802
rect 13462 15750 13480 15802
rect 11720 15738 13490 15750
rect 13596 15738 13602 15750
rect 11720 15734 13200 15738
rect 4661 15726 13200 15734
rect 2438 15706 13200 15726
rect 2274 15695 13200 15706
rect 2274 15665 2550 15695
rect 2274 15631 2280 15665
rect 2314 15631 2404 15665
rect 2438 15661 2550 15665
rect 2584 15661 3406 15695
rect 3440 15661 5062 15695
rect 5096 15661 6718 15695
rect 6752 15661 8374 15695
rect 8408 15661 10030 15695
rect 10064 15661 11686 15695
rect 11720 15686 13200 15695
rect 13252 15686 13270 15738
rect 13322 15686 13340 15738
rect 13392 15686 13410 15738
rect 13462 15686 13480 15738
rect 11720 15674 13490 15686
rect 13596 15674 13602 15686
rect 11720 15661 13200 15674
rect 2438 15634 13200 15661
rect 2438 15631 4481 15634
rect 2274 15623 4481 15631
rect 2274 15589 2550 15623
rect 2584 15589 3406 15623
rect 3440 15589 4481 15623
rect 2274 15555 2280 15589
rect 2314 15555 2404 15589
rect 2438 15582 4481 15589
rect 4533 15582 4545 15634
rect 4597 15582 4609 15634
rect 4661 15623 13200 15634
rect 4661 15589 5062 15623
rect 5096 15589 6718 15623
rect 6752 15589 8374 15623
rect 8408 15589 10030 15623
rect 10064 15589 11686 15623
rect 11720 15622 13200 15623
rect 13252 15622 13270 15674
rect 13322 15622 13340 15674
rect 13392 15622 13410 15674
rect 13462 15622 13480 15674
rect 11720 15613 13342 15622
rect 13376 15613 13490 15622
rect 11720 15610 13490 15613
rect 13596 15610 13602 15622
rect 11720 15589 13200 15610
rect 4661 15582 13200 15589
rect 2438 15558 13200 15582
rect 13252 15558 13270 15610
rect 13322 15558 13340 15610
rect 13392 15558 13410 15610
rect 13462 15558 13480 15610
rect 2438 15555 13342 15558
rect 2274 15551 13342 15555
rect 2274 15517 2550 15551
rect 2584 15517 3406 15551
rect 3440 15517 5062 15551
rect 5096 15517 6718 15551
rect 6752 15517 8374 15551
rect 8408 15517 10030 15551
rect 10064 15517 11686 15551
rect 11720 15546 13342 15551
rect 13376 15546 13490 15558
rect 13596 15546 13602 15558
rect 11720 15517 13200 15546
rect 2274 15513 13200 15517
rect 2274 15479 2280 15513
rect 2314 15479 2404 15513
rect 2438 15494 13200 15513
rect 13252 15494 13270 15546
rect 13322 15494 13340 15546
rect 13392 15494 13410 15546
rect 13462 15494 13480 15546
rect 2438 15490 13342 15494
rect 2438 15479 4481 15490
rect 2274 15445 2550 15479
rect 2584 15445 3406 15479
rect 3440 15445 4481 15479
rect 2274 15438 4481 15445
rect 4533 15438 4545 15490
rect 4597 15438 4609 15490
rect 4661 15482 13342 15490
rect 13376 15482 13490 15494
rect 13596 15482 13602 15494
rect 4661 15479 13200 15482
rect 4661 15445 5062 15479
rect 5096 15445 6718 15479
rect 6752 15445 8374 15479
rect 8408 15445 10030 15479
rect 10064 15445 11686 15479
rect 11720 15445 13200 15479
rect 4661 15438 13200 15445
rect 2274 15437 13200 15438
rect 2274 15403 2280 15437
rect 2314 15403 2404 15437
rect 2438 15430 13200 15437
rect 13252 15430 13270 15482
rect 13322 15430 13340 15482
rect 13392 15430 13410 15482
rect 13462 15430 13480 15482
rect 2438 15419 13490 15430
rect 2438 15418 13342 15419
rect 13376 15418 13490 15419
rect 13596 15418 13602 15430
rect 2438 15407 13200 15418
rect 2438 15403 2550 15407
rect 2274 15373 2550 15403
rect 2584 15373 3406 15407
rect 3440 15373 5062 15407
rect 5096 15373 6718 15407
rect 6752 15373 8374 15407
rect 8408 15373 10030 15407
rect 10064 15373 11686 15407
rect 11720 15373 13200 15407
rect 2274 15366 13200 15373
rect 13252 15366 13270 15418
rect 13322 15366 13340 15418
rect 13392 15366 13410 15418
rect 13462 15366 13480 15418
rect 2274 15361 13490 15366
rect 2274 15327 2280 15361
rect 2314 15327 2404 15361
rect 2438 15354 13490 15361
rect 13596 15354 13602 15366
rect 2438 15346 13200 15354
rect 2438 15335 4481 15346
rect 2438 15327 2550 15335
rect 2274 15301 2550 15327
rect 2584 15301 3406 15335
rect 3440 15301 4481 15335
rect 2274 15294 4481 15301
rect 4533 15294 4545 15346
rect 4597 15294 4609 15346
rect 4661 15335 13200 15346
rect 4661 15301 5062 15335
rect 5096 15301 6718 15335
rect 6752 15301 8374 15335
rect 8408 15301 10030 15335
rect 10064 15301 11686 15335
rect 11720 15302 13200 15335
rect 13252 15302 13270 15354
rect 13322 15302 13340 15354
rect 13392 15302 13410 15354
rect 13462 15302 13480 15354
rect 11720 15301 13490 15302
rect 4661 15294 13490 15301
rect 2274 15290 13490 15294
rect 13596 15290 13602 15302
rect 2274 15285 13200 15290
rect 2274 15251 2280 15285
rect 2314 15251 2404 15285
rect 2438 15263 13200 15285
rect 2438 15251 2550 15263
rect 2274 15229 2550 15251
rect 2584 15229 3406 15263
rect 3440 15229 5062 15263
rect 5096 15229 6718 15263
rect 6752 15229 8374 15263
rect 8408 15229 10030 15263
rect 10064 15229 11686 15263
rect 11720 15238 13200 15263
rect 13252 15238 13270 15290
rect 13322 15238 13340 15290
rect 13392 15238 13410 15290
rect 13462 15238 13480 15290
rect 11720 15233 13342 15238
rect 13376 15233 13490 15238
rect 11720 15229 13490 15233
rect 2274 15226 13490 15229
rect 13596 15226 13602 15238
rect 2274 15209 13200 15226
rect 2274 15175 2280 15209
rect 2314 15175 2404 15209
rect 2438 15202 13200 15209
rect 2438 15191 4481 15202
rect 2438 15175 2550 15191
rect 2274 15157 2550 15175
rect 2584 15157 3406 15191
rect 3440 15157 4481 15191
rect 2274 15150 4481 15157
rect 4533 15150 4545 15202
rect 4597 15150 4609 15202
rect 4661 15191 13200 15202
rect 4661 15157 5062 15191
rect 5096 15157 6718 15191
rect 6752 15157 8374 15191
rect 8408 15157 10030 15191
rect 10064 15157 11686 15191
rect 11720 15174 13200 15191
rect 13252 15174 13270 15226
rect 13322 15174 13340 15226
rect 13392 15174 13410 15226
rect 13462 15174 13480 15226
rect 11720 15162 13342 15174
rect 13376 15162 13490 15174
rect 13596 15162 13602 15174
rect 11720 15157 13200 15162
rect 4661 15150 13200 15157
rect 2274 15143 13200 15150
tri 13012 15048 13107 15143 ne
rect 13107 15110 13200 15143
rect 13252 15110 13270 15162
rect 13322 15110 13340 15162
rect 13392 15110 13410 15162
rect 13462 15110 13480 15162
rect 13107 15098 13490 15110
rect 13596 15098 13602 15110
rect 13107 15048 13200 15098
rect 2504 15042 4849 15048
rect 1938 14974 2056 15006
rect 1938 14940 1944 14974
rect 1978 14940 2016 14974
rect 2050 14940 2056 14974
rect 1938 14899 2056 14940
rect 1938 14865 1944 14899
rect 1978 14865 2016 14899
rect 2050 14865 2056 14899
rect 1938 14824 2056 14865
rect 1938 14790 1944 14824
rect 1978 14790 2016 14824
rect 2050 14790 2056 14824
rect 1938 14749 2056 14790
rect 1938 14715 1944 14749
rect 1978 14715 2016 14749
rect 2050 14715 2056 14749
rect 1938 14674 2056 14715
rect 1938 14640 1944 14674
rect 1978 14640 2016 14674
rect 2050 14640 2056 14674
rect 1938 14599 2056 14640
rect 1938 14565 1944 14599
rect 1978 14565 2016 14599
rect 2050 14565 2056 14599
rect 1938 14524 2056 14565
rect 1938 14490 1944 14524
rect 1978 14490 2016 14524
rect 2050 14490 2056 14524
rect 1938 14449 2056 14490
rect 1938 14415 1944 14449
rect 1978 14415 2016 14449
rect 2050 14415 2056 14449
rect 1938 14374 2056 14415
rect 1938 14340 1944 14374
rect 1978 14340 2016 14374
rect 2050 14340 2056 14374
rect 1938 14299 2056 14340
rect 1938 14265 1944 14299
rect 1978 14265 2016 14299
rect 2050 14265 2056 14299
rect 1938 14224 2056 14265
rect 1938 14190 1944 14224
rect 1978 14190 2016 14224
rect 2050 14190 2056 14224
rect 1938 14149 2056 14190
rect 1938 14115 1944 14149
rect 1978 14115 2016 14149
rect 2050 14115 2056 14149
rect 1938 14075 2056 14115
rect 1938 14041 1944 14075
rect 1978 14041 2016 14075
rect 2050 14041 2056 14075
rect 1938 14001 2056 14041
rect 1938 13967 1944 14001
rect 1978 13967 2016 14001
rect 2050 13967 2056 14001
rect 1938 13927 2056 13967
rect 1938 13893 1944 13927
rect 1978 13893 2016 13927
rect 2050 13893 2056 13927
rect 1938 13853 2056 13893
rect 1938 13819 1944 13853
rect 1978 13819 2016 13853
rect 2050 13819 2056 13853
rect 1938 13779 2056 13819
rect 1938 13745 1944 13779
rect 1978 13745 2016 13779
rect 2050 13745 2056 13779
rect 1938 13705 2056 13745
rect 1938 13671 1944 13705
rect 1978 13671 2016 13705
rect 2050 13671 2056 13705
rect 1938 13631 2056 13671
rect 1938 13597 1944 13631
rect 1978 13597 2016 13631
rect 2050 13597 2056 13631
rect 1938 13557 2056 13597
rect 1938 13523 1944 13557
rect 1978 13523 2016 13557
rect 2050 13523 2056 13557
rect 1938 13483 2056 13523
rect 1938 13449 1944 13483
rect 1978 13449 2016 13483
rect 2050 13449 2056 13483
rect 1938 13409 2056 13449
rect 1938 13375 1944 13409
rect 1978 13375 2016 13409
rect 2050 13375 2056 13409
rect 1938 13335 2056 13375
rect 1938 13301 1944 13335
rect 1978 13301 2016 13335
rect 2050 13301 2056 13335
rect 1938 13269 2056 13301
rect 2274 14987 2444 15019
rect 2274 14953 2280 14987
rect 2314 14953 2404 14987
rect 2438 14953 2444 14987
rect 2274 14912 2444 14953
rect 2274 14878 2280 14912
rect 2314 14878 2404 14912
rect 2438 14878 2444 14912
rect 2274 14837 2444 14878
rect 2274 14803 2280 14837
rect 2314 14803 2404 14837
rect 2438 14803 2444 14837
rect 2274 14762 2444 14803
rect 2274 14728 2280 14762
rect 2314 14728 2404 14762
rect 2438 14728 2444 14762
rect 2274 14687 2444 14728
rect 2274 14653 2280 14687
rect 2314 14653 2404 14687
rect 2438 14653 2444 14687
rect 2274 14612 2444 14653
rect 2274 14578 2280 14612
rect 2314 14578 2404 14612
rect 2438 14578 2444 14612
rect 2274 14537 2444 14578
rect 2274 14503 2280 14537
rect 2314 14503 2404 14537
rect 2438 14503 2444 14537
rect 2274 14462 2444 14503
rect 2274 14428 2280 14462
rect 2314 14428 2404 14462
rect 2438 14428 2444 14462
rect 2274 14387 2444 14428
rect 2274 14353 2280 14387
rect 2314 14353 2404 14387
rect 2438 14353 2444 14387
rect 2274 14312 2444 14353
rect 2274 14278 2280 14312
rect 2314 14278 2404 14312
rect 2438 14278 2444 14312
rect 2274 14237 2444 14278
rect 2274 14203 2280 14237
rect 2314 14203 2404 14237
rect 2438 14203 2444 14237
rect 2274 14162 2444 14203
rect 2274 14128 2280 14162
rect 2314 14128 2404 14162
rect 2438 14128 2444 14162
rect 2274 14087 2444 14128
rect 2274 14053 2280 14087
rect 2314 14053 2404 14087
rect 2438 14053 2444 14087
rect 2274 14012 2444 14053
rect 2274 13978 2280 14012
rect 2314 13978 2404 14012
rect 2438 13978 2444 14012
rect 2274 13937 2444 13978
rect 2274 13903 2280 13937
rect 2314 13903 2404 13937
rect 2438 13903 2444 13937
rect 2274 13862 2444 13903
rect 2274 13828 2280 13862
rect 2314 13828 2404 13862
rect 2438 13828 2444 13862
rect 2274 13787 2444 13828
rect 2274 13753 2280 13787
rect 2314 13753 2404 13787
rect 2438 13753 2444 13787
rect 2274 13712 2444 13753
rect 2274 13678 2280 13712
rect 2314 13678 2404 13712
rect 2438 13678 2444 13712
rect 2274 13636 2444 13678
rect 2274 13602 2280 13636
rect 2314 13602 2404 13636
rect 2438 13602 2444 13636
rect 2274 13560 2444 13602
rect 2274 13526 2280 13560
rect 2314 13526 2404 13560
rect 2438 13526 2444 13560
rect 2274 13484 2444 13526
rect 2274 13450 2280 13484
rect 2314 13450 2404 13484
rect 2438 13450 2444 13484
rect 2274 13408 2444 13450
rect 2274 13374 2280 13408
rect 2314 13374 2404 13408
rect 2438 13374 2444 13408
rect 2274 13332 2444 13374
rect 2274 13298 2280 13332
rect 2314 13298 2404 13332
rect 2438 13298 2444 13332
rect 2274 13266 2444 13298
rect 2504 14990 4731 15042
rect 4783 14990 4797 15042
rect 2504 14921 4849 14990
tri 13107 14956 13199 15048 ne
rect 13199 15046 13200 15048
rect 13252 15046 13270 15098
rect 13322 15046 13340 15098
rect 13392 15046 13410 15098
rect 13462 15046 13480 15098
rect 13199 15034 13490 15046
rect 13596 15034 13602 15046
rect 13199 14982 13200 15034
rect 13252 14982 13270 15034
rect 13322 14982 13340 15034
rect 13392 14982 13410 15034
rect 13462 14982 13480 15034
rect 13199 14970 13490 14982
rect 13596 14970 13602 14982
rect 2504 14869 4731 14921
rect 4783 14869 4797 14921
rect 2504 14863 4849 14869
rect 13199 14918 13200 14970
rect 13252 14918 13270 14970
rect 13322 14918 13340 14970
rect 13392 14918 13410 14970
rect 13462 14918 13480 14970
rect 13199 14906 13490 14918
rect 13596 14906 13602 14918
tri 2474 13230 2504 13260 se
rect 2504 13230 2627 14863
tri 2627 14838 2652 14863 nw
rect 13199 14854 13200 14906
rect 13252 14854 13270 14906
rect 13322 14854 13340 14906
rect 13392 14854 13410 14906
rect 13462 14854 13480 14906
rect 13199 14842 13490 14854
rect 13596 14842 13602 14854
rect 13199 14790 13200 14842
rect 13252 14790 13270 14842
rect 13322 14790 13340 14842
rect 13392 14790 13410 14842
rect 13462 14790 13480 14842
rect 13199 14778 13490 14790
rect 13596 14778 13602 14790
rect 13199 14726 13200 14778
rect 13252 14726 13270 14778
rect 13322 14726 13340 14778
rect 13392 14726 13410 14778
rect 13462 14726 13480 14778
rect 3227 14720 3345 14726
rect 3279 14668 3293 14720
rect 3227 14654 3345 14668
rect 3279 14602 3293 14654
rect 3227 14588 3345 14602
rect 3279 14536 3293 14588
rect 3227 14522 3345 14536
rect 3279 14470 3293 14522
rect 3227 14456 3345 14470
rect 3279 14404 3293 14456
rect 3227 14390 3345 14404
rect 2673 14345 2859 14357
rect 2673 14311 2679 14345
rect 2713 14311 2751 14345
rect 2785 14311 2859 14345
rect 2673 14267 2859 14311
rect 2673 14233 2679 14267
rect 2713 14233 2751 14267
rect 2785 14233 2859 14267
rect 2673 14189 2859 14233
rect 2673 14155 2679 14189
rect 2713 14155 2751 14189
rect 2785 14155 2859 14189
rect 2673 14111 2859 14155
rect 2673 14077 2679 14111
rect 2713 14077 2751 14111
rect 2785 14077 2859 14111
rect 2673 14033 2859 14077
rect 2673 13999 2679 14033
rect 2713 13999 2751 14033
rect 2785 13999 2859 14033
rect 2673 13955 2859 13999
rect 2673 13921 2679 13955
rect 2713 13921 2751 13955
rect 2785 13921 2859 13955
rect 2673 13877 2859 13921
rect 2673 13843 2679 13877
rect 2713 13843 2751 13877
rect 2785 13843 2859 13877
rect 2673 13799 2859 13843
rect 2673 13765 2679 13799
rect 2713 13765 2751 13799
rect 2785 13765 2859 13799
rect 2673 13722 2859 13765
rect 2673 13688 2679 13722
rect 2713 13688 2751 13722
rect 2785 13688 2859 13722
rect 2673 13645 2859 13688
rect 2673 13611 2679 13645
rect 2713 13611 2751 13645
rect 2785 13611 2859 13645
rect 2673 13568 2859 13611
rect 2673 13534 2679 13568
rect 2713 13534 2751 13568
rect 2785 13534 2859 13568
rect 2673 13491 2859 13534
rect 2673 13457 2679 13491
rect 2713 13457 2751 13491
rect 2785 13457 2859 13491
rect 2673 13414 2859 13457
rect 2673 13380 2679 13414
rect 2713 13380 2751 13414
rect 2785 13380 2859 13414
rect 2950 14345 3068 14357
rect 2950 14311 2956 14345
rect 2990 14311 3028 14345
rect 3062 14311 3068 14345
rect 2950 14267 3068 14311
rect 2950 14233 2956 14267
rect 2990 14233 3028 14267
rect 3062 14233 3068 14267
rect 2950 14189 3068 14233
rect 2950 14155 2956 14189
rect 2990 14155 3028 14189
rect 3062 14155 3068 14189
rect 2950 14111 3068 14155
rect 2950 14077 2956 14111
rect 2990 14077 3028 14111
rect 3062 14077 3068 14111
rect 2950 14033 3068 14077
rect 2950 13999 2956 14033
rect 2990 13999 3028 14033
rect 3062 13999 3068 14033
rect 2950 13955 3068 13999
rect 2950 13921 2956 13955
rect 2990 13921 3028 13955
rect 3062 13921 3068 13955
rect 2950 13892 3068 13921
rect 3002 13840 3016 13892
rect 2950 13826 3068 13840
rect 3002 13774 3016 13826
rect 2950 13765 2956 13774
rect 2990 13765 3028 13774
rect 3062 13765 3068 13774
rect 2950 13760 3068 13765
rect 3002 13708 3016 13760
rect 2950 13694 2956 13708
rect 2990 13694 3028 13708
rect 3062 13694 3068 13708
rect 3002 13642 3016 13694
rect 2950 13628 2956 13642
rect 2990 13628 3028 13642
rect 3062 13628 3068 13642
rect 3002 13576 3016 13628
rect 2950 13568 3068 13576
rect 2950 13562 2956 13568
rect 2990 13562 3028 13568
rect 3062 13562 3068 13568
rect 3002 13510 3016 13562
rect 2950 13495 3068 13510
rect 3002 13443 3016 13495
rect 2950 13428 3068 13443
tri 2859 13380 2889 13410 sw
rect 2673 13370 2889 13380
tri 2889 13370 2899 13380 sw
rect 3002 13376 3016 13428
rect 2673 13368 2899 13370
tri 2759 13351 2776 13368 ne
rect 2776 13351 2899 13368
tri 2899 13351 2918 13370 sw
tri 2776 13309 2818 13351 ne
tri 2627 13230 2657 13260 sw
rect 1487 13218 2781 13230
rect 1487 13184 2669 13218
rect 2703 13184 2741 13218
rect 2775 13184 2781 13218
rect 1487 13111 2781 13184
rect 1487 13077 2669 13111
rect 2703 13077 2741 13111
rect 2775 13077 2781 13111
rect 1487 13004 2781 13077
rect 1487 12970 2669 13004
rect 2703 12970 2741 13004
rect 2775 12970 2781 13004
rect 1487 12958 2781 12970
rect 1487 12889 1828 12958
tri 1828 12889 1897 12958 nw
tri 2793 12921 2818 12946 se
rect 2818 12921 2918 13351
rect 1938 12889 2056 12921
tri 2776 12904 2793 12921 se
rect 2793 12904 2918 12921
rect 1487 12855 1794 12889
tri 1794 12855 1828 12889 nw
rect 1938 12855 1944 12889
rect 1978 12855 2016 12889
rect 2050 12855 2056 12889
rect 1487 12814 1753 12855
tri 1753 12814 1794 12855 nw
rect 1938 12814 2056 12855
rect 1487 12801 1740 12814
tri 1740 12801 1753 12814 nw
rect 1487 12780 1719 12801
tri 1719 12780 1740 12801 nw
rect 1938 12780 1944 12814
rect 1978 12780 2016 12814
rect 2050 12780 2056 12814
tri 2673 12801 2776 12904 se
rect 2776 12801 2815 12904
tri 2815 12801 2918 12904 nw
rect 1487 11414 1687 12780
tri 1687 12748 1719 12780 nw
rect 1938 12739 2056 12780
rect 1938 12705 1944 12739
rect 1978 12705 2016 12739
rect 2050 12705 2056 12739
rect 1938 12664 2056 12705
rect 1938 12630 1944 12664
rect 1978 12630 2016 12664
rect 2050 12630 2056 12664
rect 1938 12589 2056 12630
rect 1938 12555 1944 12589
rect 1978 12555 2016 12589
rect 2050 12555 2056 12589
rect 1938 12514 2056 12555
rect 1938 12480 1944 12514
rect 1978 12480 2016 12514
rect 2050 12480 2056 12514
rect 1938 12439 2056 12480
rect 1938 12405 1944 12439
rect 1978 12405 2016 12439
rect 2050 12405 2056 12439
rect 1938 12364 2056 12405
rect 1938 12330 1944 12364
rect 1978 12330 2016 12364
rect 2050 12330 2056 12364
rect 1938 12289 2056 12330
rect 1938 12255 1944 12289
rect 1978 12255 2016 12289
rect 2050 12255 2056 12289
rect 1938 12214 2056 12255
rect 1938 12180 1944 12214
rect 1978 12180 2016 12214
rect 2050 12180 2056 12214
rect 1938 12139 2056 12180
rect 1938 12105 1944 12139
rect 1978 12105 2016 12139
rect 2050 12105 2056 12139
rect 1938 12064 2056 12105
rect 1938 12030 1944 12064
rect 1978 12030 2016 12064
rect 2050 12030 2056 12064
rect 1938 11989 2056 12030
rect 1938 11955 1944 11989
rect 1978 11955 2016 11989
rect 2050 11955 2056 11989
rect 1938 11914 2056 11955
rect 1938 11880 1944 11914
rect 1978 11880 2016 11914
rect 2050 11880 2056 11914
rect 1938 11839 2056 11880
rect 1938 11805 1944 11839
rect 1978 11805 2016 11839
rect 2050 11805 2056 11839
rect 1938 11764 2056 11805
rect 1938 11730 1944 11764
rect 1978 11730 2016 11764
rect 2050 11730 2056 11764
rect 1938 11689 2056 11730
rect 1938 11655 1944 11689
rect 1978 11655 2016 11689
rect 2050 11655 2056 11689
rect 1938 11614 2056 11655
rect 1938 11580 1944 11614
rect 1978 11580 2016 11614
rect 2050 11580 2056 11614
rect 1938 11539 2056 11580
rect 1938 11505 1944 11539
rect 1978 11505 2016 11539
rect 2050 11505 2056 11539
rect 1938 11464 2056 11505
rect 1938 11430 1944 11464
rect 1978 11430 2016 11464
rect 2050 11430 2056 11464
tri 1687 11414 1689 11416 sw
rect 1487 11389 1689 11414
tri 1689 11389 1714 11414 sw
rect 1938 11389 2056 11430
rect 1487 11368 1714 11389
tri 1714 11368 1735 11389 sw
rect 1487 11355 1735 11368
tri 1735 11355 1748 11368 sw
rect 1938 11355 1944 11389
rect 1978 11355 2016 11389
rect 2050 11355 2056 11389
rect 2249 12789 2791 12801
rect 2249 11891 2255 12789
rect 2361 12714 2791 12789
tri 2791 12777 2815 12801 nw
rect 2361 12680 2679 12714
rect 2713 12680 2751 12714
rect 2785 12680 2791 12714
rect 2361 12641 2791 12680
rect 2361 12607 2679 12641
rect 2713 12607 2751 12641
rect 2785 12607 2791 12641
rect 2361 12568 2791 12607
rect 2361 12534 2679 12568
rect 2713 12534 2751 12568
rect 2785 12534 2791 12568
rect 2361 12495 2791 12534
rect 2361 12461 2679 12495
rect 2713 12461 2751 12495
rect 2785 12461 2791 12495
rect 2361 12422 2791 12461
rect 2361 11891 2679 12422
rect 2249 11852 2679 11891
rect 2249 11818 2255 11852
rect 2289 11818 2327 11852
rect 2361 11818 2679 11852
rect 2249 11779 2679 11818
rect 2249 11745 2255 11779
rect 2289 11745 2327 11779
rect 2361 11745 2679 11779
rect 2249 11706 2679 11745
rect 2249 11672 2255 11706
rect 2289 11672 2327 11706
rect 2361 11672 2679 11706
rect 2249 11633 2679 11672
rect 2249 11599 2255 11633
rect 2289 11599 2327 11633
rect 2361 11599 2679 11633
rect 2249 11560 2679 11599
rect 2249 11526 2255 11560
rect 2289 11526 2327 11560
rect 2361 11526 2679 11560
rect 2249 11487 2679 11526
rect 2249 11453 2255 11487
rect 2289 11453 2327 11487
rect 2361 11453 2679 11487
rect 2249 11414 2679 11453
rect 2249 11380 2255 11414
rect 2289 11380 2327 11414
rect 2361 11380 2679 11414
rect 2785 11380 2791 12422
rect 2249 11370 2791 11380
rect 2950 12714 3068 13376
rect 2950 12680 2956 12714
rect 2990 12680 3028 12714
rect 3062 12680 3068 12714
rect 2950 12641 3068 12680
rect 2950 12607 2956 12641
rect 2990 12607 3028 12641
rect 3062 12607 3068 12641
rect 2950 12568 3068 12607
rect 2950 12534 2956 12568
rect 2990 12534 3028 12568
rect 3062 12534 3068 12568
rect 2950 12495 3068 12534
rect 2950 12461 2956 12495
rect 2990 12461 3028 12495
rect 3062 12461 3068 12495
rect 2950 12422 3068 12461
rect 2950 11892 2956 12422
rect 3062 11892 3068 12422
rect 2950 11826 2956 11840
rect 3062 11826 3068 11840
rect 2950 11760 2956 11774
rect 3062 11760 3068 11774
rect 2950 11694 2956 11708
rect 3062 11694 3068 11708
rect 2950 11628 2956 11642
rect 3062 11628 3068 11642
rect 2950 11562 2956 11576
rect 3062 11562 3068 11576
rect 2950 11495 2956 11510
rect 3062 11495 3068 11510
rect 2950 11428 2956 11443
rect 3062 11428 3068 11443
rect 3002 11376 3016 11380
tri 2791 11370 2796 11375 sw
rect 2249 11368 2796 11370
tri 2796 11368 2798 11370 sw
rect 1487 11313 1748 11355
tri 1748 11313 1790 11355 sw
rect 1938 11313 2056 11355
tri 2657 11334 2691 11368 ne
rect 1487 11279 1790 11313
tri 1790 11279 1824 11313 sw
rect 1938 11279 1944 11313
rect 1978 11279 2016 11313
rect 2050 11279 2056 11313
rect 1487 11206 1824 11279
tri 1824 11206 1897 11279 sw
rect 1938 11247 2056 11279
rect 2691 11333 2798 11368
tri 2691 11248 2776 11333 ne
rect 2776 11248 2798 11333
tri 2798 11248 2918 11368 sw
tri 2776 11247 2777 11248 ne
rect 2777 11247 2918 11248
tri 2777 11233 2791 11247 ne
rect 2791 11233 2918 11247
tri 2791 11206 2818 11233 ne
rect 1487 11194 2750 11206
rect 1487 11160 2638 11194
rect 2672 11160 2710 11194
rect 2744 11160 2750 11194
rect 1487 11087 2750 11160
rect 1487 11053 2638 11087
rect 2672 11053 2710 11087
rect 2744 11053 2750 11087
rect 1487 10980 2750 11053
rect 1487 10946 2638 10980
rect 2672 10946 2710 10980
rect 2744 10946 2750 10980
rect 1487 10934 2750 10946
rect 1487 10847 1810 10934
tri 1810 10847 1897 10934 nw
tri 2802 10879 2818 10895 se
rect 2818 10879 2918 11233
rect 1938 10847 2056 10879
tri 2776 10853 2802 10879 se
rect 2802 10853 2918 10879
rect 1487 10813 1776 10847
tri 1776 10813 1810 10847 nw
rect 1938 10813 1944 10847
rect 1978 10813 2016 10847
rect 2050 10813 2056 10847
rect 1487 10771 1734 10813
tri 1734 10771 1776 10813 nw
rect 1938 10771 2056 10813
rect 1487 10737 1700 10771
tri 1700 10737 1734 10771 nw
rect 1938 10737 1944 10771
rect 1978 10737 2016 10771
rect 2050 10737 2056 10771
rect 1487 9420 1687 10737
tri 1687 10724 1700 10737 nw
rect 1938 10695 2056 10737
tri 2649 10726 2776 10853 se
rect 2776 10730 2795 10853
tri 2795 10730 2918 10853 nw
rect 2776 10726 2791 10730
tri 2791 10726 2795 10730 nw
rect 1938 10661 1944 10695
rect 1978 10661 2016 10695
rect 2050 10661 2056 10695
rect 1938 10620 2056 10661
rect 1938 10586 1944 10620
rect 1978 10586 2016 10620
rect 2050 10586 2056 10620
rect 1938 10545 2056 10586
rect 1938 10511 1944 10545
rect 1978 10511 2016 10545
rect 2050 10511 2056 10545
rect 1938 10470 2056 10511
rect 1938 10436 1944 10470
rect 1978 10436 2016 10470
rect 2050 10436 2056 10470
rect 1938 10395 2056 10436
rect 1938 10361 1944 10395
rect 1978 10361 2016 10395
rect 2050 10361 2056 10395
rect 1938 10320 2056 10361
rect 1938 10286 1944 10320
rect 1978 10286 2016 10320
rect 2050 10286 2056 10320
rect 1938 10245 2056 10286
rect 1938 10211 1944 10245
rect 1978 10211 2016 10245
rect 2050 10211 2056 10245
rect 1938 10170 2056 10211
rect 1938 10136 1944 10170
rect 1978 10136 2016 10170
rect 2050 10136 2056 10170
rect 1938 10095 2056 10136
rect 1938 10061 1944 10095
rect 1978 10061 2016 10095
rect 2050 10061 2056 10095
rect 1938 10020 2056 10061
rect 1938 9986 1944 10020
rect 1978 9986 2016 10020
rect 2050 9986 2056 10020
rect 1938 9945 2056 9986
rect 1938 9911 1944 9945
rect 1978 9911 2016 9945
rect 2050 9911 2056 9945
rect 1938 9870 2056 9911
rect 1938 9836 1944 9870
rect 1978 9836 2016 9870
rect 2050 9836 2056 9870
rect 1938 9795 2056 9836
rect 1938 9761 1944 9795
rect 1978 9761 2016 9795
rect 2050 9761 2056 9795
rect 1938 9720 2056 9761
rect 1938 9686 1944 9720
rect 1978 9686 2016 9720
rect 2050 9686 2056 9720
rect 1938 9645 2056 9686
rect 1938 9611 1944 9645
rect 1978 9611 2016 9645
rect 2050 9611 2056 9645
rect 1938 9570 2056 9611
rect 1938 9536 1944 9570
rect 1978 9536 2016 9570
rect 2050 9536 2056 9570
rect 1938 9495 2056 9536
rect 1938 9461 1944 9495
rect 1978 9461 2016 9495
rect 2050 9461 2056 9495
tri 1687 9420 1707 9440 sw
rect 1938 9420 2056 9461
rect 1487 9416 1707 9420
tri 1707 9416 1711 9420 sw
rect 1487 9386 1711 9416
tri 1711 9386 1741 9416 sw
rect 1938 9386 1944 9420
rect 1978 9386 2016 9420
rect 2050 9386 2056 9420
rect 1487 9381 1741 9386
tri 1741 9381 1746 9386 sw
rect 1487 9380 1746 9381
tri 1746 9380 1747 9381 sw
rect 1487 9245 1747 9380
tri 1747 9245 1882 9380 sw
rect 1938 9354 2056 9386
rect 2249 10714 2791 10726
rect 2249 9600 2255 10714
rect 2361 10680 2679 10714
rect 2713 10680 2751 10714
rect 2785 10680 2791 10714
rect 2361 10641 2791 10680
rect 2361 10607 2679 10641
rect 2713 10607 2751 10641
rect 2785 10607 2791 10641
rect 2361 10568 2791 10607
rect 2361 10534 2679 10568
rect 2713 10534 2751 10568
rect 2785 10534 2791 10568
rect 2361 10495 2791 10534
rect 2361 10461 2679 10495
rect 2713 10461 2751 10495
rect 2785 10461 2791 10495
rect 2361 10422 2791 10461
rect 2361 9600 2679 10422
rect 2249 9561 2679 9600
rect 2249 9527 2255 9561
rect 2289 9527 2327 9561
rect 2361 9527 2679 9561
rect 2249 9488 2679 9527
rect 2249 9454 2255 9488
rect 2289 9454 2327 9488
rect 2361 9454 2679 9488
rect 2249 9415 2679 9454
rect 2249 9381 2255 9415
rect 2289 9381 2327 9415
rect 2361 9381 2679 9415
rect 2249 9380 2679 9381
rect 2785 9380 2791 10422
rect 2249 9366 2791 9380
rect 2950 10714 3068 11376
rect 2950 10680 2956 10714
rect 2990 10680 3028 10714
rect 3062 10680 3068 10714
rect 2950 10641 3068 10680
rect 2950 10607 2956 10641
rect 2990 10607 3028 10641
rect 3062 10607 3068 10641
rect 2950 10568 3068 10607
rect 2950 10534 2956 10568
rect 2990 10534 3028 10568
rect 3062 10534 3068 10568
rect 2950 10495 3068 10534
rect 2950 10461 2956 10495
rect 2990 10461 3028 10495
rect 3062 10461 3068 10495
rect 2950 10422 3068 10461
rect 2950 9896 2956 10422
rect 3062 9896 3068 10422
rect 2950 9830 2956 9844
rect 3062 9830 3068 9844
rect 2950 9764 2956 9778
rect 3062 9764 3068 9778
rect 2950 9698 2956 9712
rect 3062 9698 3068 9712
rect 2950 9632 2956 9646
rect 3062 9632 3068 9646
rect 2950 9566 2956 9580
rect 3062 9566 3068 9580
rect 2950 9499 2956 9514
rect 3062 9499 3068 9514
rect 2950 9432 2956 9447
rect 3062 9432 3068 9447
tri 2656 9354 2668 9366 ne
rect 2668 9354 2791 9366
tri 2668 9331 2691 9354 ne
rect 2691 9330 2791 9354
tri 2691 9245 2776 9330 ne
rect 2776 9245 2791 9330
tri 2791 9245 2918 9372 sw
rect 1487 9233 2724 9245
rect 1487 9199 2612 9233
rect 2646 9199 2684 9233
rect 2718 9199 2724 9233
tri 2776 9230 2791 9245 ne
rect 2791 9230 2918 9245
tri 2791 9203 2818 9230 ne
rect 1487 9160 2724 9199
rect 1487 9126 2612 9160
rect 2646 9126 2684 9160
rect 2718 9126 2724 9160
rect 1487 9086 2724 9126
rect 1487 9052 2612 9086
rect 2646 9052 2684 9086
rect 2718 9052 2724 9086
rect 1487 9012 2724 9052
rect 1487 8978 2612 9012
rect 2646 8978 2684 9012
rect 2718 8978 2724 9012
rect 1487 8938 2724 8978
rect 1487 8904 2612 8938
rect 2646 8904 2684 8938
rect 2718 8904 2724 8938
rect 1487 8892 2724 8904
rect 1487 7433 1687 8892
tri 1687 8748 1831 8892 nw
tri 2776 8850 2818 8892 se
rect 2818 8850 2918 9230
tri 2690 8764 2776 8850 se
rect 2776 8764 2816 8850
rect 1938 8732 2056 8764
tri 2674 8748 2690 8764 se
rect 2690 8748 2816 8764
tri 2816 8748 2918 8850 nw
tri 2662 8736 2674 8748 se
rect 2674 8736 2794 8748
rect 1938 7618 1944 8732
rect 2050 7618 2056 8732
rect 1938 7579 2056 7618
rect 1938 7545 1944 7579
rect 1978 7545 2016 7579
rect 2050 7545 2056 7579
rect 1938 7513 2056 7545
rect 2249 8726 2794 8736
tri 2794 8726 2816 8748 nw
rect 2249 8724 2791 8726
rect 2249 8690 2255 8724
rect 2289 8690 2327 8724
rect 2361 8714 2791 8724
tri 2791 8723 2794 8726 nw
rect 2361 8690 2679 8714
rect 2249 8680 2679 8690
rect 2713 8680 2751 8714
rect 2785 8680 2791 8714
rect 2249 8651 2791 8680
rect 2249 8617 2255 8651
rect 2289 8617 2327 8651
rect 2361 8641 2791 8651
rect 2361 8617 2679 8641
rect 2249 8607 2679 8617
rect 2713 8607 2751 8641
rect 2785 8607 2791 8641
rect 2249 8577 2791 8607
rect 2249 8543 2255 8577
rect 2289 8543 2327 8577
rect 2361 8568 2791 8577
rect 2361 8543 2679 8568
rect 2249 8534 2679 8543
rect 2713 8534 2751 8568
rect 2785 8534 2791 8568
rect 2249 8503 2791 8534
rect 2249 8469 2255 8503
rect 2289 8469 2327 8503
rect 2361 8495 2791 8503
rect 2361 8469 2679 8495
rect 2249 8461 2679 8469
rect 2713 8461 2751 8495
rect 2785 8461 2791 8495
rect 2249 8429 2791 8461
rect 2249 8395 2255 8429
rect 2289 8395 2327 8429
rect 2361 8422 2791 8429
rect 2361 8395 2679 8422
rect 2249 8355 2679 8395
rect 2249 8321 2255 8355
rect 2289 8321 2327 8355
rect 2361 8321 2679 8355
rect 2249 8281 2679 8321
rect 2249 8247 2255 8281
rect 2289 8247 2327 8281
rect 2361 8247 2679 8281
rect 2249 8207 2679 8247
rect 2249 8173 2255 8207
rect 2289 8173 2327 8207
rect 2361 8173 2679 8207
rect 2249 8133 2679 8173
rect 2249 8099 2255 8133
rect 2289 8099 2327 8133
rect 2361 8099 2679 8133
rect 2249 8059 2679 8099
rect 2249 8025 2255 8059
rect 2289 8025 2327 8059
rect 2361 8025 2679 8059
rect 2249 7985 2679 8025
rect 2249 7951 2255 7985
rect 2289 7951 2327 7985
rect 2361 7951 2679 7985
rect 2249 7911 2679 7951
rect 2249 7877 2255 7911
rect 2289 7877 2327 7911
rect 2361 7877 2679 7911
rect 2249 7837 2679 7877
rect 2249 7803 2255 7837
rect 2289 7803 2327 7837
rect 2361 7803 2679 7837
rect 2249 7763 2679 7803
rect 2249 7729 2255 7763
rect 2289 7729 2327 7763
rect 2361 7729 2679 7763
rect 2249 7689 2679 7729
rect 2249 7655 2255 7689
rect 2289 7655 2327 7689
rect 2361 7655 2679 7689
rect 2249 7615 2679 7655
rect 2249 7581 2255 7615
rect 2289 7581 2327 7615
rect 2361 7581 2679 7615
rect 2249 7541 2679 7581
rect 2249 7507 2255 7541
rect 2289 7507 2327 7541
rect 2361 7507 2679 7541
rect 2249 7467 2679 7507
tri 1687 7433 1705 7451 sw
rect 2249 7433 2255 7467
rect 2289 7433 2327 7467
rect 2361 7433 2679 7467
rect 1487 7393 1705 7433
tri 1705 7393 1745 7433 sw
rect 2249 7393 2679 7433
rect 1487 7368 1745 7393
tri 1745 7368 1770 7393 sw
rect 1487 7359 1770 7368
tri 1770 7359 1779 7368 sw
rect 2249 7359 2255 7393
rect 2289 7359 2327 7393
rect 2361 7380 2679 7393
rect 2785 7380 2791 8422
rect 2950 8714 3068 9380
rect 2950 8680 2956 8714
rect 2990 8680 3028 8714
rect 3062 8680 3068 8714
rect 2950 8641 3068 8680
rect 2950 8607 2956 8641
rect 2990 8607 3028 8641
rect 3062 8607 3068 8641
rect 2950 8568 3068 8607
rect 2950 8534 2956 8568
rect 2990 8534 3028 8568
rect 3062 8534 3068 8568
rect 2950 8495 3068 8534
rect 2950 8461 2956 8495
rect 2990 8461 3028 8495
rect 3062 8461 3068 8495
rect 2950 8422 3068 8461
rect 2950 7892 2956 8422
rect 3062 7892 3068 8422
rect 2950 7826 2956 7840
rect 3062 7826 3068 7840
rect 2950 7760 2956 7774
rect 3062 7760 3068 7774
rect 2950 7694 2956 7708
rect 3062 7694 3068 7708
rect 2950 7628 2956 7642
rect 3062 7628 3068 7642
rect 2950 7562 2956 7576
rect 3062 7562 3068 7576
rect 2950 7495 2956 7510
rect 3062 7495 3068 7510
rect 2950 7428 2956 7443
rect 3062 7428 3068 7443
tri 2791 7380 2825 7414 sw
rect 2361 7368 2825 7380
tri 2825 7368 2837 7380 sw
rect 3002 7376 3016 7380
rect 2361 7359 2837 7368
rect 1487 7255 1779 7359
tri 1779 7255 1883 7359 sw
rect 2249 7347 2837 7359
tri 2716 7287 2776 7347 ne
rect 2776 7287 2837 7347
tri 2837 7287 2918 7368 sw
tri 2776 7272 2791 7287 ne
rect 2791 7272 2918 7287
tri 2791 7255 2808 7272 ne
rect 2808 7255 2918 7272
rect 1487 7243 2750 7255
tri 2808 7245 2818 7255 ne
rect 1487 7209 2638 7243
rect 2672 7209 2710 7243
rect 2744 7209 2750 7243
rect 1487 7153 2750 7209
rect 1487 7119 2638 7153
rect 2672 7119 2710 7153
rect 2744 7119 2750 7153
rect 1487 7063 2750 7119
rect 1487 7029 2638 7063
rect 2672 7029 2710 7063
rect 2744 7029 2750 7063
rect 1487 6972 2750 7029
rect 1487 6938 2638 6972
rect 2672 6938 2710 6972
rect 2744 6938 2750 6972
rect 1487 6926 2750 6938
tri 2810 6926 2818 6934 se
rect 2818 6926 2918 7255
rect 1487 6820 1748 6926
tri 1748 6820 1854 6926 nw
tri 2776 6892 2810 6926 se
rect 2810 6892 2918 6926
tri 2705 6821 2776 6892 se
rect 2776 6821 2846 6892
rect 2249 6820 2846 6821
tri 2846 6820 2918 6892 nw
rect 1487 6808 1736 6820
tri 1736 6808 1748 6820 nw
rect 2249 6808 2791 6820
rect 1487 6774 1702 6808
tri 1702 6774 1736 6808 nw
rect 2249 6774 2255 6808
rect 2289 6774 2327 6808
rect 2361 6774 2791 6808
rect 1487 4837 1687 6774
tri 1687 6759 1702 6774 nw
rect 2249 6735 2791 6774
tri 2791 6765 2846 6820 nw
rect 2249 6701 2255 6735
rect 2289 6701 2327 6735
rect 2361 6714 2791 6735
rect 2361 6701 2679 6714
rect 2249 6680 2679 6701
rect 2713 6680 2751 6714
rect 2785 6680 2791 6714
rect 2249 6662 2791 6680
rect 2249 6628 2255 6662
rect 2289 6628 2327 6662
rect 2361 6641 2791 6662
rect 2361 6628 2679 6641
rect 2249 6607 2679 6628
rect 2713 6607 2751 6641
rect 2785 6607 2791 6641
rect 1938 6560 2056 6592
rect 1938 6526 1944 6560
rect 1978 6526 2016 6560
rect 2050 6526 2056 6560
rect 1938 6487 2056 6526
rect 1938 6453 1944 6487
rect 1978 6453 2016 6487
rect 2050 6453 2056 6487
rect 1938 6414 2056 6453
rect 1938 6380 1944 6414
rect 1978 6380 2016 6414
rect 2050 6380 2056 6414
rect 1938 6341 2056 6380
rect 1938 6307 1944 6341
rect 1978 6307 2016 6341
rect 2050 6307 2056 6341
rect 1938 6268 2056 6307
rect 1938 6234 1944 6268
rect 1978 6234 2016 6268
rect 2050 6234 2056 6268
rect 1938 6195 2056 6234
rect 1938 6161 1944 6195
rect 1978 6161 2016 6195
rect 2050 6161 2056 6195
rect 1938 6122 2056 6161
rect 1938 6088 1944 6122
rect 1978 6088 2016 6122
rect 2050 6088 2056 6122
rect 1938 6049 2056 6088
rect 1938 6015 1944 6049
rect 1978 6015 2016 6049
rect 2050 6015 2056 6049
rect 1938 5976 2056 6015
rect 1938 5942 1944 5976
rect 1978 5942 2016 5976
rect 2050 5942 2056 5976
rect 1938 5903 2056 5942
rect 1938 5869 1944 5903
rect 1978 5869 2016 5903
rect 2050 5869 2056 5903
rect 1938 5830 2056 5869
rect 1938 5796 1944 5830
rect 1978 5796 2016 5830
rect 2050 5796 2056 5830
rect 1938 5757 2056 5796
rect 1938 5723 1944 5757
rect 1978 5723 2016 5757
rect 2050 5723 2056 5757
rect 1938 5683 2056 5723
rect 1938 5649 1944 5683
rect 1978 5649 2016 5683
rect 2050 5649 2056 5683
rect 1938 5609 2056 5649
rect 1938 5575 1944 5609
rect 1978 5575 2016 5609
rect 2050 5575 2056 5609
rect 1938 5535 2056 5575
rect 1938 5501 1944 5535
rect 1978 5501 2016 5535
rect 2050 5501 2056 5535
rect 1938 5461 2056 5501
rect 1938 5427 1944 5461
rect 1978 5427 2016 5461
rect 2050 5427 2056 5461
rect 1938 5387 2056 5427
rect 1938 5353 1944 5387
rect 1978 5353 2016 5387
rect 2050 5353 2056 5387
rect 1938 5313 2056 5353
rect 1938 5279 1944 5313
rect 1978 5279 2016 5313
rect 2050 5279 2056 5313
rect 1938 5239 2056 5279
rect 1938 5205 1944 5239
rect 1978 5205 2016 5239
rect 2050 5205 2056 5239
rect 1938 5165 2056 5205
rect 1938 5131 1944 5165
rect 1978 5131 2016 5165
rect 2050 5131 2056 5165
rect 1938 5091 2056 5131
rect 1938 5057 1944 5091
rect 1978 5057 2016 5091
rect 2050 5057 2056 5091
rect 1938 5017 2056 5057
rect 1938 4983 1944 5017
rect 1978 4983 2016 5017
rect 2050 4983 2056 5017
rect 2249 6589 2791 6607
rect 2249 6555 2255 6589
rect 2289 6555 2327 6589
rect 2361 6568 2791 6589
rect 2361 6555 2679 6568
rect 2249 6534 2679 6555
rect 2713 6534 2751 6568
rect 2785 6534 2791 6568
rect 2249 6516 2791 6534
rect 2249 6482 2255 6516
rect 2289 6482 2327 6516
rect 2361 6495 2791 6516
rect 2361 6482 2679 6495
rect 2249 6461 2679 6482
rect 2713 6461 2751 6495
rect 2785 6461 2791 6495
rect 2249 6443 2791 6461
rect 2249 6409 2255 6443
rect 2289 6409 2327 6443
rect 2361 6422 2791 6443
rect 2361 6409 2679 6422
rect 2249 6370 2679 6409
rect 2249 6336 2255 6370
rect 2289 6336 2327 6370
rect 2361 6336 2679 6370
rect 2249 6297 2679 6336
rect 2249 6263 2255 6297
rect 2289 6263 2327 6297
rect 2361 6263 2679 6297
rect 2249 6224 2679 6263
rect 2249 6190 2255 6224
rect 2289 6190 2327 6224
rect 2361 6190 2679 6224
rect 2249 6151 2679 6190
rect 2249 6117 2255 6151
rect 2289 6117 2327 6151
rect 2361 6117 2679 6151
rect 2249 6078 2679 6117
rect 2249 6044 2255 6078
rect 2289 6044 2327 6078
rect 2361 6044 2679 6078
rect 2249 6005 2679 6044
rect 2249 5971 2255 6005
rect 2289 5971 2327 6005
rect 2361 5971 2679 6005
rect 2249 5932 2679 5971
rect 2249 5898 2255 5932
rect 2289 5898 2327 5932
rect 2361 5898 2679 5932
rect 2249 5859 2679 5898
rect 2249 5825 2255 5859
rect 2289 5825 2327 5859
rect 2361 5825 2679 5859
rect 2249 5786 2679 5825
rect 2249 5752 2255 5786
rect 2289 5752 2327 5786
rect 2361 5752 2679 5786
rect 2249 5713 2679 5752
rect 2249 5679 2255 5713
rect 2289 5679 2327 5713
rect 2361 5679 2679 5713
rect 2249 5640 2679 5679
rect 2249 5606 2255 5640
rect 2289 5606 2327 5640
rect 2361 5606 2679 5640
rect 2249 5567 2679 5606
rect 2249 5533 2255 5567
rect 2289 5533 2327 5567
rect 2361 5533 2679 5567
rect 2249 5494 2679 5533
rect 2249 5460 2255 5494
rect 2289 5460 2327 5494
rect 2361 5460 2679 5494
rect 2249 5421 2679 5460
rect 2249 5387 2255 5421
rect 2289 5387 2327 5421
rect 2361 5387 2679 5421
rect 2249 5380 2679 5387
rect 2785 5380 2791 6422
rect 2950 6714 3068 7376
rect 2950 6680 2956 6714
rect 2990 6680 3028 6714
rect 3062 6680 3068 6714
rect 2950 6641 3068 6680
rect 2950 6607 2956 6641
rect 2990 6607 3028 6641
rect 3062 6607 3068 6641
rect 2950 6568 3068 6607
rect 2950 6534 2956 6568
rect 2990 6534 3028 6568
rect 3062 6534 3068 6568
rect 2950 6495 3068 6534
rect 2950 6461 2956 6495
rect 2990 6461 3028 6495
rect 3062 6461 3068 6495
rect 2950 6422 3068 6461
rect 2950 5896 2956 6422
rect 3062 5896 3068 6422
rect 2950 5830 2956 5844
rect 3062 5830 3068 5844
rect 2950 5764 2956 5778
rect 3062 5764 3068 5778
rect 2950 5698 2956 5712
rect 3062 5698 3068 5712
rect 2950 5632 2956 5646
rect 3062 5632 3068 5646
rect 2950 5566 2956 5580
rect 3062 5566 3068 5580
rect 2950 5499 2956 5514
rect 3062 5499 3068 5514
tri 2791 5380 2858 5447 sw
rect 2950 5432 2956 5447
rect 3062 5432 3068 5447
rect 2249 5377 2858 5380
tri 2858 5377 2861 5380 sw
rect 2249 5374 2861 5377
tri 2861 5374 2864 5377 sw
rect 2249 5368 2864 5374
tri 2864 5368 2870 5374 sw
rect 2950 5368 3068 5380
rect 3279 14338 3293 14390
rect 3781 14720 3899 14726
rect 3833 14668 3847 14720
rect 3781 14654 3899 14668
rect 3833 14602 3847 14654
rect 3781 14588 3899 14602
rect 3833 14536 3847 14588
rect 3781 14522 3899 14536
rect 3833 14470 3847 14522
rect 3781 14456 3899 14470
rect 3833 14404 3847 14456
rect 3781 14390 3899 14404
rect 3227 14323 3233 14338
rect 3267 14323 3305 14338
rect 3339 14323 3345 14338
rect 3279 14271 3293 14323
rect 3227 14267 3345 14271
rect 3227 14256 3233 14267
rect 3267 14256 3305 14267
rect 3339 14256 3345 14267
rect 3279 14204 3293 14256
rect 3227 14189 3345 14204
rect 3227 14155 3233 14189
rect 3267 14155 3305 14189
rect 3339 14155 3345 14189
rect 3227 14111 3345 14155
rect 3227 14077 3233 14111
rect 3267 14077 3305 14111
rect 3339 14077 3345 14111
rect 3227 14033 3345 14077
rect 3227 13999 3233 14033
rect 3267 13999 3305 14033
rect 3339 13999 3345 14033
rect 3227 13955 3345 13999
rect 3227 13921 3233 13955
rect 3267 13921 3305 13955
rect 3339 13921 3345 13955
rect 3227 13877 3345 13921
rect 3227 13843 3233 13877
rect 3267 13843 3305 13877
rect 3339 13843 3345 13877
rect 3227 13799 3345 13843
rect 3227 13765 3233 13799
rect 3267 13765 3305 13799
rect 3339 13765 3345 13799
rect 3227 13722 3345 13765
rect 3227 13688 3233 13722
rect 3267 13688 3305 13722
rect 3339 13688 3345 13722
rect 3227 13645 3345 13688
rect 3227 13611 3233 13645
rect 3267 13611 3305 13645
rect 3339 13611 3345 13645
rect 3227 13568 3345 13611
rect 3227 13534 3233 13568
rect 3267 13534 3305 13568
rect 3339 13534 3345 13568
rect 3227 13491 3345 13534
rect 3227 13457 3233 13491
rect 3267 13457 3305 13491
rect 3339 13457 3345 13491
rect 3227 13414 3345 13457
rect 3227 13380 3233 13414
rect 3267 13380 3305 13414
rect 3339 13380 3345 13414
rect 3227 12720 3345 13380
rect 3279 12668 3293 12720
rect 3227 12654 3345 12668
rect 3279 12602 3293 12654
rect 3227 12588 3345 12602
rect 3279 12536 3293 12588
rect 3227 12534 3233 12536
rect 3267 12534 3305 12536
rect 3339 12534 3345 12536
rect 3227 12522 3345 12534
rect 3279 12470 3293 12522
rect 3227 12461 3233 12470
rect 3267 12461 3305 12470
rect 3339 12461 3345 12470
rect 3227 12456 3345 12461
rect 3279 12422 3293 12456
rect 3227 12390 3233 12404
rect 3339 12390 3345 12404
rect 3227 12323 3233 12338
rect 3339 12323 3345 12338
rect 3227 12256 3233 12271
rect 3339 12256 3345 12271
rect 3227 11380 3233 12204
rect 3339 11380 3345 12204
rect 3227 10724 3345 11380
rect 3279 10672 3293 10724
rect 3227 10658 3345 10672
rect 3279 10606 3293 10658
rect 3227 10592 3345 10606
rect 3279 10540 3293 10592
rect 3227 10534 3233 10540
rect 3267 10534 3305 10540
rect 3339 10534 3345 10540
rect 3227 10526 3345 10534
rect 3279 10474 3293 10526
rect 3227 10461 3233 10474
rect 3267 10461 3305 10474
rect 3339 10461 3345 10474
rect 3227 10460 3345 10461
rect 3279 10422 3293 10460
rect 3227 10394 3233 10408
rect 3339 10394 3345 10408
rect 3227 10327 3233 10342
rect 3339 10327 3345 10342
rect 3227 10260 3233 10275
rect 3339 10260 3345 10275
rect 3227 9380 3233 10208
rect 3339 9380 3345 10208
rect 3227 8720 3345 9380
rect 3279 8668 3293 8720
rect 3227 8654 3345 8668
rect 3279 8602 3293 8654
rect 3227 8588 3345 8602
rect 3279 8536 3293 8588
rect 3227 8534 3233 8536
rect 3267 8534 3305 8536
rect 3339 8534 3345 8536
rect 3227 8522 3345 8534
rect 3279 8470 3293 8522
rect 3227 8461 3233 8470
rect 3267 8461 3305 8470
rect 3339 8461 3345 8470
rect 3227 8456 3345 8461
rect 3279 8422 3293 8456
rect 3227 8390 3233 8404
rect 3339 8390 3345 8404
rect 3227 8323 3233 8338
rect 3339 8323 3345 8338
rect 3227 8256 3233 8271
rect 3339 8256 3345 8271
rect 3227 7380 3233 8204
rect 3339 7380 3345 8204
rect 3227 6724 3345 7380
rect 3279 6672 3293 6724
rect 3227 6658 3345 6672
rect 3279 6606 3293 6658
rect 3227 6592 3345 6606
rect 3279 6540 3293 6592
rect 3227 6534 3233 6540
rect 3267 6534 3305 6540
rect 3339 6534 3345 6540
rect 3227 6526 3345 6534
rect 3279 6474 3293 6526
rect 3227 6461 3233 6474
rect 3267 6461 3305 6474
rect 3339 6461 3345 6474
rect 3227 6460 3345 6461
rect 3279 6422 3293 6460
rect 3227 6394 3233 6408
rect 3339 6394 3345 6408
rect 3227 6327 3233 6342
rect 3339 6327 3345 6342
rect 3227 6260 3233 6275
rect 3339 6260 3345 6275
rect 3227 5380 3233 6208
rect 3339 5380 3345 6208
rect 2249 5362 2870 5368
tri 2870 5362 2876 5368 sw
rect 2249 5348 2876 5362
rect 2249 5314 2255 5348
rect 2289 5314 2327 5348
rect 2361 5338 2876 5348
tri 2876 5338 2900 5362 sw
rect 2361 5314 2900 5338
rect 2249 5304 2900 5314
tri 2900 5304 2934 5338 sw
rect 2249 5289 2934 5304
tri 2934 5289 2949 5304 sw
rect 2249 5274 2949 5289
rect 2249 5240 2255 5274
rect 2289 5240 2327 5274
rect 2361 5271 2949 5274
tri 2949 5271 2967 5289 sw
rect 2361 5265 2967 5271
tri 2967 5265 2973 5271 sw
tri 3221 5265 3227 5271 se
rect 3227 5265 3345 5380
rect 3504 14345 3622 14357
rect 3504 14311 3510 14345
rect 3544 14311 3582 14345
rect 3616 14311 3622 14345
rect 3504 14267 3622 14311
rect 3504 14233 3510 14267
rect 3544 14233 3582 14267
rect 3616 14233 3622 14267
rect 3504 14189 3622 14233
rect 3504 14155 3510 14189
rect 3544 14155 3582 14189
rect 3616 14155 3622 14189
rect 3504 14111 3622 14155
rect 3504 14077 3510 14111
rect 3544 14077 3582 14111
rect 3616 14077 3622 14111
rect 3504 14033 3622 14077
rect 3504 13999 3510 14033
rect 3544 13999 3582 14033
rect 3616 13999 3622 14033
rect 3504 13955 3622 13999
rect 3504 13921 3510 13955
rect 3544 13921 3582 13955
rect 3616 13921 3622 13955
rect 3504 13892 3622 13921
rect 3556 13840 3570 13892
rect 3504 13826 3622 13840
rect 3556 13774 3570 13826
rect 3504 13765 3510 13774
rect 3544 13765 3582 13774
rect 3616 13765 3622 13774
rect 3504 13760 3622 13765
rect 3556 13708 3570 13760
rect 3504 13694 3510 13708
rect 3544 13694 3582 13708
rect 3616 13694 3622 13708
rect 3556 13642 3570 13694
rect 3504 13628 3510 13642
rect 3544 13628 3582 13642
rect 3616 13628 3622 13642
rect 3556 13576 3570 13628
rect 3504 13568 3622 13576
rect 3504 13562 3510 13568
rect 3544 13562 3582 13568
rect 3616 13562 3622 13568
rect 3556 13510 3570 13562
rect 3504 13495 3622 13510
rect 3556 13443 3570 13495
rect 3504 13428 3622 13443
rect 3556 13376 3570 13428
rect 3504 12714 3622 13376
rect 3504 12680 3510 12714
rect 3544 12680 3582 12714
rect 3616 12680 3622 12714
rect 3504 12641 3622 12680
rect 3504 12607 3510 12641
rect 3544 12607 3582 12641
rect 3616 12607 3622 12641
rect 3504 12568 3622 12607
rect 3504 12534 3510 12568
rect 3544 12534 3582 12568
rect 3616 12534 3622 12568
rect 3504 12495 3622 12534
rect 3504 12461 3510 12495
rect 3544 12461 3582 12495
rect 3616 12461 3622 12495
rect 3504 12422 3622 12461
rect 3504 11892 3510 12422
rect 3616 11892 3622 12422
rect 3504 11826 3510 11840
rect 3616 11826 3622 11840
rect 3504 11760 3510 11774
rect 3616 11760 3622 11774
rect 3504 11694 3510 11708
rect 3616 11694 3622 11708
rect 3504 11628 3510 11642
rect 3616 11628 3622 11642
rect 3504 11562 3510 11576
rect 3616 11562 3622 11576
rect 3504 11495 3510 11510
rect 3616 11495 3622 11510
rect 3504 11428 3510 11443
rect 3616 11428 3622 11443
rect 3556 11376 3570 11380
rect 3504 10714 3622 11376
rect 3504 10680 3510 10714
rect 3544 10680 3582 10714
rect 3616 10680 3622 10714
rect 3504 10641 3622 10680
rect 3504 10607 3510 10641
rect 3544 10607 3582 10641
rect 3616 10607 3622 10641
rect 3504 10568 3622 10607
rect 3504 10534 3510 10568
rect 3544 10534 3582 10568
rect 3616 10534 3622 10568
rect 3504 10495 3622 10534
rect 3504 10461 3510 10495
rect 3544 10461 3582 10495
rect 3616 10461 3622 10495
rect 3504 10422 3622 10461
rect 3504 9896 3510 10422
rect 3616 9896 3622 10422
rect 3504 9830 3510 9844
rect 3616 9830 3622 9844
rect 3504 9764 3510 9778
rect 3616 9764 3622 9778
rect 3504 9698 3510 9712
rect 3616 9698 3622 9712
rect 3504 9632 3510 9646
rect 3616 9632 3622 9646
rect 3504 9566 3510 9580
rect 3616 9566 3622 9580
rect 3504 9499 3510 9514
rect 3616 9499 3622 9514
rect 3504 9432 3510 9447
rect 3616 9432 3622 9447
rect 3504 8714 3622 9380
rect 3504 8680 3510 8714
rect 3544 8680 3582 8714
rect 3616 8680 3622 8714
rect 3504 8641 3622 8680
rect 3504 8607 3510 8641
rect 3544 8607 3582 8641
rect 3616 8607 3622 8641
rect 3504 8568 3622 8607
rect 3504 8534 3510 8568
rect 3544 8534 3582 8568
rect 3616 8534 3622 8568
rect 3504 8495 3622 8534
rect 3504 8461 3510 8495
rect 3544 8461 3582 8495
rect 3616 8461 3622 8495
rect 3504 8422 3622 8461
rect 3504 7892 3510 8422
rect 3616 7892 3622 8422
rect 3504 7826 3510 7840
rect 3616 7826 3622 7840
rect 3504 7760 3510 7774
rect 3616 7760 3622 7774
rect 3504 7694 3510 7708
rect 3616 7694 3622 7708
rect 3504 7628 3510 7642
rect 3616 7628 3622 7642
rect 3504 7562 3510 7576
rect 3616 7562 3622 7576
rect 3504 7495 3510 7510
rect 3616 7495 3622 7510
rect 3504 7428 3510 7443
rect 3616 7428 3622 7443
rect 3556 7376 3570 7380
rect 3504 6714 3622 7376
rect 3504 6680 3510 6714
rect 3544 6680 3582 6714
rect 3616 6680 3622 6714
rect 3504 6641 3622 6680
rect 3504 6607 3510 6641
rect 3544 6607 3582 6641
rect 3616 6607 3622 6641
rect 3504 6568 3622 6607
rect 3504 6534 3510 6568
rect 3544 6534 3582 6568
rect 3616 6534 3622 6568
rect 3504 6495 3622 6534
rect 3504 6461 3510 6495
rect 3544 6461 3582 6495
rect 3616 6461 3622 6495
rect 3504 6422 3622 6461
rect 3504 5896 3510 6422
rect 3616 5896 3622 6422
rect 3504 5830 3510 5844
rect 3616 5830 3622 5844
rect 3504 5764 3510 5778
rect 3616 5764 3622 5778
rect 3504 5698 3510 5712
rect 3616 5698 3622 5712
rect 3504 5632 3510 5646
rect 3616 5632 3622 5646
rect 3504 5566 3510 5580
rect 3616 5566 3622 5580
rect 3504 5499 3510 5514
rect 3616 5499 3622 5514
rect 3504 5432 3510 5447
rect 3616 5432 3622 5447
rect 3504 5368 3622 5380
rect 3833 14338 3847 14390
rect 4335 14720 4453 14726
rect 4387 14668 4401 14720
rect 4335 14654 4453 14668
rect 4387 14602 4401 14654
rect 4335 14588 4453 14602
rect 4387 14536 4401 14588
rect 4335 14522 4453 14536
rect 4387 14470 4401 14522
rect 4335 14456 4453 14470
rect 4387 14404 4401 14456
rect 4335 14390 4453 14404
rect 3781 14323 3787 14338
rect 3821 14323 3859 14338
rect 3893 14323 3899 14338
rect 3833 14271 3847 14323
rect 3781 14267 3899 14271
rect 3781 14256 3787 14267
rect 3821 14256 3859 14267
rect 3893 14256 3899 14267
rect 3833 14204 3847 14256
rect 3781 14189 3899 14204
rect 3781 14155 3787 14189
rect 3821 14155 3859 14189
rect 3893 14155 3899 14189
rect 3781 14111 3899 14155
rect 3781 14077 3787 14111
rect 3821 14077 3859 14111
rect 3893 14077 3899 14111
rect 3781 14033 3899 14077
rect 3781 13999 3787 14033
rect 3821 13999 3859 14033
rect 3893 13999 3899 14033
rect 3781 13955 3899 13999
rect 3781 13921 3787 13955
rect 3821 13921 3859 13955
rect 3893 13921 3899 13955
rect 3781 13877 3899 13921
rect 3781 13843 3787 13877
rect 3821 13843 3859 13877
rect 3893 13843 3899 13877
rect 3781 13799 3899 13843
rect 3781 13765 3787 13799
rect 3821 13765 3859 13799
rect 3893 13765 3899 13799
rect 3781 13722 3899 13765
rect 3781 13688 3787 13722
rect 3821 13688 3859 13722
rect 3893 13688 3899 13722
rect 3781 13645 3899 13688
rect 3781 13611 3787 13645
rect 3821 13611 3859 13645
rect 3893 13611 3899 13645
rect 3781 13568 3899 13611
rect 3781 13534 3787 13568
rect 3821 13534 3859 13568
rect 3893 13534 3899 13568
rect 3781 13491 3899 13534
rect 3781 13457 3787 13491
rect 3821 13457 3859 13491
rect 3893 13457 3899 13491
rect 3781 13414 3899 13457
rect 3781 13380 3787 13414
rect 3821 13380 3859 13414
rect 3893 13380 3899 13414
rect 3781 12720 3899 13380
rect 3833 12668 3847 12720
rect 3781 12654 3899 12668
rect 3833 12602 3847 12654
rect 3781 12588 3899 12602
rect 3833 12536 3847 12588
rect 3781 12534 3787 12536
rect 3821 12534 3859 12536
rect 3893 12534 3899 12536
rect 3781 12522 3899 12534
rect 3833 12470 3847 12522
rect 3781 12461 3787 12470
rect 3821 12461 3859 12470
rect 3893 12461 3899 12470
rect 3781 12456 3899 12461
rect 3833 12422 3847 12456
rect 3781 12390 3787 12404
rect 3893 12390 3899 12404
rect 3781 12323 3787 12338
rect 3893 12323 3899 12338
rect 3781 12256 3787 12271
rect 3893 12256 3899 12271
rect 3781 11380 3787 12204
rect 3893 11380 3899 12204
rect 3781 10724 3899 11380
rect 3833 10672 3847 10724
rect 3781 10658 3899 10672
rect 3833 10606 3847 10658
rect 3781 10592 3899 10606
rect 3833 10540 3847 10592
rect 3781 10534 3787 10540
rect 3821 10534 3859 10540
rect 3893 10534 3899 10540
rect 3781 10526 3899 10534
rect 3833 10474 3847 10526
rect 3781 10461 3787 10474
rect 3821 10461 3859 10474
rect 3893 10461 3899 10474
rect 3781 10460 3899 10461
rect 3833 10422 3847 10460
rect 3781 10394 3787 10408
rect 3893 10394 3899 10408
rect 3781 10327 3787 10342
rect 3893 10327 3899 10342
rect 3781 10260 3787 10275
rect 3893 10260 3899 10275
rect 3781 9380 3787 10208
rect 3893 9380 3899 10208
rect 3781 8720 3899 9380
rect 3833 8668 3847 8720
rect 3781 8654 3899 8668
rect 3833 8602 3847 8654
rect 3781 8588 3899 8602
rect 3833 8536 3847 8588
rect 3781 8534 3787 8536
rect 3821 8534 3859 8536
rect 3893 8534 3899 8536
rect 3781 8522 3899 8534
rect 3833 8470 3847 8522
rect 3781 8461 3787 8470
rect 3821 8461 3859 8470
rect 3893 8461 3899 8470
rect 3781 8456 3899 8461
rect 3833 8422 3847 8456
rect 3781 8390 3787 8404
rect 3893 8390 3899 8404
rect 3781 8323 3787 8338
rect 3893 8323 3899 8338
rect 3781 8256 3787 8271
rect 3893 8256 3899 8271
rect 3781 7380 3787 8204
rect 3893 7380 3899 8204
rect 3781 6724 3899 7380
rect 3833 6672 3847 6724
rect 3781 6658 3899 6672
rect 3833 6606 3847 6658
rect 3781 6592 3899 6606
rect 3833 6540 3847 6592
rect 3781 6534 3787 6540
rect 3821 6534 3859 6540
rect 3893 6534 3899 6540
rect 3781 6526 3899 6534
rect 3833 6474 3847 6526
rect 3781 6461 3787 6474
rect 3821 6461 3859 6474
rect 3893 6461 3899 6474
rect 3781 6460 3899 6461
rect 3833 6422 3847 6460
rect 3781 6394 3787 6408
rect 3893 6394 3899 6408
rect 3781 6327 3787 6342
rect 3893 6327 3899 6342
rect 3781 6260 3787 6275
rect 3893 6260 3899 6275
rect 3781 5380 3787 6208
rect 3893 5380 3899 6208
tri 3345 5265 3351 5271 sw
tri 3775 5265 3781 5271 se
rect 3781 5265 3899 5380
rect 4058 14345 4176 14357
rect 4058 14311 4064 14345
rect 4098 14311 4136 14345
rect 4170 14311 4176 14345
rect 4058 14267 4176 14311
rect 4058 14233 4064 14267
rect 4098 14233 4136 14267
rect 4170 14233 4176 14267
rect 4058 14189 4176 14233
rect 4058 14155 4064 14189
rect 4098 14155 4136 14189
rect 4170 14155 4176 14189
rect 4058 14111 4176 14155
rect 4058 14077 4064 14111
rect 4098 14077 4136 14111
rect 4170 14077 4176 14111
rect 4058 14033 4176 14077
rect 4058 13999 4064 14033
rect 4098 13999 4136 14033
rect 4170 13999 4176 14033
rect 4058 13955 4176 13999
rect 4058 13921 4064 13955
rect 4098 13921 4136 13955
rect 4170 13921 4176 13955
rect 4058 13892 4176 13921
rect 4110 13840 4124 13892
rect 4058 13826 4176 13840
rect 4110 13774 4124 13826
rect 4058 13765 4064 13774
rect 4098 13765 4136 13774
rect 4170 13765 4176 13774
rect 4058 13760 4176 13765
rect 4110 13708 4124 13760
rect 4058 13694 4064 13708
rect 4098 13694 4136 13708
rect 4170 13694 4176 13708
rect 4110 13642 4124 13694
rect 4058 13628 4064 13642
rect 4098 13628 4136 13642
rect 4170 13628 4176 13642
rect 4110 13576 4124 13628
rect 4058 13568 4176 13576
rect 4058 13562 4064 13568
rect 4098 13562 4136 13568
rect 4170 13562 4176 13568
rect 4110 13510 4124 13562
rect 4058 13495 4176 13510
rect 4110 13443 4124 13495
rect 4058 13428 4176 13443
rect 4110 13376 4124 13428
rect 4058 12714 4176 13376
rect 4058 12680 4064 12714
rect 4098 12680 4136 12714
rect 4170 12680 4176 12714
rect 4058 12641 4176 12680
rect 4058 12607 4064 12641
rect 4098 12607 4136 12641
rect 4170 12607 4176 12641
rect 4058 12568 4176 12607
rect 4058 12534 4064 12568
rect 4098 12534 4136 12568
rect 4170 12534 4176 12568
rect 4058 12495 4176 12534
rect 4058 12461 4064 12495
rect 4098 12461 4136 12495
rect 4170 12461 4176 12495
rect 4058 12422 4176 12461
rect 4058 11892 4064 12422
rect 4170 11892 4176 12422
rect 4058 11826 4064 11840
rect 4170 11826 4176 11840
rect 4058 11760 4064 11774
rect 4170 11760 4176 11774
rect 4058 11694 4064 11708
rect 4170 11694 4176 11708
rect 4058 11628 4064 11642
rect 4170 11628 4176 11642
rect 4058 11562 4064 11576
rect 4170 11562 4176 11576
rect 4058 11495 4064 11510
rect 4170 11495 4176 11510
rect 4058 11428 4064 11443
rect 4170 11428 4176 11443
rect 4110 11376 4124 11380
rect 4058 10714 4176 11376
rect 4058 10680 4064 10714
rect 4098 10680 4136 10714
rect 4170 10680 4176 10714
rect 4058 10641 4176 10680
rect 4058 10607 4064 10641
rect 4098 10607 4136 10641
rect 4170 10607 4176 10641
rect 4058 10568 4176 10607
rect 4058 10534 4064 10568
rect 4098 10534 4136 10568
rect 4170 10534 4176 10568
rect 4058 10495 4176 10534
rect 4058 10461 4064 10495
rect 4098 10461 4136 10495
rect 4170 10461 4176 10495
rect 4058 10422 4176 10461
rect 4058 9896 4064 10422
rect 4170 9896 4176 10422
rect 4058 9830 4064 9844
rect 4170 9830 4176 9844
rect 4058 9764 4064 9778
rect 4170 9764 4176 9778
rect 4058 9698 4064 9712
rect 4170 9698 4176 9712
rect 4058 9632 4064 9646
rect 4170 9632 4176 9646
rect 4058 9566 4064 9580
rect 4170 9566 4176 9580
rect 4058 9499 4064 9514
rect 4170 9499 4176 9514
rect 4058 9432 4064 9447
rect 4170 9432 4176 9447
rect 4058 8714 4176 9380
rect 4058 8680 4064 8714
rect 4098 8680 4136 8714
rect 4170 8680 4176 8714
rect 4058 8641 4176 8680
rect 4058 8607 4064 8641
rect 4098 8607 4136 8641
rect 4170 8607 4176 8641
rect 4058 8568 4176 8607
rect 4058 8534 4064 8568
rect 4098 8534 4136 8568
rect 4170 8534 4176 8568
rect 4058 8495 4176 8534
rect 4058 8461 4064 8495
rect 4098 8461 4136 8495
rect 4170 8461 4176 8495
rect 4058 8422 4176 8461
rect 4058 7892 4064 8422
rect 4170 7892 4176 8422
rect 4058 7826 4064 7840
rect 4170 7826 4176 7840
rect 4058 7760 4064 7774
rect 4170 7760 4176 7774
rect 4058 7694 4064 7708
rect 4170 7694 4176 7708
rect 4058 7628 4064 7642
rect 4170 7628 4176 7642
rect 4058 7562 4064 7576
rect 4170 7562 4176 7576
rect 4058 7495 4064 7510
rect 4170 7495 4176 7510
rect 4058 7428 4064 7443
rect 4170 7428 4176 7443
rect 4110 7376 4124 7380
rect 4058 6714 4176 7376
rect 4058 6680 4064 6714
rect 4098 6680 4136 6714
rect 4170 6680 4176 6714
rect 4058 6641 4176 6680
rect 4058 6607 4064 6641
rect 4098 6607 4136 6641
rect 4170 6607 4176 6641
rect 4058 6568 4176 6607
rect 4058 6534 4064 6568
rect 4098 6534 4136 6568
rect 4170 6534 4176 6568
rect 4058 6495 4176 6534
rect 4058 6461 4064 6495
rect 4098 6461 4136 6495
rect 4170 6461 4176 6495
rect 4058 6422 4176 6461
rect 4058 5896 4064 6422
rect 4170 5896 4176 6422
rect 4058 5830 4064 5844
rect 4170 5830 4176 5844
rect 4058 5764 4064 5778
rect 4170 5764 4176 5778
rect 4058 5698 4064 5712
rect 4170 5698 4176 5712
rect 4058 5632 4064 5646
rect 4170 5632 4176 5646
rect 4058 5566 4064 5580
rect 4170 5566 4176 5580
rect 4058 5499 4064 5514
rect 4170 5499 4176 5514
rect 4058 5432 4064 5447
rect 4170 5432 4176 5447
rect 4058 5368 4176 5380
rect 4387 14338 4401 14390
rect 4889 14720 5007 14726
rect 4941 14668 4955 14720
rect 4889 14654 5007 14668
rect 4941 14602 4955 14654
rect 4889 14588 5007 14602
rect 4941 14536 4955 14588
rect 4889 14522 5007 14536
rect 4941 14470 4955 14522
rect 4889 14456 5007 14470
rect 4941 14404 4955 14456
rect 4889 14390 5007 14404
rect 4335 14323 4341 14338
rect 4375 14323 4413 14338
rect 4447 14323 4453 14338
rect 4387 14271 4401 14323
rect 4335 14267 4453 14271
rect 4335 14256 4341 14267
rect 4375 14256 4413 14267
rect 4447 14256 4453 14267
rect 4387 14204 4401 14256
rect 4335 14189 4453 14204
rect 4335 14155 4341 14189
rect 4375 14155 4413 14189
rect 4447 14155 4453 14189
rect 4335 14111 4453 14155
rect 4335 14077 4341 14111
rect 4375 14077 4413 14111
rect 4447 14077 4453 14111
rect 4335 14033 4453 14077
rect 4335 13999 4341 14033
rect 4375 13999 4413 14033
rect 4447 13999 4453 14033
rect 4335 13955 4453 13999
rect 4335 13921 4341 13955
rect 4375 13921 4413 13955
rect 4447 13921 4453 13955
rect 4335 13877 4453 13921
rect 4335 13843 4341 13877
rect 4375 13843 4413 13877
rect 4447 13843 4453 13877
rect 4335 13799 4453 13843
rect 4335 13765 4341 13799
rect 4375 13765 4413 13799
rect 4447 13765 4453 13799
rect 4335 13722 4453 13765
rect 4335 13688 4341 13722
rect 4375 13688 4413 13722
rect 4447 13688 4453 13722
rect 4335 13645 4453 13688
rect 4335 13611 4341 13645
rect 4375 13611 4413 13645
rect 4447 13611 4453 13645
rect 4335 13568 4453 13611
rect 4335 13534 4341 13568
rect 4375 13534 4413 13568
rect 4447 13534 4453 13568
rect 4335 13491 4453 13534
rect 4335 13457 4341 13491
rect 4375 13457 4413 13491
rect 4447 13457 4453 13491
rect 4335 13414 4453 13457
rect 4335 13380 4341 13414
rect 4375 13380 4413 13414
rect 4447 13380 4453 13414
rect 4335 12720 4453 13380
rect 4387 12668 4401 12720
rect 4335 12654 4453 12668
rect 4387 12602 4401 12654
rect 4335 12588 4453 12602
rect 4387 12536 4401 12588
rect 4335 12534 4341 12536
rect 4375 12534 4413 12536
rect 4447 12534 4453 12536
rect 4335 12522 4453 12534
rect 4387 12470 4401 12522
rect 4335 12461 4341 12470
rect 4375 12461 4413 12470
rect 4447 12461 4453 12470
rect 4335 12456 4453 12461
rect 4387 12422 4401 12456
rect 4335 12390 4341 12404
rect 4447 12390 4453 12404
rect 4335 12323 4341 12338
rect 4447 12323 4453 12338
rect 4335 12256 4341 12271
rect 4447 12256 4453 12271
rect 4335 11380 4341 12204
rect 4447 11380 4453 12204
rect 4335 10724 4453 11380
rect 4387 10672 4401 10724
rect 4335 10658 4453 10672
rect 4387 10606 4401 10658
rect 4335 10592 4453 10606
rect 4387 10540 4401 10592
rect 4335 10534 4341 10540
rect 4375 10534 4413 10540
rect 4447 10534 4453 10540
rect 4335 10526 4453 10534
rect 4387 10474 4401 10526
rect 4335 10461 4341 10474
rect 4375 10461 4413 10474
rect 4447 10461 4453 10474
rect 4335 10460 4453 10461
rect 4387 10422 4401 10460
rect 4335 10394 4341 10408
rect 4447 10394 4453 10408
rect 4335 10327 4341 10342
rect 4447 10327 4453 10342
rect 4335 10260 4341 10275
rect 4447 10260 4453 10275
rect 4335 9380 4341 10208
rect 4447 9380 4453 10208
rect 4335 8720 4453 9380
rect 4387 8668 4401 8720
rect 4335 8654 4453 8668
rect 4387 8602 4401 8654
rect 4335 8588 4453 8602
rect 4387 8536 4401 8588
rect 4335 8534 4341 8536
rect 4375 8534 4413 8536
rect 4447 8534 4453 8536
rect 4335 8522 4453 8534
rect 4387 8470 4401 8522
rect 4335 8461 4341 8470
rect 4375 8461 4413 8470
rect 4447 8461 4453 8470
rect 4335 8456 4453 8461
rect 4387 8422 4401 8456
rect 4335 8390 4341 8404
rect 4447 8390 4453 8404
rect 4335 8323 4341 8338
rect 4447 8323 4453 8338
rect 4335 8256 4341 8271
rect 4447 8256 4453 8271
rect 4335 7380 4341 8204
rect 4447 7380 4453 8204
rect 4335 6724 4453 7380
rect 4387 6672 4401 6724
rect 4335 6658 4453 6672
rect 4387 6606 4401 6658
rect 4335 6592 4453 6606
rect 4387 6540 4401 6592
rect 4335 6534 4341 6540
rect 4375 6534 4413 6540
rect 4447 6534 4453 6540
rect 4335 6526 4453 6534
rect 4387 6474 4401 6526
rect 4335 6461 4341 6474
rect 4375 6461 4413 6474
rect 4447 6461 4453 6474
rect 4335 6460 4453 6461
rect 4387 6422 4401 6460
rect 4335 6394 4341 6408
rect 4447 6394 4453 6408
rect 4335 6327 4341 6342
rect 4447 6327 4453 6342
rect 4335 6260 4341 6275
rect 4447 6260 4453 6275
rect 4335 5380 4341 6208
rect 4447 5380 4453 6208
tri 3899 5265 3905 5271 sw
tri 4329 5265 4335 5271 se
rect 4335 5265 4453 5380
rect 4612 14345 4730 14357
rect 4612 14311 4618 14345
rect 4652 14311 4690 14345
rect 4724 14311 4730 14345
rect 4612 14267 4730 14311
rect 4612 14233 4618 14267
rect 4652 14233 4690 14267
rect 4724 14233 4730 14267
rect 4612 14189 4730 14233
rect 4612 14155 4618 14189
rect 4652 14155 4690 14189
rect 4724 14155 4730 14189
rect 4612 14111 4730 14155
rect 4612 14077 4618 14111
rect 4652 14077 4690 14111
rect 4724 14077 4730 14111
rect 4612 14033 4730 14077
rect 4612 13999 4618 14033
rect 4652 13999 4690 14033
rect 4724 13999 4730 14033
rect 4612 13955 4730 13999
rect 4612 13921 4618 13955
rect 4652 13921 4690 13955
rect 4724 13921 4730 13955
rect 4612 13892 4730 13921
rect 4664 13840 4678 13892
rect 4612 13826 4730 13840
rect 4664 13774 4678 13826
rect 4612 13765 4618 13774
rect 4652 13765 4690 13774
rect 4724 13765 4730 13774
rect 4612 13760 4730 13765
rect 4664 13708 4678 13760
rect 4612 13694 4618 13708
rect 4652 13694 4690 13708
rect 4724 13694 4730 13708
rect 4664 13642 4678 13694
rect 4612 13628 4618 13642
rect 4652 13628 4690 13642
rect 4724 13628 4730 13642
rect 4664 13576 4678 13628
rect 4612 13568 4730 13576
rect 4612 13562 4618 13568
rect 4652 13562 4690 13568
rect 4724 13562 4730 13568
rect 4664 13510 4678 13562
rect 4612 13495 4730 13510
rect 4664 13443 4678 13495
rect 4612 13428 4730 13443
rect 4664 13376 4678 13428
rect 4612 12714 4730 13376
rect 4612 12680 4618 12714
rect 4652 12680 4690 12714
rect 4724 12680 4730 12714
rect 4612 12641 4730 12680
rect 4612 12607 4618 12641
rect 4652 12607 4690 12641
rect 4724 12607 4730 12641
rect 4612 12568 4730 12607
rect 4612 12534 4618 12568
rect 4652 12534 4690 12568
rect 4724 12534 4730 12568
rect 4612 12495 4730 12534
rect 4612 12461 4618 12495
rect 4652 12461 4690 12495
rect 4724 12461 4730 12495
rect 4612 12422 4730 12461
rect 4612 11892 4618 12422
rect 4724 11892 4730 12422
rect 4612 11826 4618 11840
rect 4724 11826 4730 11840
rect 4612 11760 4618 11774
rect 4724 11760 4730 11774
rect 4612 11694 4618 11708
rect 4724 11694 4730 11708
rect 4612 11628 4618 11642
rect 4724 11628 4730 11642
rect 4612 11562 4618 11576
rect 4724 11562 4730 11576
rect 4612 11495 4618 11510
rect 4724 11495 4730 11510
rect 4612 11428 4618 11443
rect 4724 11428 4730 11443
rect 4664 11376 4678 11380
rect 4612 10714 4730 11376
rect 4612 10680 4618 10714
rect 4652 10680 4690 10714
rect 4724 10680 4730 10714
rect 4612 10641 4730 10680
rect 4612 10607 4618 10641
rect 4652 10607 4690 10641
rect 4724 10607 4730 10641
rect 4612 10568 4730 10607
rect 4612 10534 4618 10568
rect 4652 10534 4690 10568
rect 4724 10534 4730 10568
rect 4612 10495 4730 10534
rect 4612 10461 4618 10495
rect 4652 10461 4690 10495
rect 4724 10461 4730 10495
rect 4612 10422 4730 10461
rect 4612 9896 4618 10422
rect 4724 9896 4730 10422
rect 4612 9830 4618 9844
rect 4724 9830 4730 9844
rect 4612 9764 4618 9778
rect 4724 9764 4730 9778
rect 4612 9698 4618 9712
rect 4724 9698 4730 9712
rect 4612 9632 4618 9646
rect 4724 9632 4730 9646
rect 4612 9566 4618 9580
rect 4724 9566 4730 9580
rect 4612 9499 4618 9514
rect 4724 9499 4730 9514
rect 4612 9432 4618 9447
rect 4724 9432 4730 9447
rect 4612 8714 4730 9380
rect 4612 8680 4618 8714
rect 4652 8680 4690 8714
rect 4724 8680 4730 8714
rect 4612 8641 4730 8680
rect 4612 8607 4618 8641
rect 4652 8607 4690 8641
rect 4724 8607 4730 8641
rect 4612 8568 4730 8607
rect 4612 8534 4618 8568
rect 4652 8534 4690 8568
rect 4724 8534 4730 8568
rect 4612 8495 4730 8534
rect 4612 8461 4618 8495
rect 4652 8461 4690 8495
rect 4724 8461 4730 8495
rect 4612 8422 4730 8461
rect 4612 7892 4618 8422
rect 4724 7892 4730 8422
rect 4612 7826 4618 7840
rect 4724 7826 4730 7840
rect 4612 7760 4618 7774
rect 4724 7760 4730 7774
rect 4612 7694 4618 7708
rect 4724 7694 4730 7708
rect 4612 7628 4618 7642
rect 4724 7628 4730 7642
rect 4612 7562 4618 7576
rect 4724 7562 4730 7576
rect 4612 7495 4618 7510
rect 4724 7495 4730 7510
rect 4612 7428 4618 7443
rect 4724 7428 4730 7443
rect 4664 7376 4678 7380
rect 4612 6714 4730 7376
rect 4612 6680 4618 6714
rect 4652 6680 4690 6714
rect 4724 6680 4730 6714
rect 4612 6641 4730 6680
rect 4612 6607 4618 6641
rect 4652 6607 4690 6641
rect 4724 6607 4730 6641
rect 4612 6568 4730 6607
rect 4612 6534 4618 6568
rect 4652 6534 4690 6568
rect 4724 6534 4730 6568
rect 4612 6495 4730 6534
rect 4612 6461 4618 6495
rect 4652 6461 4690 6495
rect 4724 6461 4730 6495
rect 4612 6422 4730 6461
rect 4612 5896 4618 6422
rect 4724 5896 4730 6422
rect 4612 5830 4618 5844
rect 4724 5830 4730 5844
rect 4612 5764 4618 5778
rect 4724 5764 4730 5778
rect 4612 5698 4618 5712
rect 4724 5698 4730 5712
rect 4612 5632 4618 5646
rect 4724 5632 4730 5646
rect 4612 5566 4618 5580
rect 4724 5566 4730 5580
rect 4612 5499 4618 5514
rect 4724 5499 4730 5514
rect 4612 5432 4618 5447
rect 4724 5432 4730 5447
rect 4612 5368 4730 5380
rect 4941 14338 4955 14390
rect 5443 14720 5561 14726
rect 5495 14668 5509 14720
rect 5443 14654 5561 14668
rect 5495 14602 5509 14654
rect 5443 14588 5561 14602
rect 5495 14536 5509 14588
rect 5443 14522 5561 14536
rect 5495 14470 5509 14522
rect 5443 14456 5561 14470
rect 5495 14404 5509 14456
rect 5443 14390 5561 14404
rect 4889 14323 4895 14338
rect 4929 14323 4967 14338
rect 5001 14323 5007 14338
rect 4941 14271 4955 14323
rect 4889 14267 5007 14271
rect 4889 14256 4895 14267
rect 4929 14256 4967 14267
rect 5001 14256 5007 14267
rect 4941 14204 4955 14256
rect 4889 14189 5007 14204
rect 4889 14155 4895 14189
rect 4929 14155 4967 14189
rect 5001 14155 5007 14189
rect 4889 14111 5007 14155
rect 4889 14077 4895 14111
rect 4929 14077 4967 14111
rect 5001 14077 5007 14111
rect 4889 14033 5007 14077
rect 4889 13999 4895 14033
rect 4929 13999 4967 14033
rect 5001 13999 5007 14033
rect 4889 13955 5007 13999
rect 4889 13921 4895 13955
rect 4929 13921 4967 13955
rect 5001 13921 5007 13955
rect 4889 13877 5007 13921
rect 4889 13843 4895 13877
rect 4929 13843 4967 13877
rect 5001 13843 5007 13877
rect 4889 13799 5007 13843
rect 4889 13765 4895 13799
rect 4929 13765 4967 13799
rect 5001 13765 5007 13799
rect 4889 13722 5007 13765
rect 4889 13688 4895 13722
rect 4929 13688 4967 13722
rect 5001 13688 5007 13722
rect 4889 13645 5007 13688
rect 4889 13611 4895 13645
rect 4929 13611 4967 13645
rect 5001 13611 5007 13645
rect 4889 13568 5007 13611
rect 4889 13534 4895 13568
rect 4929 13534 4967 13568
rect 5001 13534 5007 13568
rect 4889 13491 5007 13534
rect 4889 13457 4895 13491
rect 4929 13457 4967 13491
rect 5001 13457 5007 13491
rect 4889 13414 5007 13457
rect 4889 13380 4895 13414
rect 4929 13380 4967 13414
rect 5001 13380 5007 13414
rect 4889 12720 5007 13380
rect 4941 12668 4955 12720
rect 4889 12654 5007 12668
rect 4941 12602 4955 12654
rect 4889 12588 5007 12602
rect 4941 12536 4955 12588
rect 4889 12534 4895 12536
rect 4929 12534 4967 12536
rect 5001 12534 5007 12536
rect 4889 12522 5007 12534
rect 4941 12470 4955 12522
rect 4889 12461 4895 12470
rect 4929 12461 4967 12470
rect 5001 12461 5007 12470
rect 4889 12456 5007 12461
rect 4941 12422 4955 12456
rect 4889 12390 4895 12404
rect 5001 12390 5007 12404
rect 4889 12323 4895 12338
rect 5001 12323 5007 12338
rect 4889 12256 4895 12271
rect 5001 12256 5007 12271
rect 4889 11380 4895 12204
rect 5001 11380 5007 12204
rect 4889 10724 5007 11380
rect 4941 10672 4955 10724
rect 4889 10658 5007 10672
rect 4941 10606 4955 10658
rect 4889 10592 5007 10606
rect 4941 10540 4955 10592
rect 4889 10534 4895 10540
rect 4929 10534 4967 10540
rect 5001 10534 5007 10540
rect 4889 10526 5007 10534
rect 4941 10474 4955 10526
rect 4889 10461 4895 10474
rect 4929 10461 4967 10474
rect 5001 10461 5007 10474
rect 4889 10460 5007 10461
rect 4941 10422 4955 10460
rect 4889 10394 4895 10408
rect 5001 10394 5007 10408
rect 4889 10327 4895 10342
rect 5001 10327 5007 10342
rect 4889 10260 4895 10275
rect 5001 10260 5007 10275
rect 4889 9380 4895 10208
rect 5001 9380 5007 10208
rect 4889 8720 5007 9380
rect 4941 8668 4955 8720
rect 4889 8654 5007 8668
rect 4941 8602 4955 8654
rect 4889 8588 5007 8602
rect 4941 8536 4955 8588
rect 4889 8534 4895 8536
rect 4929 8534 4967 8536
rect 5001 8534 5007 8536
rect 4889 8522 5007 8534
rect 4941 8470 4955 8522
rect 4889 8461 4895 8470
rect 4929 8461 4967 8470
rect 5001 8461 5007 8470
rect 4889 8456 5007 8461
rect 4941 8422 4955 8456
rect 4889 8390 4895 8404
rect 5001 8390 5007 8404
rect 4889 8323 4895 8338
rect 5001 8323 5007 8338
rect 4889 8256 4895 8271
rect 5001 8256 5007 8271
rect 4889 7380 4895 8204
rect 5001 7380 5007 8204
rect 4889 6724 5007 7380
rect 4941 6672 4955 6724
rect 4889 6658 5007 6672
rect 4941 6606 4955 6658
rect 4889 6592 5007 6606
rect 4941 6540 4955 6592
rect 4889 6534 4895 6540
rect 4929 6534 4967 6540
rect 5001 6534 5007 6540
rect 4889 6526 5007 6534
rect 4941 6474 4955 6526
rect 4889 6461 4895 6474
rect 4929 6461 4967 6474
rect 5001 6461 5007 6474
rect 4889 6460 5007 6461
rect 4941 6422 4955 6460
rect 4889 6394 4895 6408
rect 5001 6394 5007 6408
rect 4889 6327 4895 6342
rect 5001 6327 5007 6342
rect 4889 6260 4895 6275
rect 5001 6260 5007 6275
rect 4889 5380 4895 6208
rect 5001 5380 5007 6208
tri 4453 5265 4459 5271 sw
tri 4883 5265 4889 5271 se
rect 4889 5265 5007 5380
rect 5166 14345 5284 14357
rect 5166 14311 5172 14345
rect 5206 14311 5244 14345
rect 5278 14311 5284 14345
rect 5166 14267 5284 14311
rect 5166 14233 5172 14267
rect 5206 14233 5244 14267
rect 5278 14233 5284 14267
rect 5166 14189 5284 14233
rect 5166 14155 5172 14189
rect 5206 14155 5244 14189
rect 5278 14155 5284 14189
rect 5166 14111 5284 14155
rect 5166 14077 5172 14111
rect 5206 14077 5244 14111
rect 5278 14077 5284 14111
rect 5166 14033 5284 14077
rect 5166 13999 5172 14033
rect 5206 13999 5244 14033
rect 5278 13999 5284 14033
rect 5166 13955 5284 13999
rect 5166 13921 5172 13955
rect 5206 13921 5244 13955
rect 5278 13921 5284 13955
rect 5166 13892 5284 13921
rect 5218 13840 5232 13892
rect 5166 13826 5284 13840
rect 5218 13774 5232 13826
rect 5166 13765 5172 13774
rect 5206 13765 5244 13774
rect 5278 13765 5284 13774
rect 5166 13760 5284 13765
rect 5218 13708 5232 13760
rect 5166 13694 5172 13708
rect 5206 13694 5244 13708
rect 5278 13694 5284 13708
rect 5218 13642 5232 13694
rect 5166 13628 5172 13642
rect 5206 13628 5244 13642
rect 5278 13628 5284 13642
rect 5218 13576 5232 13628
rect 5166 13568 5284 13576
rect 5166 13562 5172 13568
rect 5206 13562 5244 13568
rect 5278 13562 5284 13568
rect 5218 13510 5232 13562
rect 5166 13495 5284 13510
rect 5218 13443 5232 13495
rect 5166 13428 5284 13443
rect 5218 13376 5232 13428
rect 5166 12714 5284 13376
rect 5166 12680 5172 12714
rect 5206 12680 5244 12714
rect 5278 12680 5284 12714
rect 5166 12641 5284 12680
rect 5166 12607 5172 12641
rect 5206 12607 5244 12641
rect 5278 12607 5284 12641
rect 5166 12568 5284 12607
rect 5166 12534 5172 12568
rect 5206 12534 5244 12568
rect 5278 12534 5284 12568
rect 5166 12495 5284 12534
rect 5166 12461 5172 12495
rect 5206 12461 5244 12495
rect 5278 12461 5284 12495
rect 5166 12422 5284 12461
rect 5166 11892 5172 12422
rect 5278 11892 5284 12422
rect 5166 11826 5172 11840
rect 5278 11826 5284 11840
rect 5166 11760 5172 11774
rect 5278 11760 5284 11774
rect 5166 11694 5172 11708
rect 5278 11694 5284 11708
rect 5166 11628 5172 11642
rect 5278 11628 5284 11642
rect 5166 11562 5172 11576
rect 5278 11562 5284 11576
rect 5166 11495 5172 11510
rect 5278 11495 5284 11510
rect 5166 11428 5172 11443
rect 5278 11428 5284 11443
rect 5218 11376 5232 11380
rect 5166 10714 5284 11376
rect 5166 10680 5172 10714
rect 5206 10680 5244 10714
rect 5278 10680 5284 10714
rect 5166 10641 5284 10680
rect 5166 10607 5172 10641
rect 5206 10607 5244 10641
rect 5278 10607 5284 10641
rect 5166 10568 5284 10607
rect 5166 10534 5172 10568
rect 5206 10534 5244 10568
rect 5278 10534 5284 10568
rect 5166 10495 5284 10534
rect 5166 10461 5172 10495
rect 5206 10461 5244 10495
rect 5278 10461 5284 10495
rect 5166 10422 5284 10461
rect 5166 9896 5172 10422
rect 5278 9896 5284 10422
rect 5166 9830 5172 9844
rect 5278 9830 5284 9844
rect 5166 9764 5172 9778
rect 5278 9764 5284 9778
rect 5166 9698 5172 9712
rect 5278 9698 5284 9712
rect 5166 9632 5172 9646
rect 5278 9632 5284 9646
rect 5166 9566 5172 9580
rect 5278 9566 5284 9580
rect 5166 9499 5172 9514
rect 5278 9499 5284 9514
rect 5166 9432 5172 9447
rect 5278 9432 5284 9447
rect 5166 8714 5284 9380
rect 5166 8680 5172 8714
rect 5206 8680 5244 8714
rect 5278 8680 5284 8714
rect 5166 8641 5284 8680
rect 5166 8607 5172 8641
rect 5206 8607 5244 8641
rect 5278 8607 5284 8641
rect 5166 8568 5284 8607
rect 5166 8534 5172 8568
rect 5206 8534 5244 8568
rect 5278 8534 5284 8568
rect 5166 8495 5284 8534
rect 5166 8461 5172 8495
rect 5206 8461 5244 8495
rect 5278 8461 5284 8495
rect 5166 8422 5284 8461
rect 5166 7892 5172 8422
rect 5278 7892 5284 8422
rect 5166 7826 5172 7840
rect 5278 7826 5284 7840
rect 5166 7760 5172 7774
rect 5278 7760 5284 7774
rect 5166 7694 5172 7708
rect 5278 7694 5284 7708
rect 5166 7628 5172 7642
rect 5278 7628 5284 7642
rect 5166 7562 5172 7576
rect 5278 7562 5284 7576
rect 5166 7495 5172 7510
rect 5278 7495 5284 7510
rect 5166 7428 5172 7443
rect 5278 7428 5284 7443
rect 5218 7376 5232 7380
rect 5166 6714 5284 7376
rect 5166 6680 5172 6714
rect 5206 6680 5244 6714
rect 5278 6680 5284 6714
rect 5166 6641 5284 6680
rect 5166 6607 5172 6641
rect 5206 6607 5244 6641
rect 5278 6607 5284 6641
rect 5166 6568 5284 6607
rect 5166 6534 5172 6568
rect 5206 6534 5244 6568
rect 5278 6534 5284 6568
rect 5166 6495 5284 6534
rect 5166 6461 5172 6495
rect 5206 6461 5244 6495
rect 5278 6461 5284 6495
rect 5166 6422 5284 6461
rect 5166 5896 5172 6422
rect 5278 5896 5284 6422
rect 5166 5830 5172 5844
rect 5278 5830 5284 5844
rect 5166 5764 5172 5778
rect 5278 5764 5284 5778
rect 5166 5698 5172 5712
rect 5278 5698 5284 5712
rect 5166 5632 5172 5646
rect 5278 5632 5284 5646
rect 5166 5566 5172 5580
rect 5278 5566 5284 5580
rect 5166 5499 5172 5514
rect 5278 5499 5284 5514
rect 5166 5432 5172 5447
rect 5278 5432 5284 5447
rect 5166 5368 5284 5380
rect 5495 14338 5509 14390
rect 5997 14720 6115 14726
rect 6049 14668 6063 14720
rect 5997 14654 6115 14668
rect 6049 14602 6063 14654
rect 5997 14588 6115 14602
rect 6049 14536 6063 14588
rect 5997 14522 6115 14536
rect 6049 14470 6063 14522
rect 5997 14456 6115 14470
rect 6049 14404 6063 14456
rect 5997 14390 6115 14404
rect 5443 14323 5449 14338
rect 5483 14323 5521 14338
rect 5555 14323 5561 14338
rect 5495 14271 5509 14323
rect 5443 14267 5561 14271
rect 5443 14256 5449 14267
rect 5483 14256 5521 14267
rect 5555 14256 5561 14267
rect 5495 14204 5509 14256
rect 5443 14189 5561 14204
rect 5443 14155 5449 14189
rect 5483 14155 5521 14189
rect 5555 14155 5561 14189
rect 5443 14111 5561 14155
rect 5443 14077 5449 14111
rect 5483 14077 5521 14111
rect 5555 14077 5561 14111
rect 5443 14033 5561 14077
rect 5443 13999 5449 14033
rect 5483 13999 5521 14033
rect 5555 13999 5561 14033
rect 5443 13955 5561 13999
rect 5443 13921 5449 13955
rect 5483 13921 5521 13955
rect 5555 13921 5561 13955
rect 5443 13877 5561 13921
rect 5443 13843 5449 13877
rect 5483 13843 5521 13877
rect 5555 13843 5561 13877
rect 5443 13799 5561 13843
rect 5443 13765 5449 13799
rect 5483 13765 5521 13799
rect 5555 13765 5561 13799
rect 5443 13722 5561 13765
rect 5443 13688 5449 13722
rect 5483 13688 5521 13722
rect 5555 13688 5561 13722
rect 5443 13645 5561 13688
rect 5443 13611 5449 13645
rect 5483 13611 5521 13645
rect 5555 13611 5561 13645
rect 5443 13568 5561 13611
rect 5443 13534 5449 13568
rect 5483 13534 5521 13568
rect 5555 13534 5561 13568
rect 5443 13491 5561 13534
rect 5443 13457 5449 13491
rect 5483 13457 5521 13491
rect 5555 13457 5561 13491
rect 5443 13414 5561 13457
rect 5443 13380 5449 13414
rect 5483 13380 5521 13414
rect 5555 13380 5561 13414
rect 5443 12720 5561 13380
rect 5495 12668 5509 12720
rect 5443 12654 5561 12668
rect 5495 12602 5509 12654
rect 5443 12588 5561 12602
rect 5495 12536 5509 12588
rect 5443 12534 5449 12536
rect 5483 12534 5521 12536
rect 5555 12534 5561 12536
rect 5443 12522 5561 12534
rect 5495 12470 5509 12522
rect 5443 12461 5449 12470
rect 5483 12461 5521 12470
rect 5555 12461 5561 12470
rect 5443 12456 5561 12461
rect 5495 12422 5509 12456
rect 5443 12390 5449 12404
rect 5555 12390 5561 12404
rect 5443 12323 5449 12338
rect 5555 12323 5561 12338
rect 5443 12256 5449 12271
rect 5555 12256 5561 12271
rect 5443 11380 5449 12204
rect 5555 11380 5561 12204
rect 5443 10724 5561 11380
rect 5495 10672 5509 10724
rect 5443 10658 5561 10672
rect 5495 10606 5509 10658
rect 5443 10592 5561 10606
rect 5495 10540 5509 10592
rect 5443 10534 5449 10540
rect 5483 10534 5521 10540
rect 5555 10534 5561 10540
rect 5443 10526 5561 10534
rect 5495 10474 5509 10526
rect 5443 10461 5449 10474
rect 5483 10461 5521 10474
rect 5555 10461 5561 10474
rect 5443 10460 5561 10461
rect 5495 10422 5509 10460
rect 5443 10394 5449 10408
rect 5555 10394 5561 10408
rect 5443 10327 5449 10342
rect 5555 10327 5561 10342
rect 5443 10260 5449 10275
rect 5555 10260 5561 10275
rect 5443 9380 5449 10208
rect 5555 9380 5561 10208
rect 5443 8720 5561 9380
rect 5495 8668 5509 8720
rect 5443 8654 5561 8668
rect 5495 8602 5509 8654
rect 5443 8588 5561 8602
rect 5495 8536 5509 8588
rect 5443 8534 5449 8536
rect 5483 8534 5521 8536
rect 5555 8534 5561 8536
rect 5443 8522 5561 8534
rect 5495 8470 5509 8522
rect 5443 8461 5449 8470
rect 5483 8461 5521 8470
rect 5555 8461 5561 8470
rect 5443 8456 5561 8461
rect 5495 8422 5509 8456
rect 5443 8390 5449 8404
rect 5555 8390 5561 8404
rect 5443 8323 5449 8338
rect 5555 8323 5561 8338
rect 5443 8256 5449 8271
rect 5555 8256 5561 8271
rect 5443 7380 5449 8204
rect 5555 7380 5561 8204
rect 5443 6724 5561 7380
rect 5495 6672 5509 6724
rect 5443 6658 5561 6672
rect 5495 6606 5509 6658
rect 5443 6592 5561 6606
rect 5495 6540 5509 6592
rect 5443 6534 5449 6540
rect 5483 6534 5521 6540
rect 5555 6534 5561 6540
rect 5443 6526 5561 6534
rect 5495 6474 5509 6526
rect 5443 6461 5449 6474
rect 5483 6461 5521 6474
rect 5555 6461 5561 6474
rect 5443 6460 5561 6461
rect 5495 6422 5509 6460
rect 5443 6394 5449 6408
rect 5555 6394 5561 6408
rect 5443 6327 5449 6342
rect 5555 6327 5561 6342
rect 5443 6260 5449 6275
rect 5555 6260 5561 6275
rect 5443 5380 5449 6208
rect 5555 5380 5561 6208
tri 5007 5265 5013 5271 sw
tri 5437 5265 5443 5271 se
rect 5443 5265 5561 5380
rect 5720 14345 5838 14357
rect 5720 14311 5726 14345
rect 5760 14311 5798 14345
rect 5832 14311 5838 14345
rect 5720 14267 5838 14311
rect 5720 14233 5726 14267
rect 5760 14233 5798 14267
rect 5832 14233 5838 14267
rect 5720 14189 5838 14233
rect 5720 14155 5726 14189
rect 5760 14155 5798 14189
rect 5832 14155 5838 14189
rect 5720 14111 5838 14155
rect 5720 14077 5726 14111
rect 5760 14077 5798 14111
rect 5832 14077 5838 14111
rect 5720 14033 5838 14077
rect 5720 13999 5726 14033
rect 5760 13999 5798 14033
rect 5832 13999 5838 14033
rect 5720 13955 5838 13999
rect 5720 13921 5726 13955
rect 5760 13921 5798 13955
rect 5832 13921 5838 13955
rect 5720 13892 5838 13921
rect 5772 13840 5786 13892
rect 5720 13826 5838 13840
rect 5772 13774 5786 13826
rect 5720 13765 5726 13774
rect 5760 13765 5798 13774
rect 5832 13765 5838 13774
rect 5720 13760 5838 13765
rect 5772 13708 5786 13760
rect 5720 13694 5726 13708
rect 5760 13694 5798 13708
rect 5832 13694 5838 13708
rect 5772 13642 5786 13694
rect 5720 13628 5726 13642
rect 5760 13628 5798 13642
rect 5832 13628 5838 13642
rect 5772 13576 5786 13628
rect 5720 13568 5838 13576
rect 5720 13562 5726 13568
rect 5760 13562 5798 13568
rect 5832 13562 5838 13568
rect 5772 13510 5786 13562
rect 5720 13495 5838 13510
rect 5772 13443 5786 13495
rect 5720 13428 5838 13443
rect 5772 13376 5786 13428
rect 5720 12714 5838 13376
rect 5720 12680 5726 12714
rect 5760 12680 5798 12714
rect 5832 12680 5838 12714
rect 5720 12641 5838 12680
rect 5720 12607 5726 12641
rect 5760 12607 5798 12641
rect 5832 12607 5838 12641
rect 5720 12568 5838 12607
rect 5720 12534 5726 12568
rect 5760 12534 5798 12568
rect 5832 12534 5838 12568
rect 5720 12495 5838 12534
rect 5720 12461 5726 12495
rect 5760 12461 5798 12495
rect 5832 12461 5838 12495
rect 5720 12422 5838 12461
rect 5720 11892 5726 12422
rect 5832 11892 5838 12422
rect 5720 11826 5726 11840
rect 5832 11826 5838 11840
rect 5720 11760 5726 11774
rect 5832 11760 5838 11774
rect 5720 11694 5726 11708
rect 5832 11694 5838 11708
rect 5720 11628 5726 11642
rect 5832 11628 5838 11642
rect 5720 11562 5726 11576
rect 5832 11562 5838 11576
rect 5720 11495 5726 11510
rect 5832 11495 5838 11510
rect 5720 11428 5726 11443
rect 5832 11428 5838 11443
rect 5772 11376 5786 11380
rect 5720 10714 5838 11376
rect 5720 10680 5726 10714
rect 5760 10680 5798 10714
rect 5832 10680 5838 10714
rect 5720 10641 5838 10680
rect 5720 10607 5726 10641
rect 5760 10607 5798 10641
rect 5832 10607 5838 10641
rect 5720 10568 5838 10607
rect 5720 10534 5726 10568
rect 5760 10534 5798 10568
rect 5832 10534 5838 10568
rect 5720 10495 5838 10534
rect 5720 10461 5726 10495
rect 5760 10461 5798 10495
rect 5832 10461 5838 10495
rect 5720 10422 5838 10461
rect 5720 9896 5726 10422
rect 5832 9896 5838 10422
rect 5720 9830 5726 9844
rect 5832 9830 5838 9844
rect 5720 9764 5726 9778
rect 5832 9764 5838 9778
rect 5720 9698 5726 9712
rect 5832 9698 5838 9712
rect 5720 9632 5726 9646
rect 5832 9632 5838 9646
rect 5720 9566 5726 9580
rect 5832 9566 5838 9580
rect 5720 9499 5726 9514
rect 5832 9499 5838 9514
rect 5720 9432 5726 9447
rect 5832 9432 5838 9447
rect 5720 8714 5838 9380
rect 5720 8680 5726 8714
rect 5760 8680 5798 8714
rect 5832 8680 5838 8714
rect 5720 8641 5838 8680
rect 5720 8607 5726 8641
rect 5760 8607 5798 8641
rect 5832 8607 5838 8641
rect 5720 8568 5838 8607
rect 5720 8534 5726 8568
rect 5760 8534 5798 8568
rect 5832 8534 5838 8568
rect 5720 8495 5838 8534
rect 5720 8461 5726 8495
rect 5760 8461 5798 8495
rect 5832 8461 5838 8495
rect 5720 8422 5838 8461
rect 5720 7892 5726 8422
rect 5832 7892 5838 8422
rect 5720 7826 5726 7840
rect 5832 7826 5838 7840
rect 5720 7760 5726 7774
rect 5832 7760 5838 7774
rect 5720 7694 5726 7708
rect 5832 7694 5838 7708
rect 5720 7628 5726 7642
rect 5832 7628 5838 7642
rect 5720 7562 5726 7576
rect 5832 7562 5838 7576
rect 5720 7495 5726 7510
rect 5832 7495 5838 7510
rect 5720 7428 5726 7443
rect 5832 7428 5838 7443
rect 5772 7376 5786 7380
rect 5720 6714 5838 7376
rect 5720 6680 5726 6714
rect 5760 6680 5798 6714
rect 5832 6680 5838 6714
rect 5720 6641 5838 6680
rect 5720 6607 5726 6641
rect 5760 6607 5798 6641
rect 5832 6607 5838 6641
rect 5720 6568 5838 6607
rect 5720 6534 5726 6568
rect 5760 6534 5798 6568
rect 5832 6534 5838 6568
rect 5720 6495 5838 6534
rect 5720 6461 5726 6495
rect 5760 6461 5798 6495
rect 5832 6461 5838 6495
rect 5720 6422 5838 6461
rect 5720 5896 5726 6422
rect 5832 5896 5838 6422
rect 5720 5830 5726 5844
rect 5832 5830 5838 5844
rect 5720 5764 5726 5778
rect 5832 5764 5838 5778
rect 5720 5698 5726 5712
rect 5832 5698 5838 5712
rect 5720 5632 5726 5646
rect 5832 5632 5838 5646
rect 5720 5566 5726 5580
rect 5832 5566 5838 5580
rect 5720 5499 5726 5514
rect 5832 5499 5838 5514
rect 5720 5432 5726 5447
rect 5832 5432 5838 5447
rect 5720 5368 5838 5380
rect 6049 14338 6063 14390
rect 6551 14720 6669 14726
rect 6603 14668 6617 14720
rect 6551 14654 6669 14668
rect 6603 14602 6617 14654
rect 6551 14588 6669 14602
rect 6603 14536 6617 14588
rect 6551 14522 6669 14536
rect 6603 14470 6617 14522
rect 6551 14456 6669 14470
rect 6603 14404 6617 14456
rect 6551 14390 6669 14404
rect 5997 14323 6003 14338
rect 6037 14323 6075 14338
rect 6109 14323 6115 14338
rect 6049 14271 6063 14323
rect 5997 14267 6115 14271
rect 5997 14256 6003 14267
rect 6037 14256 6075 14267
rect 6109 14256 6115 14267
rect 6049 14204 6063 14256
rect 5997 14189 6115 14204
rect 5997 14155 6003 14189
rect 6037 14155 6075 14189
rect 6109 14155 6115 14189
rect 5997 14111 6115 14155
rect 5997 14077 6003 14111
rect 6037 14077 6075 14111
rect 6109 14077 6115 14111
rect 5997 14033 6115 14077
rect 5997 13999 6003 14033
rect 6037 13999 6075 14033
rect 6109 13999 6115 14033
rect 5997 13955 6115 13999
rect 5997 13921 6003 13955
rect 6037 13921 6075 13955
rect 6109 13921 6115 13955
rect 5997 13877 6115 13921
rect 5997 13843 6003 13877
rect 6037 13843 6075 13877
rect 6109 13843 6115 13877
rect 5997 13799 6115 13843
rect 5997 13765 6003 13799
rect 6037 13765 6075 13799
rect 6109 13765 6115 13799
rect 5997 13722 6115 13765
rect 5997 13688 6003 13722
rect 6037 13688 6075 13722
rect 6109 13688 6115 13722
rect 5997 13645 6115 13688
rect 5997 13611 6003 13645
rect 6037 13611 6075 13645
rect 6109 13611 6115 13645
rect 5997 13568 6115 13611
rect 5997 13534 6003 13568
rect 6037 13534 6075 13568
rect 6109 13534 6115 13568
rect 5997 13491 6115 13534
rect 5997 13457 6003 13491
rect 6037 13457 6075 13491
rect 6109 13457 6115 13491
rect 5997 13414 6115 13457
rect 5997 13380 6003 13414
rect 6037 13380 6075 13414
rect 6109 13380 6115 13414
rect 5997 12720 6115 13380
rect 6049 12668 6063 12720
rect 5997 12654 6115 12668
rect 6049 12602 6063 12654
rect 5997 12588 6115 12602
rect 6049 12536 6063 12588
rect 5997 12534 6003 12536
rect 6037 12534 6075 12536
rect 6109 12534 6115 12536
rect 5997 12522 6115 12534
rect 6049 12470 6063 12522
rect 5997 12461 6003 12470
rect 6037 12461 6075 12470
rect 6109 12461 6115 12470
rect 5997 12456 6115 12461
rect 6049 12422 6063 12456
rect 5997 12390 6003 12404
rect 6109 12390 6115 12404
rect 5997 12323 6003 12338
rect 6109 12323 6115 12338
rect 5997 12256 6003 12271
rect 6109 12256 6115 12271
rect 5997 11380 6003 12204
rect 6109 11380 6115 12204
rect 5997 10724 6115 11380
rect 6049 10672 6063 10724
rect 5997 10658 6115 10672
rect 6049 10606 6063 10658
rect 5997 10592 6115 10606
rect 6049 10540 6063 10592
rect 5997 10534 6003 10540
rect 6037 10534 6075 10540
rect 6109 10534 6115 10540
rect 5997 10526 6115 10534
rect 6049 10474 6063 10526
rect 5997 10461 6003 10474
rect 6037 10461 6075 10474
rect 6109 10461 6115 10474
rect 5997 10460 6115 10461
rect 6049 10422 6063 10460
rect 5997 10394 6003 10408
rect 6109 10394 6115 10408
rect 5997 10327 6003 10342
rect 6109 10327 6115 10342
rect 5997 10260 6003 10275
rect 6109 10260 6115 10275
rect 5997 9380 6003 10208
rect 6109 9380 6115 10208
rect 5997 8720 6115 9380
rect 6049 8668 6063 8720
rect 5997 8654 6115 8668
rect 6049 8602 6063 8654
rect 5997 8588 6115 8602
rect 6049 8536 6063 8588
rect 5997 8534 6003 8536
rect 6037 8534 6075 8536
rect 6109 8534 6115 8536
rect 5997 8522 6115 8534
rect 6049 8470 6063 8522
rect 5997 8461 6003 8470
rect 6037 8461 6075 8470
rect 6109 8461 6115 8470
rect 5997 8456 6115 8461
rect 6049 8422 6063 8456
rect 5997 8390 6003 8404
rect 6109 8390 6115 8404
rect 5997 8323 6003 8338
rect 6109 8323 6115 8338
rect 5997 8256 6003 8271
rect 6109 8256 6115 8271
rect 5997 7380 6003 8204
rect 6109 7380 6115 8204
rect 5997 6724 6115 7380
rect 6049 6672 6063 6724
rect 5997 6658 6115 6672
rect 6049 6606 6063 6658
rect 5997 6592 6115 6606
rect 6049 6540 6063 6592
rect 5997 6534 6003 6540
rect 6037 6534 6075 6540
rect 6109 6534 6115 6540
rect 5997 6526 6115 6534
rect 6049 6474 6063 6526
rect 5997 6461 6003 6474
rect 6037 6461 6075 6474
rect 6109 6461 6115 6474
rect 5997 6460 6115 6461
rect 6049 6422 6063 6460
rect 5997 6394 6003 6408
rect 6109 6394 6115 6408
rect 5997 6327 6003 6342
rect 6109 6327 6115 6342
rect 5997 6260 6003 6275
rect 6109 6260 6115 6275
rect 5997 5380 6003 6208
rect 6109 5380 6115 6208
tri 5561 5265 5567 5271 sw
tri 5991 5265 5997 5271 se
rect 5997 5265 6115 5380
rect 6274 14345 6392 14357
rect 6274 14311 6280 14345
rect 6314 14311 6352 14345
rect 6386 14311 6392 14345
rect 6274 14267 6392 14311
rect 6274 14233 6280 14267
rect 6314 14233 6352 14267
rect 6386 14233 6392 14267
rect 6274 14189 6392 14233
rect 6274 14155 6280 14189
rect 6314 14155 6352 14189
rect 6386 14155 6392 14189
rect 6274 14111 6392 14155
rect 6274 14077 6280 14111
rect 6314 14077 6352 14111
rect 6386 14077 6392 14111
rect 6274 14033 6392 14077
rect 6274 13999 6280 14033
rect 6314 13999 6352 14033
rect 6386 13999 6392 14033
rect 6274 13955 6392 13999
rect 6274 13921 6280 13955
rect 6314 13921 6352 13955
rect 6386 13921 6392 13955
rect 6274 13892 6392 13921
rect 6326 13840 6340 13892
rect 6274 13826 6392 13840
rect 6326 13774 6340 13826
rect 6274 13765 6280 13774
rect 6314 13765 6352 13774
rect 6386 13765 6392 13774
rect 6274 13760 6392 13765
rect 6326 13708 6340 13760
rect 6274 13694 6280 13708
rect 6314 13694 6352 13708
rect 6386 13694 6392 13708
rect 6326 13642 6340 13694
rect 6274 13628 6280 13642
rect 6314 13628 6352 13642
rect 6386 13628 6392 13642
rect 6326 13576 6340 13628
rect 6274 13568 6392 13576
rect 6274 13562 6280 13568
rect 6314 13562 6352 13568
rect 6386 13562 6392 13568
rect 6326 13510 6340 13562
rect 6274 13495 6392 13510
rect 6326 13443 6340 13495
rect 6274 13428 6392 13443
rect 6326 13376 6340 13428
rect 6274 12714 6392 13376
rect 6274 12680 6280 12714
rect 6314 12680 6352 12714
rect 6386 12680 6392 12714
rect 6274 12641 6392 12680
rect 6274 12607 6280 12641
rect 6314 12607 6352 12641
rect 6386 12607 6392 12641
rect 6274 12568 6392 12607
rect 6274 12534 6280 12568
rect 6314 12534 6352 12568
rect 6386 12534 6392 12568
rect 6274 12495 6392 12534
rect 6274 12461 6280 12495
rect 6314 12461 6352 12495
rect 6386 12461 6392 12495
rect 6274 12422 6392 12461
rect 6274 11892 6280 12422
rect 6386 11892 6392 12422
rect 6274 11826 6280 11840
rect 6386 11826 6392 11840
rect 6274 11760 6280 11774
rect 6386 11760 6392 11774
rect 6274 11694 6280 11708
rect 6386 11694 6392 11708
rect 6274 11628 6280 11642
rect 6386 11628 6392 11642
rect 6274 11562 6280 11576
rect 6386 11562 6392 11576
rect 6274 11495 6280 11510
rect 6386 11495 6392 11510
rect 6274 11428 6280 11443
rect 6386 11428 6392 11443
rect 6326 11376 6340 11380
rect 6274 10714 6392 11376
rect 6274 10680 6280 10714
rect 6314 10680 6352 10714
rect 6386 10680 6392 10714
rect 6274 10641 6392 10680
rect 6274 10607 6280 10641
rect 6314 10607 6352 10641
rect 6386 10607 6392 10641
rect 6274 10568 6392 10607
rect 6274 10534 6280 10568
rect 6314 10534 6352 10568
rect 6386 10534 6392 10568
rect 6274 10495 6392 10534
rect 6274 10461 6280 10495
rect 6314 10461 6352 10495
rect 6386 10461 6392 10495
rect 6274 10422 6392 10461
rect 6274 9896 6280 10422
rect 6386 9896 6392 10422
rect 6274 9830 6280 9844
rect 6386 9830 6392 9844
rect 6274 9764 6280 9778
rect 6386 9764 6392 9778
rect 6274 9698 6280 9712
rect 6386 9698 6392 9712
rect 6274 9632 6280 9646
rect 6386 9632 6392 9646
rect 6274 9566 6280 9580
rect 6386 9566 6392 9580
rect 6274 9499 6280 9514
rect 6386 9499 6392 9514
rect 6274 9432 6280 9447
rect 6386 9432 6392 9447
rect 6274 8714 6392 9380
rect 6274 8680 6280 8714
rect 6314 8680 6352 8714
rect 6386 8680 6392 8714
rect 6274 8641 6392 8680
rect 6274 8607 6280 8641
rect 6314 8607 6352 8641
rect 6386 8607 6392 8641
rect 6274 8568 6392 8607
rect 6274 8534 6280 8568
rect 6314 8534 6352 8568
rect 6386 8534 6392 8568
rect 6274 8495 6392 8534
rect 6274 8461 6280 8495
rect 6314 8461 6352 8495
rect 6386 8461 6392 8495
rect 6274 8422 6392 8461
rect 6274 7892 6280 8422
rect 6386 7892 6392 8422
rect 6274 7826 6280 7840
rect 6386 7826 6392 7840
rect 6274 7760 6280 7774
rect 6386 7760 6392 7774
rect 6274 7694 6280 7708
rect 6386 7694 6392 7708
rect 6274 7628 6280 7642
rect 6386 7628 6392 7642
rect 6274 7562 6280 7576
rect 6386 7562 6392 7576
rect 6274 7495 6280 7510
rect 6386 7495 6392 7510
rect 6274 7428 6280 7443
rect 6386 7428 6392 7443
rect 6326 7376 6340 7380
rect 6274 6714 6392 7376
rect 6274 6680 6280 6714
rect 6314 6680 6352 6714
rect 6386 6680 6392 6714
rect 6274 6641 6392 6680
rect 6274 6607 6280 6641
rect 6314 6607 6352 6641
rect 6386 6607 6392 6641
rect 6274 6568 6392 6607
rect 6274 6534 6280 6568
rect 6314 6534 6352 6568
rect 6386 6534 6392 6568
rect 6274 6495 6392 6534
rect 6274 6461 6280 6495
rect 6314 6461 6352 6495
rect 6386 6461 6392 6495
rect 6274 6422 6392 6461
rect 6274 5896 6280 6422
rect 6386 5896 6392 6422
rect 6274 5830 6280 5844
rect 6386 5830 6392 5844
rect 6274 5764 6280 5778
rect 6386 5764 6392 5778
rect 6274 5698 6280 5712
rect 6386 5698 6392 5712
rect 6274 5632 6280 5646
rect 6386 5632 6392 5646
rect 6274 5566 6280 5580
rect 6386 5566 6392 5580
rect 6274 5499 6280 5514
rect 6386 5499 6392 5514
rect 6274 5432 6280 5447
rect 6386 5432 6392 5447
rect 6274 5368 6392 5380
rect 6603 14338 6617 14390
rect 7105 14720 7223 14726
rect 7157 14668 7171 14720
rect 7105 14654 7223 14668
rect 7157 14602 7171 14654
rect 7105 14588 7223 14602
rect 7157 14536 7171 14588
rect 7105 14522 7223 14536
rect 7157 14470 7171 14522
rect 7105 14456 7223 14470
rect 7157 14404 7171 14456
rect 7105 14390 7223 14404
rect 6551 14323 6557 14338
rect 6591 14323 6629 14338
rect 6663 14323 6669 14338
rect 6603 14271 6617 14323
rect 6551 14267 6669 14271
rect 6551 14256 6557 14267
rect 6591 14256 6629 14267
rect 6663 14256 6669 14267
rect 6603 14204 6617 14256
rect 6551 14189 6669 14204
rect 6551 14155 6557 14189
rect 6591 14155 6629 14189
rect 6663 14155 6669 14189
rect 6551 14111 6669 14155
rect 6551 14077 6557 14111
rect 6591 14077 6629 14111
rect 6663 14077 6669 14111
rect 6551 14033 6669 14077
rect 6551 13999 6557 14033
rect 6591 13999 6629 14033
rect 6663 13999 6669 14033
rect 6551 13955 6669 13999
rect 6551 13921 6557 13955
rect 6591 13921 6629 13955
rect 6663 13921 6669 13955
rect 6551 13877 6669 13921
rect 6551 13843 6557 13877
rect 6591 13843 6629 13877
rect 6663 13843 6669 13877
rect 6551 13799 6669 13843
rect 6551 13765 6557 13799
rect 6591 13765 6629 13799
rect 6663 13765 6669 13799
rect 6551 13722 6669 13765
rect 6551 13688 6557 13722
rect 6591 13688 6629 13722
rect 6663 13688 6669 13722
rect 6551 13645 6669 13688
rect 6551 13611 6557 13645
rect 6591 13611 6629 13645
rect 6663 13611 6669 13645
rect 6551 13568 6669 13611
rect 6551 13534 6557 13568
rect 6591 13534 6629 13568
rect 6663 13534 6669 13568
rect 6551 13491 6669 13534
rect 6551 13457 6557 13491
rect 6591 13457 6629 13491
rect 6663 13457 6669 13491
rect 6551 13414 6669 13457
rect 6551 13380 6557 13414
rect 6591 13380 6629 13414
rect 6663 13380 6669 13414
rect 6551 12720 6669 13380
rect 6603 12668 6617 12720
rect 6551 12654 6669 12668
rect 6603 12602 6617 12654
rect 6551 12588 6669 12602
rect 6603 12536 6617 12588
rect 6551 12534 6557 12536
rect 6591 12534 6629 12536
rect 6663 12534 6669 12536
rect 6551 12522 6669 12534
rect 6603 12470 6617 12522
rect 6551 12461 6557 12470
rect 6591 12461 6629 12470
rect 6663 12461 6669 12470
rect 6551 12456 6669 12461
rect 6603 12422 6617 12456
rect 6551 12390 6557 12404
rect 6663 12390 6669 12404
rect 6551 12323 6557 12338
rect 6663 12323 6669 12338
rect 6551 12256 6557 12271
rect 6663 12256 6669 12271
rect 6551 11380 6557 12204
rect 6663 11380 6669 12204
rect 6551 10724 6669 11380
rect 6603 10672 6617 10724
rect 6551 10658 6669 10672
rect 6603 10606 6617 10658
rect 6551 10592 6669 10606
rect 6603 10540 6617 10592
rect 6551 10534 6557 10540
rect 6591 10534 6629 10540
rect 6663 10534 6669 10540
rect 6551 10526 6669 10534
rect 6603 10474 6617 10526
rect 6551 10461 6557 10474
rect 6591 10461 6629 10474
rect 6663 10461 6669 10474
rect 6551 10460 6669 10461
rect 6603 10422 6617 10460
rect 6551 10394 6557 10408
rect 6663 10394 6669 10408
rect 6551 10327 6557 10342
rect 6663 10327 6669 10342
rect 6551 10260 6557 10275
rect 6663 10260 6669 10275
rect 6551 9380 6557 10208
rect 6663 9380 6669 10208
rect 6551 8720 6669 9380
rect 6603 8668 6617 8720
rect 6551 8654 6669 8668
rect 6603 8602 6617 8654
rect 6551 8588 6669 8602
rect 6603 8536 6617 8588
rect 6551 8534 6557 8536
rect 6591 8534 6629 8536
rect 6663 8534 6669 8536
rect 6551 8522 6669 8534
rect 6603 8470 6617 8522
rect 6551 8461 6557 8470
rect 6591 8461 6629 8470
rect 6663 8461 6669 8470
rect 6551 8456 6669 8461
rect 6603 8422 6617 8456
rect 6551 8390 6557 8404
rect 6663 8390 6669 8404
rect 6551 8323 6557 8338
rect 6663 8323 6669 8338
rect 6551 8256 6557 8271
rect 6663 8256 6669 8271
rect 6551 7380 6557 8204
rect 6663 7380 6669 8204
rect 6551 6724 6669 7380
rect 6603 6672 6617 6724
rect 6551 6658 6669 6672
rect 6603 6606 6617 6658
rect 6551 6592 6669 6606
rect 6603 6540 6617 6592
rect 6551 6534 6557 6540
rect 6591 6534 6629 6540
rect 6663 6534 6669 6540
rect 6551 6526 6669 6534
rect 6603 6474 6617 6526
rect 6551 6461 6557 6474
rect 6591 6461 6629 6474
rect 6663 6461 6669 6474
rect 6551 6460 6669 6461
rect 6603 6422 6617 6460
rect 6551 6394 6557 6408
rect 6663 6394 6669 6408
rect 6551 6327 6557 6342
rect 6663 6327 6669 6342
rect 6551 6260 6557 6275
rect 6663 6260 6669 6275
rect 6551 5380 6557 6208
rect 6663 5380 6669 6208
tri 6115 5265 6121 5271 sw
tri 6545 5265 6551 5271 se
rect 6551 5265 6669 5380
rect 6828 14345 6946 14357
rect 6828 14311 6834 14345
rect 6868 14311 6906 14345
rect 6940 14311 6946 14345
rect 6828 14267 6946 14311
rect 6828 14233 6834 14267
rect 6868 14233 6906 14267
rect 6940 14233 6946 14267
rect 6828 14189 6946 14233
rect 6828 14155 6834 14189
rect 6868 14155 6906 14189
rect 6940 14155 6946 14189
rect 6828 14111 6946 14155
rect 6828 14077 6834 14111
rect 6868 14077 6906 14111
rect 6940 14077 6946 14111
rect 6828 14033 6946 14077
rect 6828 13999 6834 14033
rect 6868 13999 6906 14033
rect 6940 13999 6946 14033
rect 6828 13955 6946 13999
rect 6828 13921 6834 13955
rect 6868 13921 6906 13955
rect 6940 13921 6946 13955
rect 6828 13892 6946 13921
rect 6880 13840 6894 13892
rect 6828 13826 6946 13840
rect 6880 13774 6894 13826
rect 6828 13765 6834 13774
rect 6868 13765 6906 13774
rect 6940 13765 6946 13774
rect 6828 13760 6946 13765
rect 6880 13708 6894 13760
rect 6828 13694 6834 13708
rect 6868 13694 6906 13708
rect 6940 13694 6946 13708
rect 6880 13642 6894 13694
rect 6828 13628 6834 13642
rect 6868 13628 6906 13642
rect 6940 13628 6946 13642
rect 6880 13576 6894 13628
rect 6828 13568 6946 13576
rect 6828 13562 6834 13568
rect 6868 13562 6906 13568
rect 6940 13562 6946 13568
rect 6880 13510 6894 13562
rect 6828 13495 6946 13510
rect 6880 13443 6894 13495
rect 6828 13428 6946 13443
rect 6880 13376 6894 13428
rect 6828 12714 6946 13376
rect 6828 12680 6834 12714
rect 6868 12680 6906 12714
rect 6940 12680 6946 12714
rect 6828 12641 6946 12680
rect 6828 12607 6834 12641
rect 6868 12607 6906 12641
rect 6940 12607 6946 12641
rect 6828 12568 6946 12607
rect 6828 12534 6834 12568
rect 6868 12534 6906 12568
rect 6940 12534 6946 12568
rect 6828 12495 6946 12534
rect 6828 12461 6834 12495
rect 6868 12461 6906 12495
rect 6940 12461 6946 12495
rect 6828 12422 6946 12461
rect 6828 11892 6834 12422
rect 6940 11892 6946 12422
rect 6828 11826 6834 11840
rect 6940 11826 6946 11840
rect 6828 11760 6834 11774
rect 6940 11760 6946 11774
rect 6828 11694 6834 11708
rect 6940 11694 6946 11708
rect 6828 11628 6834 11642
rect 6940 11628 6946 11642
rect 6828 11562 6834 11576
rect 6940 11562 6946 11576
rect 6828 11495 6834 11510
rect 6940 11495 6946 11510
rect 6828 11428 6834 11443
rect 6940 11428 6946 11443
rect 6880 11376 6894 11380
rect 6828 10714 6946 11376
rect 6828 10680 6834 10714
rect 6868 10680 6906 10714
rect 6940 10680 6946 10714
rect 6828 10641 6946 10680
rect 6828 10607 6834 10641
rect 6868 10607 6906 10641
rect 6940 10607 6946 10641
rect 6828 10568 6946 10607
rect 6828 10534 6834 10568
rect 6868 10534 6906 10568
rect 6940 10534 6946 10568
rect 6828 10495 6946 10534
rect 6828 10461 6834 10495
rect 6868 10461 6906 10495
rect 6940 10461 6946 10495
rect 6828 10422 6946 10461
rect 6828 9896 6834 10422
rect 6940 9896 6946 10422
rect 6828 9830 6834 9844
rect 6940 9830 6946 9844
rect 6828 9764 6834 9778
rect 6940 9764 6946 9778
rect 6828 9698 6834 9712
rect 6940 9698 6946 9712
rect 6828 9632 6834 9646
rect 6940 9632 6946 9646
rect 6828 9566 6834 9580
rect 6940 9566 6946 9580
rect 6828 9499 6834 9514
rect 6940 9499 6946 9514
rect 6828 9432 6834 9447
rect 6940 9432 6946 9447
rect 6828 8714 6946 9380
rect 6828 8680 6834 8714
rect 6868 8680 6906 8714
rect 6940 8680 6946 8714
rect 6828 8641 6946 8680
rect 6828 8607 6834 8641
rect 6868 8607 6906 8641
rect 6940 8607 6946 8641
rect 6828 8568 6946 8607
rect 6828 8534 6834 8568
rect 6868 8534 6906 8568
rect 6940 8534 6946 8568
rect 6828 8495 6946 8534
rect 6828 8461 6834 8495
rect 6868 8461 6906 8495
rect 6940 8461 6946 8495
rect 6828 8422 6946 8461
rect 6828 7892 6834 8422
rect 6940 7892 6946 8422
rect 6828 7826 6834 7840
rect 6940 7826 6946 7840
rect 6828 7760 6834 7774
rect 6940 7760 6946 7774
rect 6828 7694 6834 7708
rect 6940 7694 6946 7708
rect 6828 7628 6834 7642
rect 6940 7628 6946 7642
rect 6828 7562 6834 7576
rect 6940 7562 6946 7576
rect 6828 7495 6834 7510
rect 6940 7495 6946 7510
rect 6828 7428 6834 7443
rect 6940 7428 6946 7443
rect 6880 7376 6894 7380
rect 6828 6714 6946 7376
rect 6828 6680 6834 6714
rect 6868 6680 6906 6714
rect 6940 6680 6946 6714
rect 6828 6641 6946 6680
rect 6828 6607 6834 6641
rect 6868 6607 6906 6641
rect 6940 6607 6946 6641
rect 6828 6568 6946 6607
rect 6828 6534 6834 6568
rect 6868 6534 6906 6568
rect 6940 6534 6946 6568
rect 6828 6495 6946 6534
rect 6828 6461 6834 6495
rect 6868 6461 6906 6495
rect 6940 6461 6946 6495
rect 6828 6422 6946 6461
rect 6828 5896 6834 6422
rect 6940 5896 6946 6422
rect 6828 5830 6834 5844
rect 6940 5830 6946 5844
rect 6828 5764 6834 5778
rect 6940 5764 6946 5778
rect 6828 5698 6834 5712
rect 6940 5698 6946 5712
rect 6828 5632 6834 5646
rect 6940 5632 6946 5646
rect 6828 5566 6834 5580
rect 6940 5566 6946 5580
rect 6828 5499 6834 5514
rect 6940 5499 6946 5514
rect 6828 5432 6834 5447
rect 6940 5432 6946 5447
rect 6828 5368 6946 5380
rect 7157 14338 7171 14390
rect 7659 14720 7777 14726
rect 7711 14668 7725 14720
rect 7659 14654 7777 14668
rect 7711 14602 7725 14654
rect 7659 14588 7777 14602
rect 7711 14536 7725 14588
rect 7659 14522 7777 14536
rect 7711 14470 7725 14522
rect 7659 14456 7777 14470
rect 7711 14404 7725 14456
rect 7659 14390 7777 14404
rect 7105 14323 7111 14338
rect 7145 14323 7183 14338
rect 7217 14323 7223 14338
rect 7157 14271 7171 14323
rect 7105 14267 7223 14271
rect 7105 14256 7111 14267
rect 7145 14256 7183 14267
rect 7217 14256 7223 14267
rect 7157 14204 7171 14256
rect 7105 14189 7223 14204
rect 7105 14155 7111 14189
rect 7145 14155 7183 14189
rect 7217 14155 7223 14189
rect 7105 14111 7223 14155
rect 7105 14077 7111 14111
rect 7145 14077 7183 14111
rect 7217 14077 7223 14111
rect 7105 14033 7223 14077
rect 7105 13999 7111 14033
rect 7145 13999 7183 14033
rect 7217 13999 7223 14033
rect 7105 13955 7223 13999
rect 7105 13921 7111 13955
rect 7145 13921 7183 13955
rect 7217 13921 7223 13955
rect 7105 13877 7223 13921
rect 7105 13843 7111 13877
rect 7145 13843 7183 13877
rect 7217 13843 7223 13877
rect 7105 13799 7223 13843
rect 7105 13765 7111 13799
rect 7145 13765 7183 13799
rect 7217 13765 7223 13799
rect 7105 13722 7223 13765
rect 7105 13688 7111 13722
rect 7145 13688 7183 13722
rect 7217 13688 7223 13722
rect 7105 13645 7223 13688
rect 7105 13611 7111 13645
rect 7145 13611 7183 13645
rect 7217 13611 7223 13645
rect 7105 13568 7223 13611
rect 7105 13534 7111 13568
rect 7145 13534 7183 13568
rect 7217 13534 7223 13568
rect 7105 13491 7223 13534
rect 7105 13457 7111 13491
rect 7145 13457 7183 13491
rect 7217 13457 7223 13491
rect 7105 13414 7223 13457
rect 7105 13380 7111 13414
rect 7145 13380 7183 13414
rect 7217 13380 7223 13414
rect 7105 12720 7223 13380
rect 7157 12668 7171 12720
rect 7105 12654 7223 12668
rect 7157 12602 7171 12654
rect 7105 12588 7223 12602
rect 7157 12536 7171 12588
rect 7105 12534 7111 12536
rect 7145 12534 7183 12536
rect 7217 12534 7223 12536
rect 7105 12522 7223 12534
rect 7157 12470 7171 12522
rect 7105 12461 7111 12470
rect 7145 12461 7183 12470
rect 7217 12461 7223 12470
rect 7105 12456 7223 12461
rect 7157 12422 7171 12456
rect 7105 12390 7111 12404
rect 7217 12390 7223 12404
rect 7105 12323 7111 12338
rect 7217 12323 7223 12338
rect 7105 12256 7111 12271
rect 7217 12256 7223 12271
rect 7105 11380 7111 12204
rect 7217 11380 7223 12204
rect 7105 10724 7223 11380
rect 7157 10672 7171 10724
rect 7105 10658 7223 10672
rect 7157 10606 7171 10658
rect 7105 10592 7223 10606
rect 7157 10540 7171 10592
rect 7105 10534 7111 10540
rect 7145 10534 7183 10540
rect 7217 10534 7223 10540
rect 7105 10526 7223 10534
rect 7157 10474 7171 10526
rect 7105 10461 7111 10474
rect 7145 10461 7183 10474
rect 7217 10461 7223 10474
rect 7105 10460 7223 10461
rect 7157 10422 7171 10460
rect 7105 10394 7111 10408
rect 7217 10394 7223 10408
rect 7105 10327 7111 10342
rect 7217 10327 7223 10342
rect 7105 10260 7111 10275
rect 7217 10260 7223 10275
rect 7105 9380 7111 10208
rect 7217 9380 7223 10208
rect 7105 8720 7223 9380
rect 7157 8668 7171 8720
rect 7105 8654 7223 8668
rect 7157 8602 7171 8654
rect 7105 8588 7223 8602
rect 7157 8536 7171 8588
rect 7105 8534 7111 8536
rect 7145 8534 7183 8536
rect 7217 8534 7223 8536
rect 7105 8522 7223 8534
rect 7157 8470 7171 8522
rect 7105 8461 7111 8470
rect 7145 8461 7183 8470
rect 7217 8461 7223 8470
rect 7105 8456 7223 8461
rect 7157 8422 7171 8456
rect 7105 8390 7111 8404
rect 7217 8390 7223 8404
rect 7105 8323 7111 8338
rect 7217 8323 7223 8338
rect 7105 8256 7111 8271
rect 7217 8256 7223 8271
rect 7105 7380 7111 8204
rect 7217 7380 7223 8204
rect 7105 6724 7223 7380
rect 7157 6672 7171 6724
rect 7105 6658 7223 6672
rect 7157 6606 7171 6658
rect 7105 6592 7223 6606
rect 7157 6540 7171 6592
rect 7105 6534 7111 6540
rect 7145 6534 7183 6540
rect 7217 6534 7223 6540
rect 7105 6526 7223 6534
rect 7157 6474 7171 6526
rect 7105 6461 7111 6474
rect 7145 6461 7183 6474
rect 7217 6461 7223 6474
rect 7105 6460 7223 6461
rect 7157 6422 7171 6460
rect 7105 6394 7111 6408
rect 7217 6394 7223 6408
rect 7105 6327 7111 6342
rect 7217 6327 7223 6342
rect 7105 6260 7111 6275
rect 7217 6260 7223 6275
rect 7105 5380 7111 6208
rect 7217 5380 7223 6208
tri 6669 5265 6675 5271 sw
tri 7099 5265 7105 5271 se
rect 7105 5265 7223 5380
rect 7382 14345 7500 14357
rect 7382 14311 7388 14345
rect 7422 14311 7460 14345
rect 7494 14311 7500 14345
rect 7382 14267 7500 14311
rect 7382 14233 7388 14267
rect 7422 14233 7460 14267
rect 7494 14233 7500 14267
rect 7382 14189 7500 14233
rect 7382 14155 7388 14189
rect 7422 14155 7460 14189
rect 7494 14155 7500 14189
rect 7382 14111 7500 14155
rect 7382 14077 7388 14111
rect 7422 14077 7460 14111
rect 7494 14077 7500 14111
rect 7382 14033 7500 14077
rect 7382 13999 7388 14033
rect 7422 13999 7460 14033
rect 7494 13999 7500 14033
rect 7382 13955 7500 13999
rect 7382 13921 7388 13955
rect 7422 13921 7460 13955
rect 7494 13921 7500 13955
rect 7382 13892 7500 13921
rect 7434 13840 7448 13892
rect 7382 13826 7500 13840
rect 7434 13774 7448 13826
rect 7382 13765 7388 13774
rect 7422 13765 7460 13774
rect 7494 13765 7500 13774
rect 7382 13760 7500 13765
rect 7434 13708 7448 13760
rect 7382 13694 7388 13708
rect 7422 13694 7460 13708
rect 7494 13694 7500 13708
rect 7434 13642 7448 13694
rect 7382 13628 7388 13642
rect 7422 13628 7460 13642
rect 7494 13628 7500 13642
rect 7434 13576 7448 13628
rect 7382 13568 7500 13576
rect 7382 13562 7388 13568
rect 7422 13562 7460 13568
rect 7494 13562 7500 13568
rect 7434 13510 7448 13562
rect 7382 13495 7500 13510
rect 7434 13443 7448 13495
rect 7382 13428 7500 13443
rect 7434 13376 7448 13428
rect 7382 12714 7500 13376
rect 7382 12680 7388 12714
rect 7422 12680 7460 12714
rect 7494 12680 7500 12714
rect 7382 12641 7500 12680
rect 7382 12607 7388 12641
rect 7422 12607 7460 12641
rect 7494 12607 7500 12641
rect 7382 12568 7500 12607
rect 7382 12534 7388 12568
rect 7422 12534 7460 12568
rect 7494 12534 7500 12568
rect 7382 12495 7500 12534
rect 7382 12461 7388 12495
rect 7422 12461 7460 12495
rect 7494 12461 7500 12495
rect 7382 12422 7500 12461
rect 7382 11892 7388 12422
rect 7494 11892 7500 12422
rect 7382 11826 7388 11840
rect 7494 11826 7500 11840
rect 7382 11760 7388 11774
rect 7494 11760 7500 11774
rect 7382 11694 7388 11708
rect 7494 11694 7500 11708
rect 7382 11628 7388 11642
rect 7494 11628 7500 11642
rect 7382 11562 7388 11576
rect 7494 11562 7500 11576
rect 7382 11495 7388 11510
rect 7494 11495 7500 11510
rect 7382 11428 7388 11443
rect 7494 11428 7500 11443
rect 7434 11376 7448 11380
rect 7382 10714 7500 11376
rect 7382 10680 7388 10714
rect 7422 10680 7460 10714
rect 7494 10680 7500 10714
rect 7382 10641 7500 10680
rect 7382 10607 7388 10641
rect 7422 10607 7460 10641
rect 7494 10607 7500 10641
rect 7382 10568 7500 10607
rect 7382 10534 7388 10568
rect 7422 10534 7460 10568
rect 7494 10534 7500 10568
rect 7382 10495 7500 10534
rect 7382 10461 7388 10495
rect 7422 10461 7460 10495
rect 7494 10461 7500 10495
rect 7382 10422 7500 10461
rect 7382 9896 7388 10422
rect 7494 9896 7500 10422
rect 7382 9830 7388 9844
rect 7494 9830 7500 9844
rect 7382 9764 7388 9778
rect 7494 9764 7500 9778
rect 7382 9698 7388 9712
rect 7494 9698 7500 9712
rect 7382 9632 7388 9646
rect 7494 9632 7500 9646
rect 7382 9566 7388 9580
rect 7494 9566 7500 9580
rect 7382 9499 7388 9514
rect 7494 9499 7500 9514
rect 7382 9432 7388 9447
rect 7494 9432 7500 9447
rect 7382 8714 7500 9380
rect 7382 8680 7388 8714
rect 7422 8680 7460 8714
rect 7494 8680 7500 8714
rect 7382 8641 7500 8680
rect 7382 8607 7388 8641
rect 7422 8607 7460 8641
rect 7494 8607 7500 8641
rect 7382 8568 7500 8607
rect 7382 8534 7388 8568
rect 7422 8534 7460 8568
rect 7494 8534 7500 8568
rect 7382 8495 7500 8534
rect 7382 8461 7388 8495
rect 7422 8461 7460 8495
rect 7494 8461 7500 8495
rect 7382 8422 7500 8461
rect 7382 7892 7388 8422
rect 7494 7892 7500 8422
rect 7382 7826 7388 7840
rect 7494 7826 7500 7840
rect 7382 7760 7388 7774
rect 7494 7760 7500 7774
rect 7382 7694 7388 7708
rect 7494 7694 7500 7708
rect 7382 7628 7388 7642
rect 7494 7628 7500 7642
rect 7382 7562 7388 7576
rect 7494 7562 7500 7576
rect 7382 7495 7388 7510
rect 7494 7495 7500 7510
rect 7382 7428 7388 7443
rect 7494 7428 7500 7443
rect 7434 7376 7448 7380
rect 7382 6714 7500 7376
rect 7382 6680 7388 6714
rect 7422 6680 7460 6714
rect 7494 6680 7500 6714
rect 7382 6641 7500 6680
rect 7382 6607 7388 6641
rect 7422 6607 7460 6641
rect 7494 6607 7500 6641
rect 7382 6568 7500 6607
rect 7382 6534 7388 6568
rect 7422 6534 7460 6568
rect 7494 6534 7500 6568
rect 7382 6495 7500 6534
rect 7382 6461 7388 6495
rect 7422 6461 7460 6495
rect 7494 6461 7500 6495
rect 7382 6422 7500 6461
rect 7382 5896 7388 6422
rect 7494 5896 7500 6422
rect 7382 5830 7388 5844
rect 7494 5830 7500 5844
rect 7382 5764 7388 5778
rect 7494 5764 7500 5778
rect 7382 5698 7388 5712
rect 7494 5698 7500 5712
rect 7382 5632 7388 5646
rect 7494 5632 7500 5646
rect 7382 5566 7388 5580
rect 7494 5566 7500 5580
rect 7382 5499 7388 5514
rect 7494 5499 7500 5514
rect 7382 5432 7388 5447
rect 7494 5432 7500 5447
rect 7382 5368 7500 5380
rect 7711 14338 7725 14390
rect 8213 14720 8331 14726
rect 8265 14668 8279 14720
rect 8213 14654 8331 14668
rect 8265 14602 8279 14654
rect 8213 14588 8331 14602
rect 8265 14536 8279 14588
rect 8213 14522 8331 14536
rect 8265 14470 8279 14522
rect 8213 14456 8331 14470
rect 8265 14404 8279 14456
rect 8213 14390 8331 14404
rect 7659 14323 7665 14338
rect 7699 14323 7737 14338
rect 7771 14323 7777 14338
rect 7711 14271 7725 14323
rect 7659 14267 7777 14271
rect 7659 14256 7665 14267
rect 7699 14256 7737 14267
rect 7771 14256 7777 14267
rect 7711 14204 7725 14256
rect 7659 14189 7777 14204
rect 7659 14155 7665 14189
rect 7699 14155 7737 14189
rect 7771 14155 7777 14189
rect 7659 14111 7777 14155
rect 7659 14077 7665 14111
rect 7699 14077 7737 14111
rect 7771 14077 7777 14111
rect 7659 14033 7777 14077
rect 7659 13999 7665 14033
rect 7699 13999 7737 14033
rect 7771 13999 7777 14033
rect 7659 13955 7777 13999
rect 7659 13921 7665 13955
rect 7699 13921 7737 13955
rect 7771 13921 7777 13955
rect 7659 13877 7777 13921
rect 7659 13843 7665 13877
rect 7699 13843 7737 13877
rect 7771 13843 7777 13877
rect 7659 13799 7777 13843
rect 7659 13765 7665 13799
rect 7699 13765 7737 13799
rect 7771 13765 7777 13799
rect 7659 13722 7777 13765
rect 7659 13688 7665 13722
rect 7699 13688 7737 13722
rect 7771 13688 7777 13722
rect 7659 13645 7777 13688
rect 7659 13611 7665 13645
rect 7699 13611 7737 13645
rect 7771 13611 7777 13645
rect 7659 13568 7777 13611
rect 7659 13534 7665 13568
rect 7699 13534 7737 13568
rect 7771 13534 7777 13568
rect 7659 13491 7777 13534
rect 7659 13457 7665 13491
rect 7699 13457 7737 13491
rect 7771 13457 7777 13491
rect 7659 13414 7777 13457
rect 7659 13380 7665 13414
rect 7699 13380 7737 13414
rect 7771 13380 7777 13414
rect 7659 12720 7777 13380
rect 7711 12668 7725 12720
rect 7659 12654 7777 12668
rect 7711 12602 7725 12654
rect 7659 12588 7777 12602
rect 7711 12536 7725 12588
rect 7659 12534 7665 12536
rect 7699 12534 7737 12536
rect 7771 12534 7777 12536
rect 7659 12522 7777 12534
rect 7711 12470 7725 12522
rect 7659 12461 7665 12470
rect 7699 12461 7737 12470
rect 7771 12461 7777 12470
rect 7659 12456 7777 12461
rect 7711 12422 7725 12456
rect 7659 12390 7665 12404
rect 7771 12390 7777 12404
rect 7659 12323 7665 12338
rect 7771 12323 7777 12338
rect 7659 12256 7665 12271
rect 7771 12256 7777 12271
rect 7659 11380 7665 12204
rect 7771 11380 7777 12204
rect 7659 10724 7777 11380
rect 7711 10672 7725 10724
rect 7659 10658 7777 10672
rect 7711 10606 7725 10658
rect 7659 10592 7777 10606
rect 7711 10540 7725 10592
rect 7659 10534 7665 10540
rect 7699 10534 7737 10540
rect 7771 10534 7777 10540
rect 7659 10526 7777 10534
rect 7711 10474 7725 10526
rect 7659 10461 7665 10474
rect 7699 10461 7737 10474
rect 7771 10461 7777 10474
rect 7659 10460 7777 10461
rect 7711 10422 7725 10460
rect 7659 10394 7665 10408
rect 7771 10394 7777 10408
rect 7659 10327 7665 10342
rect 7771 10327 7777 10342
rect 7659 10260 7665 10275
rect 7771 10260 7777 10275
rect 7659 9380 7665 10208
rect 7771 9380 7777 10208
rect 7659 8720 7777 9380
rect 7711 8668 7725 8720
rect 7659 8654 7777 8668
rect 7711 8602 7725 8654
rect 7659 8588 7777 8602
rect 7711 8536 7725 8588
rect 7659 8534 7665 8536
rect 7699 8534 7737 8536
rect 7771 8534 7777 8536
rect 7659 8522 7777 8534
rect 7711 8470 7725 8522
rect 7659 8461 7665 8470
rect 7699 8461 7737 8470
rect 7771 8461 7777 8470
rect 7659 8456 7777 8461
rect 7711 8422 7725 8456
rect 7659 8390 7665 8404
rect 7771 8390 7777 8404
rect 7659 8323 7665 8338
rect 7771 8323 7777 8338
rect 7659 8256 7665 8271
rect 7771 8256 7777 8271
rect 7659 7380 7665 8204
rect 7771 7380 7777 8204
rect 7659 6724 7777 7380
rect 7711 6672 7725 6724
rect 7659 6658 7777 6672
rect 7711 6606 7725 6658
rect 7659 6592 7777 6606
rect 7711 6540 7725 6592
rect 7659 6534 7665 6540
rect 7699 6534 7737 6540
rect 7771 6534 7777 6540
rect 7659 6526 7777 6534
rect 7711 6474 7725 6526
rect 7659 6461 7665 6474
rect 7699 6461 7737 6474
rect 7771 6461 7777 6474
rect 7659 6460 7777 6461
rect 7711 6422 7725 6460
rect 7659 6394 7665 6408
rect 7771 6394 7777 6408
rect 7659 6327 7665 6342
rect 7771 6327 7777 6342
rect 7659 6260 7665 6275
rect 7771 6260 7777 6275
rect 7659 5380 7665 6208
rect 7771 5380 7777 6208
tri 7223 5265 7229 5271 sw
tri 7653 5265 7659 5271 se
rect 7659 5265 7777 5380
rect 7936 14345 8054 14357
rect 7936 14311 7942 14345
rect 7976 14311 8014 14345
rect 8048 14311 8054 14345
rect 7936 14267 8054 14311
rect 7936 14233 7942 14267
rect 7976 14233 8014 14267
rect 8048 14233 8054 14267
rect 7936 14189 8054 14233
rect 7936 14155 7942 14189
rect 7976 14155 8014 14189
rect 8048 14155 8054 14189
rect 7936 14111 8054 14155
rect 7936 14077 7942 14111
rect 7976 14077 8014 14111
rect 8048 14077 8054 14111
rect 7936 14033 8054 14077
rect 7936 13999 7942 14033
rect 7976 13999 8014 14033
rect 8048 13999 8054 14033
rect 7936 13955 8054 13999
rect 7936 13921 7942 13955
rect 7976 13921 8014 13955
rect 8048 13921 8054 13955
rect 7936 13892 8054 13921
rect 7988 13840 8002 13892
rect 7936 13826 8054 13840
rect 7988 13774 8002 13826
rect 7936 13765 7942 13774
rect 7976 13765 8014 13774
rect 8048 13765 8054 13774
rect 7936 13760 8054 13765
rect 7988 13708 8002 13760
rect 7936 13694 7942 13708
rect 7976 13694 8014 13708
rect 8048 13694 8054 13708
rect 7988 13642 8002 13694
rect 7936 13628 7942 13642
rect 7976 13628 8014 13642
rect 8048 13628 8054 13642
rect 7988 13576 8002 13628
rect 7936 13568 8054 13576
rect 7936 13562 7942 13568
rect 7976 13562 8014 13568
rect 8048 13562 8054 13568
rect 7988 13510 8002 13562
rect 7936 13495 8054 13510
rect 7988 13443 8002 13495
rect 7936 13428 8054 13443
rect 7988 13376 8002 13428
rect 7936 12714 8054 13376
rect 7936 12680 7942 12714
rect 7976 12680 8014 12714
rect 8048 12680 8054 12714
rect 7936 12641 8054 12680
rect 7936 12607 7942 12641
rect 7976 12607 8014 12641
rect 8048 12607 8054 12641
rect 7936 12568 8054 12607
rect 7936 12534 7942 12568
rect 7976 12534 8014 12568
rect 8048 12534 8054 12568
rect 7936 12495 8054 12534
rect 7936 12461 7942 12495
rect 7976 12461 8014 12495
rect 8048 12461 8054 12495
rect 7936 12422 8054 12461
rect 7936 11892 7942 12422
rect 8048 11892 8054 12422
rect 7936 11826 7942 11840
rect 8048 11826 8054 11840
rect 7936 11760 7942 11774
rect 8048 11760 8054 11774
rect 7936 11694 7942 11708
rect 8048 11694 8054 11708
rect 7936 11628 7942 11642
rect 8048 11628 8054 11642
rect 7936 11562 7942 11576
rect 8048 11562 8054 11576
rect 7936 11495 7942 11510
rect 8048 11495 8054 11510
rect 7936 11428 7942 11443
rect 8048 11428 8054 11443
rect 7988 11376 8002 11380
rect 7936 10714 8054 11376
rect 7936 10680 7942 10714
rect 7976 10680 8014 10714
rect 8048 10680 8054 10714
rect 7936 10641 8054 10680
rect 7936 10607 7942 10641
rect 7976 10607 8014 10641
rect 8048 10607 8054 10641
rect 7936 10568 8054 10607
rect 7936 10534 7942 10568
rect 7976 10534 8014 10568
rect 8048 10534 8054 10568
rect 7936 10495 8054 10534
rect 7936 10461 7942 10495
rect 7976 10461 8014 10495
rect 8048 10461 8054 10495
rect 7936 10422 8054 10461
rect 7936 9896 7942 10422
rect 8048 9896 8054 10422
rect 7936 9830 7942 9844
rect 8048 9830 8054 9844
rect 7936 9764 7942 9778
rect 8048 9764 8054 9778
rect 7936 9698 7942 9712
rect 8048 9698 8054 9712
rect 7936 9632 7942 9646
rect 8048 9632 8054 9646
rect 7936 9566 7942 9580
rect 8048 9566 8054 9580
rect 7936 9499 7942 9514
rect 8048 9499 8054 9514
rect 7936 9432 7942 9447
rect 8048 9432 8054 9447
rect 7936 8714 8054 9380
rect 7936 8680 7942 8714
rect 7976 8680 8014 8714
rect 8048 8680 8054 8714
rect 7936 8641 8054 8680
rect 7936 8607 7942 8641
rect 7976 8607 8014 8641
rect 8048 8607 8054 8641
rect 7936 8568 8054 8607
rect 7936 8534 7942 8568
rect 7976 8534 8014 8568
rect 8048 8534 8054 8568
rect 7936 8495 8054 8534
rect 7936 8461 7942 8495
rect 7976 8461 8014 8495
rect 8048 8461 8054 8495
rect 7936 8422 8054 8461
rect 7936 7892 7942 8422
rect 8048 7892 8054 8422
rect 7936 7826 7942 7840
rect 8048 7826 8054 7840
rect 7936 7760 7942 7774
rect 8048 7760 8054 7774
rect 7936 7694 7942 7708
rect 8048 7694 8054 7708
rect 7936 7628 7942 7642
rect 8048 7628 8054 7642
rect 7936 7562 7942 7576
rect 8048 7562 8054 7576
rect 7936 7495 7942 7510
rect 8048 7495 8054 7510
rect 7936 7428 7942 7443
rect 8048 7428 8054 7443
rect 7988 7376 8002 7380
rect 7936 6714 8054 7376
rect 7936 6680 7942 6714
rect 7976 6680 8014 6714
rect 8048 6680 8054 6714
rect 7936 6641 8054 6680
rect 7936 6607 7942 6641
rect 7976 6607 8014 6641
rect 8048 6607 8054 6641
rect 7936 6568 8054 6607
rect 7936 6534 7942 6568
rect 7976 6534 8014 6568
rect 8048 6534 8054 6568
rect 7936 6495 8054 6534
rect 7936 6461 7942 6495
rect 7976 6461 8014 6495
rect 8048 6461 8054 6495
rect 7936 6422 8054 6461
rect 7936 5896 7942 6422
rect 8048 5896 8054 6422
rect 7936 5830 7942 5844
rect 8048 5830 8054 5844
rect 7936 5764 7942 5778
rect 8048 5764 8054 5778
rect 7936 5698 7942 5712
rect 8048 5698 8054 5712
rect 7936 5632 7942 5646
rect 8048 5632 8054 5646
rect 7936 5566 7942 5580
rect 8048 5566 8054 5580
rect 7936 5499 7942 5514
rect 8048 5499 8054 5514
rect 7936 5432 7942 5447
rect 8048 5432 8054 5447
rect 7936 5368 8054 5380
rect 8265 14338 8279 14390
rect 8767 14720 8885 14726
rect 8819 14668 8833 14720
rect 8767 14654 8885 14668
rect 8819 14602 8833 14654
rect 8767 14588 8885 14602
rect 8819 14536 8833 14588
rect 8767 14522 8885 14536
rect 8819 14470 8833 14522
rect 8767 14456 8885 14470
rect 8819 14404 8833 14456
rect 8767 14390 8885 14404
rect 8213 14323 8219 14338
rect 8253 14323 8291 14338
rect 8325 14323 8331 14338
rect 8265 14271 8279 14323
rect 8213 14267 8331 14271
rect 8213 14256 8219 14267
rect 8253 14256 8291 14267
rect 8325 14256 8331 14267
rect 8265 14204 8279 14256
rect 8213 14189 8331 14204
rect 8213 14155 8219 14189
rect 8253 14155 8291 14189
rect 8325 14155 8331 14189
rect 8213 14111 8331 14155
rect 8213 14077 8219 14111
rect 8253 14077 8291 14111
rect 8325 14077 8331 14111
rect 8213 14033 8331 14077
rect 8213 13999 8219 14033
rect 8253 13999 8291 14033
rect 8325 13999 8331 14033
rect 8213 13955 8331 13999
rect 8213 13921 8219 13955
rect 8253 13921 8291 13955
rect 8325 13921 8331 13955
rect 8213 13877 8331 13921
rect 8213 13843 8219 13877
rect 8253 13843 8291 13877
rect 8325 13843 8331 13877
rect 8213 13799 8331 13843
rect 8213 13765 8219 13799
rect 8253 13765 8291 13799
rect 8325 13765 8331 13799
rect 8213 13722 8331 13765
rect 8213 13688 8219 13722
rect 8253 13688 8291 13722
rect 8325 13688 8331 13722
rect 8213 13645 8331 13688
rect 8213 13611 8219 13645
rect 8253 13611 8291 13645
rect 8325 13611 8331 13645
rect 8213 13568 8331 13611
rect 8213 13534 8219 13568
rect 8253 13534 8291 13568
rect 8325 13534 8331 13568
rect 8213 13491 8331 13534
rect 8213 13457 8219 13491
rect 8253 13457 8291 13491
rect 8325 13457 8331 13491
rect 8213 13414 8331 13457
rect 8213 13380 8219 13414
rect 8253 13380 8291 13414
rect 8325 13380 8331 13414
rect 8213 12720 8331 13380
rect 8265 12668 8279 12720
rect 8213 12654 8331 12668
rect 8265 12602 8279 12654
rect 8213 12588 8331 12602
rect 8265 12536 8279 12588
rect 8213 12534 8219 12536
rect 8253 12534 8291 12536
rect 8325 12534 8331 12536
rect 8213 12522 8331 12534
rect 8265 12470 8279 12522
rect 8213 12461 8219 12470
rect 8253 12461 8291 12470
rect 8325 12461 8331 12470
rect 8213 12456 8331 12461
rect 8265 12422 8279 12456
rect 8213 12390 8219 12404
rect 8325 12390 8331 12404
rect 8213 12323 8219 12338
rect 8325 12323 8331 12338
rect 8213 12256 8219 12271
rect 8325 12256 8331 12271
rect 8213 11380 8219 12204
rect 8325 11380 8331 12204
rect 8213 10724 8331 11380
rect 8265 10672 8279 10724
rect 8213 10658 8331 10672
rect 8265 10606 8279 10658
rect 8213 10592 8331 10606
rect 8265 10540 8279 10592
rect 8213 10534 8219 10540
rect 8253 10534 8291 10540
rect 8325 10534 8331 10540
rect 8213 10526 8331 10534
rect 8265 10474 8279 10526
rect 8213 10461 8219 10474
rect 8253 10461 8291 10474
rect 8325 10461 8331 10474
rect 8213 10460 8331 10461
rect 8265 10422 8279 10460
rect 8213 10394 8219 10408
rect 8325 10394 8331 10408
rect 8213 10327 8219 10342
rect 8325 10327 8331 10342
rect 8213 10260 8219 10275
rect 8325 10260 8331 10275
rect 8213 9380 8219 10208
rect 8325 9380 8331 10208
rect 8213 8720 8331 9380
rect 8265 8668 8279 8720
rect 8213 8654 8331 8668
rect 8265 8602 8279 8654
rect 8213 8588 8331 8602
rect 8265 8536 8279 8588
rect 8213 8534 8219 8536
rect 8253 8534 8291 8536
rect 8325 8534 8331 8536
rect 8213 8522 8331 8534
rect 8265 8470 8279 8522
rect 8213 8461 8219 8470
rect 8253 8461 8291 8470
rect 8325 8461 8331 8470
rect 8213 8456 8331 8461
rect 8265 8422 8279 8456
rect 8213 8390 8219 8404
rect 8325 8390 8331 8404
rect 8213 8323 8219 8338
rect 8325 8323 8331 8338
rect 8213 8256 8219 8271
rect 8325 8256 8331 8271
rect 8213 7380 8219 8204
rect 8325 7380 8331 8204
rect 8213 6724 8331 7380
rect 8265 6672 8279 6724
rect 8213 6658 8331 6672
rect 8265 6606 8279 6658
rect 8213 6592 8331 6606
rect 8265 6540 8279 6592
rect 8213 6534 8219 6540
rect 8253 6534 8291 6540
rect 8325 6534 8331 6540
rect 8213 6526 8331 6534
rect 8265 6474 8279 6526
rect 8213 6461 8219 6474
rect 8253 6461 8291 6474
rect 8325 6461 8331 6474
rect 8213 6460 8331 6461
rect 8265 6422 8279 6460
rect 8213 6394 8219 6408
rect 8325 6394 8331 6408
rect 8213 6327 8219 6342
rect 8325 6327 8331 6342
rect 8213 6260 8219 6275
rect 8325 6260 8331 6275
rect 8213 5380 8219 6208
rect 8325 5380 8331 6208
tri 7777 5265 7783 5271 sw
tri 8207 5265 8213 5271 se
rect 8213 5265 8331 5380
rect 8490 14345 8608 14357
rect 8490 14311 8496 14345
rect 8530 14311 8568 14345
rect 8602 14311 8608 14345
rect 8490 14267 8608 14311
rect 8490 14233 8496 14267
rect 8530 14233 8568 14267
rect 8602 14233 8608 14267
rect 8490 14189 8608 14233
rect 8490 14155 8496 14189
rect 8530 14155 8568 14189
rect 8602 14155 8608 14189
rect 8490 14111 8608 14155
rect 8490 14077 8496 14111
rect 8530 14077 8568 14111
rect 8602 14077 8608 14111
rect 8490 14033 8608 14077
rect 8490 13999 8496 14033
rect 8530 13999 8568 14033
rect 8602 13999 8608 14033
rect 8490 13955 8608 13999
rect 8490 13921 8496 13955
rect 8530 13921 8568 13955
rect 8602 13921 8608 13955
rect 8490 13892 8608 13921
rect 8542 13840 8556 13892
rect 8490 13826 8608 13840
rect 8542 13774 8556 13826
rect 8490 13765 8496 13774
rect 8530 13765 8568 13774
rect 8602 13765 8608 13774
rect 8490 13760 8608 13765
rect 8542 13708 8556 13760
rect 8490 13694 8496 13708
rect 8530 13694 8568 13708
rect 8602 13694 8608 13708
rect 8542 13642 8556 13694
rect 8490 13628 8496 13642
rect 8530 13628 8568 13642
rect 8602 13628 8608 13642
rect 8542 13576 8556 13628
rect 8490 13568 8608 13576
rect 8490 13562 8496 13568
rect 8530 13562 8568 13568
rect 8602 13562 8608 13568
rect 8542 13510 8556 13562
rect 8490 13495 8608 13510
rect 8542 13443 8556 13495
rect 8490 13428 8608 13443
rect 8542 13376 8556 13428
rect 8490 12714 8608 13376
rect 8490 12680 8496 12714
rect 8530 12680 8568 12714
rect 8602 12680 8608 12714
rect 8490 12641 8608 12680
rect 8490 12607 8496 12641
rect 8530 12607 8568 12641
rect 8602 12607 8608 12641
rect 8490 12568 8608 12607
rect 8490 12534 8496 12568
rect 8530 12534 8568 12568
rect 8602 12534 8608 12568
rect 8490 12495 8608 12534
rect 8490 12461 8496 12495
rect 8530 12461 8568 12495
rect 8602 12461 8608 12495
rect 8490 12422 8608 12461
rect 8490 11892 8496 12422
rect 8602 11892 8608 12422
rect 8490 11826 8496 11840
rect 8602 11826 8608 11840
rect 8490 11760 8496 11774
rect 8602 11760 8608 11774
rect 8490 11694 8496 11708
rect 8602 11694 8608 11708
rect 8490 11628 8496 11642
rect 8602 11628 8608 11642
rect 8490 11562 8496 11576
rect 8602 11562 8608 11576
rect 8490 11495 8496 11510
rect 8602 11495 8608 11510
rect 8490 11428 8496 11443
rect 8602 11428 8608 11443
rect 8542 11376 8556 11380
rect 8490 10714 8608 11376
rect 8490 10680 8496 10714
rect 8530 10680 8568 10714
rect 8602 10680 8608 10714
rect 8490 10641 8608 10680
rect 8490 10607 8496 10641
rect 8530 10607 8568 10641
rect 8602 10607 8608 10641
rect 8490 10568 8608 10607
rect 8490 10534 8496 10568
rect 8530 10534 8568 10568
rect 8602 10534 8608 10568
rect 8490 10495 8608 10534
rect 8490 10461 8496 10495
rect 8530 10461 8568 10495
rect 8602 10461 8608 10495
rect 8490 10422 8608 10461
rect 8490 9896 8496 10422
rect 8602 9896 8608 10422
rect 8490 9830 8496 9844
rect 8602 9830 8608 9844
rect 8490 9764 8496 9778
rect 8602 9764 8608 9778
rect 8490 9698 8496 9712
rect 8602 9698 8608 9712
rect 8490 9632 8496 9646
rect 8602 9632 8608 9646
rect 8490 9566 8496 9580
rect 8602 9566 8608 9580
rect 8490 9499 8496 9514
rect 8602 9499 8608 9514
rect 8490 9432 8496 9447
rect 8602 9432 8608 9447
rect 8490 8714 8608 9380
rect 8490 8680 8496 8714
rect 8530 8680 8568 8714
rect 8602 8680 8608 8714
rect 8490 8641 8608 8680
rect 8490 8607 8496 8641
rect 8530 8607 8568 8641
rect 8602 8607 8608 8641
rect 8490 8568 8608 8607
rect 8490 8534 8496 8568
rect 8530 8534 8568 8568
rect 8602 8534 8608 8568
rect 8490 8495 8608 8534
rect 8490 8461 8496 8495
rect 8530 8461 8568 8495
rect 8602 8461 8608 8495
rect 8490 8422 8608 8461
rect 8490 7892 8496 8422
rect 8602 7892 8608 8422
rect 8490 7826 8496 7840
rect 8602 7826 8608 7840
rect 8490 7760 8496 7774
rect 8602 7760 8608 7774
rect 8490 7694 8496 7708
rect 8602 7694 8608 7708
rect 8490 7628 8496 7642
rect 8602 7628 8608 7642
rect 8490 7562 8496 7576
rect 8602 7562 8608 7576
rect 8490 7495 8496 7510
rect 8602 7495 8608 7510
rect 8490 7428 8496 7443
rect 8602 7428 8608 7443
rect 8542 7376 8556 7380
rect 8490 6714 8608 7376
rect 8490 6680 8496 6714
rect 8530 6680 8568 6714
rect 8602 6680 8608 6714
rect 8490 6641 8608 6680
rect 8490 6607 8496 6641
rect 8530 6607 8568 6641
rect 8602 6607 8608 6641
rect 8490 6568 8608 6607
rect 8490 6534 8496 6568
rect 8530 6534 8568 6568
rect 8602 6534 8608 6568
rect 8490 6495 8608 6534
rect 8490 6461 8496 6495
rect 8530 6461 8568 6495
rect 8602 6461 8608 6495
rect 8490 6422 8608 6461
rect 8490 5896 8496 6422
rect 8602 5896 8608 6422
rect 8490 5830 8496 5844
rect 8602 5830 8608 5844
rect 8490 5764 8496 5778
rect 8602 5764 8608 5778
rect 8490 5698 8496 5712
rect 8602 5698 8608 5712
rect 8490 5632 8496 5646
rect 8602 5632 8608 5646
rect 8490 5566 8496 5580
rect 8602 5566 8608 5580
rect 8490 5499 8496 5514
rect 8602 5499 8608 5514
rect 8490 5432 8496 5447
rect 8602 5432 8608 5447
rect 8490 5368 8608 5380
rect 8819 14338 8833 14390
rect 9321 14720 9439 14726
rect 9373 14668 9387 14720
rect 9321 14654 9439 14668
rect 9373 14602 9387 14654
rect 9321 14588 9439 14602
rect 9373 14536 9387 14588
rect 9321 14522 9439 14536
rect 9373 14470 9387 14522
rect 9321 14456 9439 14470
rect 9373 14404 9387 14456
rect 9321 14390 9439 14404
rect 8767 14323 8773 14338
rect 8807 14323 8845 14338
rect 8879 14323 8885 14338
rect 8819 14271 8833 14323
rect 8767 14267 8885 14271
rect 8767 14256 8773 14267
rect 8807 14256 8845 14267
rect 8879 14256 8885 14267
rect 8819 14204 8833 14256
rect 8767 14189 8885 14204
rect 8767 14155 8773 14189
rect 8807 14155 8845 14189
rect 8879 14155 8885 14189
rect 8767 14111 8885 14155
rect 8767 14077 8773 14111
rect 8807 14077 8845 14111
rect 8879 14077 8885 14111
rect 8767 14033 8885 14077
rect 8767 13999 8773 14033
rect 8807 13999 8845 14033
rect 8879 13999 8885 14033
rect 8767 13955 8885 13999
rect 8767 13921 8773 13955
rect 8807 13921 8845 13955
rect 8879 13921 8885 13955
rect 8767 13877 8885 13921
rect 8767 13843 8773 13877
rect 8807 13843 8845 13877
rect 8879 13843 8885 13877
rect 8767 13799 8885 13843
rect 8767 13765 8773 13799
rect 8807 13765 8845 13799
rect 8879 13765 8885 13799
rect 8767 13722 8885 13765
rect 8767 13688 8773 13722
rect 8807 13688 8845 13722
rect 8879 13688 8885 13722
rect 8767 13645 8885 13688
rect 8767 13611 8773 13645
rect 8807 13611 8845 13645
rect 8879 13611 8885 13645
rect 8767 13568 8885 13611
rect 8767 13534 8773 13568
rect 8807 13534 8845 13568
rect 8879 13534 8885 13568
rect 8767 13491 8885 13534
rect 8767 13457 8773 13491
rect 8807 13457 8845 13491
rect 8879 13457 8885 13491
rect 8767 13414 8885 13457
rect 8767 13380 8773 13414
rect 8807 13380 8845 13414
rect 8879 13380 8885 13414
rect 8767 12720 8885 13380
rect 8819 12668 8833 12720
rect 8767 12654 8885 12668
rect 8819 12602 8833 12654
rect 8767 12588 8885 12602
rect 8819 12536 8833 12588
rect 8767 12534 8773 12536
rect 8807 12534 8845 12536
rect 8879 12534 8885 12536
rect 8767 12522 8885 12534
rect 8819 12470 8833 12522
rect 8767 12461 8773 12470
rect 8807 12461 8845 12470
rect 8879 12461 8885 12470
rect 8767 12456 8885 12461
rect 8819 12422 8833 12456
rect 8767 12390 8773 12404
rect 8879 12390 8885 12404
rect 8767 12323 8773 12338
rect 8879 12323 8885 12338
rect 8767 12256 8773 12271
rect 8879 12256 8885 12271
rect 8767 11380 8773 12204
rect 8879 11380 8885 12204
rect 8767 10724 8885 11380
rect 8819 10672 8833 10724
rect 8767 10658 8885 10672
rect 8819 10606 8833 10658
rect 8767 10592 8885 10606
rect 8819 10540 8833 10592
rect 8767 10534 8773 10540
rect 8807 10534 8845 10540
rect 8879 10534 8885 10540
rect 8767 10526 8885 10534
rect 8819 10474 8833 10526
rect 8767 10461 8773 10474
rect 8807 10461 8845 10474
rect 8879 10461 8885 10474
rect 8767 10460 8885 10461
rect 8819 10422 8833 10460
rect 8767 10394 8773 10408
rect 8879 10394 8885 10408
rect 8767 10327 8773 10342
rect 8879 10327 8885 10342
rect 8767 10260 8773 10275
rect 8879 10260 8885 10275
rect 8767 9380 8773 10208
rect 8879 9380 8885 10208
rect 8767 8720 8885 9380
rect 8819 8668 8833 8720
rect 8767 8654 8885 8668
rect 8819 8602 8833 8654
rect 8767 8588 8885 8602
rect 8819 8536 8833 8588
rect 8767 8534 8773 8536
rect 8807 8534 8845 8536
rect 8879 8534 8885 8536
rect 8767 8522 8885 8534
rect 8819 8470 8833 8522
rect 8767 8461 8773 8470
rect 8807 8461 8845 8470
rect 8879 8461 8885 8470
rect 8767 8456 8885 8461
rect 8819 8422 8833 8456
rect 8767 8390 8773 8404
rect 8879 8390 8885 8404
rect 8767 8323 8773 8338
rect 8879 8323 8885 8338
rect 8767 8256 8773 8271
rect 8879 8256 8885 8271
rect 8767 7380 8773 8204
rect 8879 7380 8885 8204
rect 8767 6724 8885 7380
rect 8819 6672 8833 6724
rect 8767 6658 8885 6672
rect 8819 6606 8833 6658
rect 8767 6592 8885 6606
rect 8819 6540 8833 6592
rect 8767 6534 8773 6540
rect 8807 6534 8845 6540
rect 8879 6534 8885 6540
rect 8767 6526 8885 6534
rect 8819 6474 8833 6526
rect 8767 6461 8773 6474
rect 8807 6461 8845 6474
rect 8879 6461 8885 6474
rect 8767 6460 8885 6461
rect 8819 6422 8833 6460
rect 8767 6394 8773 6408
rect 8879 6394 8885 6408
rect 8767 6327 8773 6342
rect 8879 6327 8885 6342
rect 8767 6260 8773 6275
rect 8879 6260 8885 6275
rect 8767 5380 8773 6208
rect 8879 5380 8885 6208
tri 8331 5265 8337 5271 sw
tri 8761 5265 8767 5271 se
rect 8767 5265 8885 5380
rect 9044 14345 9162 14357
rect 9044 14311 9050 14345
rect 9084 14311 9122 14345
rect 9156 14311 9162 14345
rect 9044 14267 9162 14311
rect 9044 14233 9050 14267
rect 9084 14233 9122 14267
rect 9156 14233 9162 14267
rect 9044 14189 9162 14233
rect 9044 14155 9050 14189
rect 9084 14155 9122 14189
rect 9156 14155 9162 14189
rect 9044 14111 9162 14155
rect 9044 14077 9050 14111
rect 9084 14077 9122 14111
rect 9156 14077 9162 14111
rect 9044 14033 9162 14077
rect 9044 13999 9050 14033
rect 9084 13999 9122 14033
rect 9156 13999 9162 14033
rect 9044 13955 9162 13999
rect 9044 13921 9050 13955
rect 9084 13921 9122 13955
rect 9156 13921 9162 13955
rect 9044 13892 9162 13921
rect 9096 13840 9110 13892
rect 9044 13826 9162 13840
rect 9096 13774 9110 13826
rect 9044 13765 9050 13774
rect 9084 13765 9122 13774
rect 9156 13765 9162 13774
rect 9044 13760 9162 13765
rect 9096 13708 9110 13760
rect 9044 13694 9050 13708
rect 9084 13694 9122 13708
rect 9156 13694 9162 13708
rect 9096 13642 9110 13694
rect 9044 13628 9050 13642
rect 9084 13628 9122 13642
rect 9156 13628 9162 13642
rect 9096 13576 9110 13628
rect 9044 13568 9162 13576
rect 9044 13562 9050 13568
rect 9084 13562 9122 13568
rect 9156 13562 9162 13568
rect 9096 13510 9110 13562
rect 9044 13495 9162 13510
rect 9096 13443 9110 13495
rect 9044 13428 9162 13443
rect 9096 13376 9110 13428
rect 9044 12714 9162 13376
rect 9044 12680 9050 12714
rect 9084 12680 9122 12714
rect 9156 12680 9162 12714
rect 9044 12641 9162 12680
rect 9044 12607 9050 12641
rect 9084 12607 9122 12641
rect 9156 12607 9162 12641
rect 9044 12568 9162 12607
rect 9044 12534 9050 12568
rect 9084 12534 9122 12568
rect 9156 12534 9162 12568
rect 9044 12495 9162 12534
rect 9044 12461 9050 12495
rect 9084 12461 9122 12495
rect 9156 12461 9162 12495
rect 9044 12422 9162 12461
rect 9044 11892 9050 12422
rect 9156 11892 9162 12422
rect 9044 11826 9050 11840
rect 9156 11826 9162 11840
rect 9044 11760 9050 11774
rect 9156 11760 9162 11774
rect 9044 11694 9050 11708
rect 9156 11694 9162 11708
rect 9044 11628 9050 11642
rect 9156 11628 9162 11642
rect 9044 11562 9050 11576
rect 9156 11562 9162 11576
rect 9044 11495 9050 11510
rect 9156 11495 9162 11510
rect 9044 11428 9050 11443
rect 9156 11428 9162 11443
rect 9096 11376 9110 11380
rect 9044 10714 9162 11376
rect 9044 10680 9050 10714
rect 9084 10680 9122 10714
rect 9156 10680 9162 10714
rect 9044 10641 9162 10680
rect 9044 10607 9050 10641
rect 9084 10607 9122 10641
rect 9156 10607 9162 10641
rect 9044 10568 9162 10607
rect 9044 10534 9050 10568
rect 9084 10534 9122 10568
rect 9156 10534 9162 10568
rect 9044 10495 9162 10534
rect 9044 10461 9050 10495
rect 9084 10461 9122 10495
rect 9156 10461 9162 10495
rect 9044 10422 9162 10461
rect 9044 9896 9050 10422
rect 9156 9896 9162 10422
rect 9044 9830 9050 9844
rect 9156 9830 9162 9844
rect 9044 9764 9050 9778
rect 9156 9764 9162 9778
rect 9044 9698 9050 9712
rect 9156 9698 9162 9712
rect 9044 9632 9050 9646
rect 9156 9632 9162 9646
rect 9044 9566 9050 9580
rect 9156 9566 9162 9580
rect 9044 9499 9050 9514
rect 9156 9499 9162 9514
rect 9044 9432 9050 9447
rect 9156 9432 9162 9447
rect 9044 8714 9162 9380
rect 9044 8680 9050 8714
rect 9084 8680 9122 8714
rect 9156 8680 9162 8714
rect 9044 8641 9162 8680
rect 9044 8607 9050 8641
rect 9084 8607 9122 8641
rect 9156 8607 9162 8641
rect 9044 8568 9162 8607
rect 9044 8534 9050 8568
rect 9084 8534 9122 8568
rect 9156 8534 9162 8568
rect 9044 8495 9162 8534
rect 9044 8461 9050 8495
rect 9084 8461 9122 8495
rect 9156 8461 9162 8495
rect 9044 8422 9162 8461
rect 9044 7892 9050 8422
rect 9156 7892 9162 8422
rect 9044 7826 9050 7840
rect 9156 7826 9162 7840
rect 9044 7760 9050 7774
rect 9156 7760 9162 7774
rect 9044 7694 9050 7708
rect 9156 7694 9162 7708
rect 9044 7628 9050 7642
rect 9156 7628 9162 7642
rect 9044 7562 9050 7576
rect 9156 7562 9162 7576
rect 9044 7495 9050 7510
rect 9156 7495 9162 7510
rect 9044 7428 9050 7443
rect 9156 7428 9162 7443
rect 9096 7376 9110 7380
rect 9044 6714 9162 7376
rect 9044 6680 9050 6714
rect 9084 6680 9122 6714
rect 9156 6680 9162 6714
rect 9044 6641 9162 6680
rect 9044 6607 9050 6641
rect 9084 6607 9122 6641
rect 9156 6607 9162 6641
rect 9044 6568 9162 6607
rect 9044 6534 9050 6568
rect 9084 6534 9122 6568
rect 9156 6534 9162 6568
rect 9044 6495 9162 6534
rect 9044 6461 9050 6495
rect 9084 6461 9122 6495
rect 9156 6461 9162 6495
rect 9044 6422 9162 6461
rect 9044 5896 9050 6422
rect 9156 5896 9162 6422
rect 9044 5830 9050 5844
rect 9156 5830 9162 5844
rect 9044 5764 9050 5778
rect 9156 5764 9162 5778
rect 9044 5698 9050 5712
rect 9156 5698 9162 5712
rect 9044 5632 9050 5646
rect 9156 5632 9162 5646
rect 9044 5566 9050 5580
rect 9156 5566 9162 5580
rect 9044 5499 9050 5514
rect 9156 5499 9162 5514
rect 9044 5432 9050 5447
rect 9156 5432 9162 5447
rect 9044 5368 9162 5380
rect 9373 14338 9387 14390
rect 9875 14720 9993 14726
rect 9927 14668 9941 14720
rect 9875 14654 9993 14668
rect 9927 14602 9941 14654
rect 9875 14588 9993 14602
rect 9927 14536 9941 14588
rect 9875 14522 9993 14536
rect 9927 14470 9941 14522
rect 9875 14456 9993 14470
rect 9927 14404 9941 14456
rect 9875 14390 9993 14404
rect 9321 14323 9327 14338
rect 9361 14323 9399 14338
rect 9433 14323 9439 14338
rect 9373 14271 9387 14323
rect 9321 14267 9439 14271
rect 9321 14256 9327 14267
rect 9361 14256 9399 14267
rect 9433 14256 9439 14267
rect 9373 14204 9387 14256
rect 9321 14189 9439 14204
rect 9321 14155 9327 14189
rect 9361 14155 9399 14189
rect 9433 14155 9439 14189
rect 9321 14111 9439 14155
rect 9321 14077 9327 14111
rect 9361 14077 9399 14111
rect 9433 14077 9439 14111
rect 9321 14033 9439 14077
rect 9321 13999 9327 14033
rect 9361 13999 9399 14033
rect 9433 13999 9439 14033
rect 9321 13955 9439 13999
rect 9321 13921 9327 13955
rect 9361 13921 9399 13955
rect 9433 13921 9439 13955
rect 9321 13877 9439 13921
rect 9321 13843 9327 13877
rect 9361 13843 9399 13877
rect 9433 13843 9439 13877
rect 9321 13799 9439 13843
rect 9321 13765 9327 13799
rect 9361 13765 9399 13799
rect 9433 13765 9439 13799
rect 9321 13722 9439 13765
rect 9321 13688 9327 13722
rect 9361 13688 9399 13722
rect 9433 13688 9439 13722
rect 9321 13645 9439 13688
rect 9321 13611 9327 13645
rect 9361 13611 9399 13645
rect 9433 13611 9439 13645
rect 9321 13568 9439 13611
rect 9321 13534 9327 13568
rect 9361 13534 9399 13568
rect 9433 13534 9439 13568
rect 9321 13491 9439 13534
rect 9321 13457 9327 13491
rect 9361 13457 9399 13491
rect 9433 13457 9439 13491
rect 9321 13414 9439 13457
rect 9321 13380 9327 13414
rect 9361 13380 9399 13414
rect 9433 13380 9439 13414
rect 9321 12720 9439 13380
rect 9373 12668 9387 12720
rect 9321 12654 9439 12668
rect 9373 12602 9387 12654
rect 9321 12588 9439 12602
rect 9373 12536 9387 12588
rect 9321 12534 9327 12536
rect 9361 12534 9399 12536
rect 9433 12534 9439 12536
rect 9321 12522 9439 12534
rect 9373 12470 9387 12522
rect 9321 12461 9327 12470
rect 9361 12461 9399 12470
rect 9433 12461 9439 12470
rect 9321 12456 9439 12461
rect 9373 12422 9387 12456
rect 9321 12390 9327 12404
rect 9433 12390 9439 12404
rect 9321 12323 9327 12338
rect 9433 12323 9439 12338
rect 9321 12256 9327 12271
rect 9433 12256 9439 12271
rect 9321 11380 9327 12204
rect 9433 11380 9439 12204
rect 9321 10724 9439 11380
rect 9373 10672 9387 10724
rect 9321 10658 9439 10672
rect 9373 10606 9387 10658
rect 9321 10592 9439 10606
rect 9373 10540 9387 10592
rect 9321 10534 9327 10540
rect 9361 10534 9399 10540
rect 9433 10534 9439 10540
rect 9321 10526 9439 10534
rect 9373 10474 9387 10526
rect 9321 10461 9327 10474
rect 9361 10461 9399 10474
rect 9433 10461 9439 10474
rect 9321 10460 9439 10461
rect 9373 10422 9387 10460
rect 9321 10394 9327 10408
rect 9433 10394 9439 10408
rect 9321 10327 9327 10342
rect 9433 10327 9439 10342
rect 9321 10260 9327 10275
rect 9433 10260 9439 10275
rect 9321 9380 9327 10208
rect 9433 9380 9439 10208
rect 9321 8720 9439 9380
rect 9373 8668 9387 8720
rect 9321 8654 9439 8668
rect 9373 8602 9387 8654
rect 9321 8588 9439 8602
rect 9373 8536 9387 8588
rect 9321 8534 9327 8536
rect 9361 8534 9399 8536
rect 9433 8534 9439 8536
rect 9321 8522 9439 8534
rect 9373 8470 9387 8522
rect 9321 8461 9327 8470
rect 9361 8461 9399 8470
rect 9433 8461 9439 8470
rect 9321 8456 9439 8461
rect 9373 8422 9387 8456
rect 9321 8390 9327 8404
rect 9433 8390 9439 8404
rect 9321 8323 9327 8338
rect 9433 8323 9439 8338
rect 9321 8256 9327 8271
rect 9433 8256 9439 8271
rect 9321 7380 9327 8204
rect 9433 7380 9439 8204
rect 9321 6724 9439 7380
rect 9373 6672 9387 6724
rect 9321 6658 9439 6672
rect 9373 6606 9387 6658
rect 9321 6592 9439 6606
rect 9373 6540 9387 6592
rect 9321 6534 9327 6540
rect 9361 6534 9399 6540
rect 9433 6534 9439 6540
rect 9321 6526 9439 6534
rect 9373 6474 9387 6526
rect 9321 6461 9327 6474
rect 9361 6461 9399 6474
rect 9433 6461 9439 6474
rect 9321 6460 9439 6461
rect 9373 6422 9387 6460
rect 9321 6394 9327 6408
rect 9433 6394 9439 6408
rect 9321 6327 9327 6342
rect 9433 6327 9439 6342
rect 9321 6260 9327 6275
rect 9433 6260 9439 6275
rect 9321 5380 9327 6208
rect 9433 5380 9439 6208
tri 8885 5265 8891 5271 sw
tri 9315 5265 9321 5271 se
rect 9321 5265 9439 5380
rect 9598 14345 9716 14357
rect 9598 14311 9604 14345
rect 9638 14311 9676 14345
rect 9710 14311 9716 14345
rect 9598 14267 9716 14311
rect 9598 14233 9604 14267
rect 9638 14233 9676 14267
rect 9710 14233 9716 14267
rect 9598 14189 9716 14233
rect 9598 14155 9604 14189
rect 9638 14155 9676 14189
rect 9710 14155 9716 14189
rect 9598 14111 9716 14155
rect 9598 14077 9604 14111
rect 9638 14077 9676 14111
rect 9710 14077 9716 14111
rect 9598 14033 9716 14077
rect 9598 13999 9604 14033
rect 9638 13999 9676 14033
rect 9710 13999 9716 14033
rect 9598 13955 9716 13999
rect 9598 13921 9604 13955
rect 9638 13921 9676 13955
rect 9710 13921 9716 13955
rect 9598 13892 9716 13921
rect 9650 13840 9664 13892
rect 9598 13826 9716 13840
rect 9650 13774 9664 13826
rect 9598 13765 9604 13774
rect 9638 13765 9676 13774
rect 9710 13765 9716 13774
rect 9598 13760 9716 13765
rect 9650 13708 9664 13760
rect 9598 13694 9604 13708
rect 9638 13694 9676 13708
rect 9710 13694 9716 13708
rect 9650 13642 9664 13694
rect 9598 13628 9604 13642
rect 9638 13628 9676 13642
rect 9710 13628 9716 13642
rect 9650 13576 9664 13628
rect 9598 13568 9716 13576
rect 9598 13562 9604 13568
rect 9638 13562 9676 13568
rect 9710 13562 9716 13568
rect 9650 13510 9664 13562
rect 9598 13495 9716 13510
rect 9650 13443 9664 13495
rect 9598 13428 9716 13443
rect 9650 13376 9664 13428
rect 9598 12714 9716 13376
rect 9598 12680 9604 12714
rect 9638 12680 9676 12714
rect 9710 12680 9716 12714
rect 9598 12641 9716 12680
rect 9598 12607 9604 12641
rect 9638 12607 9676 12641
rect 9710 12607 9716 12641
rect 9598 12568 9716 12607
rect 9598 12534 9604 12568
rect 9638 12534 9676 12568
rect 9710 12534 9716 12568
rect 9598 12495 9716 12534
rect 9598 12461 9604 12495
rect 9638 12461 9676 12495
rect 9710 12461 9716 12495
rect 9598 12422 9716 12461
rect 9598 11892 9604 12422
rect 9710 11892 9716 12422
rect 9598 11826 9604 11840
rect 9710 11826 9716 11840
rect 9598 11760 9604 11774
rect 9710 11760 9716 11774
rect 9598 11694 9604 11708
rect 9710 11694 9716 11708
rect 9598 11628 9604 11642
rect 9710 11628 9716 11642
rect 9598 11562 9604 11576
rect 9710 11562 9716 11576
rect 9598 11495 9604 11510
rect 9710 11495 9716 11510
rect 9598 11428 9604 11443
rect 9710 11428 9716 11443
rect 9650 11376 9664 11380
rect 9598 10714 9716 11376
rect 9598 10680 9604 10714
rect 9638 10680 9676 10714
rect 9710 10680 9716 10714
rect 9598 10641 9716 10680
rect 9598 10607 9604 10641
rect 9638 10607 9676 10641
rect 9710 10607 9716 10641
rect 9598 10568 9716 10607
rect 9598 10534 9604 10568
rect 9638 10534 9676 10568
rect 9710 10534 9716 10568
rect 9598 10495 9716 10534
rect 9598 10461 9604 10495
rect 9638 10461 9676 10495
rect 9710 10461 9716 10495
rect 9598 10422 9716 10461
rect 9598 9896 9604 10422
rect 9710 9896 9716 10422
rect 9598 9830 9604 9844
rect 9710 9830 9716 9844
rect 9598 9764 9604 9778
rect 9710 9764 9716 9778
rect 9598 9698 9604 9712
rect 9710 9698 9716 9712
rect 9598 9632 9604 9646
rect 9710 9632 9716 9646
rect 9598 9566 9604 9580
rect 9710 9566 9716 9580
rect 9598 9499 9604 9514
rect 9710 9499 9716 9514
rect 9598 9432 9604 9447
rect 9710 9432 9716 9447
rect 9598 8714 9716 9380
rect 9598 8680 9604 8714
rect 9638 8680 9676 8714
rect 9710 8680 9716 8714
rect 9598 8641 9716 8680
rect 9598 8607 9604 8641
rect 9638 8607 9676 8641
rect 9710 8607 9716 8641
rect 9598 8568 9716 8607
rect 9598 8534 9604 8568
rect 9638 8534 9676 8568
rect 9710 8534 9716 8568
rect 9598 8495 9716 8534
rect 9598 8461 9604 8495
rect 9638 8461 9676 8495
rect 9710 8461 9716 8495
rect 9598 8422 9716 8461
rect 9598 7892 9604 8422
rect 9710 7892 9716 8422
rect 9598 7826 9604 7840
rect 9710 7826 9716 7840
rect 9598 7760 9604 7774
rect 9710 7760 9716 7774
rect 9598 7694 9604 7708
rect 9710 7694 9716 7708
rect 9598 7628 9604 7642
rect 9710 7628 9716 7642
rect 9598 7562 9604 7576
rect 9710 7562 9716 7576
rect 9598 7495 9604 7510
rect 9710 7495 9716 7510
rect 9598 7428 9604 7443
rect 9710 7428 9716 7443
rect 9650 7376 9664 7380
rect 9598 6714 9716 7376
rect 9598 6680 9604 6714
rect 9638 6680 9676 6714
rect 9710 6680 9716 6714
rect 9598 6641 9716 6680
rect 9598 6607 9604 6641
rect 9638 6607 9676 6641
rect 9710 6607 9716 6641
rect 9598 6568 9716 6607
rect 9598 6534 9604 6568
rect 9638 6534 9676 6568
rect 9710 6534 9716 6568
rect 9598 6495 9716 6534
rect 9598 6461 9604 6495
rect 9638 6461 9676 6495
rect 9710 6461 9716 6495
rect 9598 6422 9716 6461
rect 9598 5896 9604 6422
rect 9710 5896 9716 6422
rect 9598 5830 9604 5844
rect 9710 5830 9716 5844
rect 9598 5764 9604 5778
rect 9710 5764 9716 5778
rect 9598 5698 9604 5712
rect 9710 5698 9716 5712
rect 9598 5632 9604 5646
rect 9710 5632 9716 5646
rect 9598 5566 9604 5580
rect 9710 5566 9716 5580
rect 9598 5499 9604 5514
rect 9710 5499 9716 5514
rect 9598 5432 9604 5447
rect 9710 5432 9716 5447
rect 9598 5368 9716 5380
rect 9927 14338 9941 14390
rect 10429 14720 10547 14726
rect 10481 14668 10495 14720
rect 10429 14654 10547 14668
rect 10481 14602 10495 14654
rect 10429 14588 10547 14602
rect 10481 14536 10495 14588
rect 10429 14522 10547 14536
rect 10481 14470 10495 14522
rect 10429 14456 10547 14470
rect 10481 14404 10495 14456
rect 10429 14390 10547 14404
rect 9875 14323 9881 14338
rect 9915 14323 9953 14338
rect 9987 14323 9993 14338
rect 9927 14271 9941 14323
rect 9875 14267 9993 14271
rect 9875 14256 9881 14267
rect 9915 14256 9953 14267
rect 9987 14256 9993 14267
rect 9927 14204 9941 14256
rect 9875 14189 9993 14204
rect 9875 14155 9881 14189
rect 9915 14155 9953 14189
rect 9987 14155 9993 14189
rect 9875 14111 9993 14155
rect 9875 14077 9881 14111
rect 9915 14077 9953 14111
rect 9987 14077 9993 14111
rect 9875 14033 9993 14077
rect 9875 13999 9881 14033
rect 9915 13999 9953 14033
rect 9987 13999 9993 14033
rect 9875 13955 9993 13999
rect 9875 13921 9881 13955
rect 9915 13921 9953 13955
rect 9987 13921 9993 13955
rect 9875 13877 9993 13921
rect 9875 13843 9881 13877
rect 9915 13843 9953 13877
rect 9987 13843 9993 13877
rect 9875 13799 9993 13843
rect 9875 13765 9881 13799
rect 9915 13765 9953 13799
rect 9987 13765 9993 13799
rect 9875 13722 9993 13765
rect 9875 13688 9881 13722
rect 9915 13688 9953 13722
rect 9987 13688 9993 13722
rect 9875 13645 9993 13688
rect 9875 13611 9881 13645
rect 9915 13611 9953 13645
rect 9987 13611 9993 13645
rect 9875 13568 9993 13611
rect 9875 13534 9881 13568
rect 9915 13534 9953 13568
rect 9987 13534 9993 13568
rect 9875 13491 9993 13534
rect 9875 13457 9881 13491
rect 9915 13457 9953 13491
rect 9987 13457 9993 13491
rect 9875 13414 9993 13457
rect 9875 13380 9881 13414
rect 9915 13380 9953 13414
rect 9987 13380 9993 13414
rect 9875 12720 9993 13380
rect 9927 12668 9941 12720
rect 9875 12654 9993 12668
rect 9927 12602 9941 12654
rect 9875 12588 9993 12602
rect 9927 12536 9941 12588
rect 9875 12534 9881 12536
rect 9915 12534 9953 12536
rect 9987 12534 9993 12536
rect 9875 12522 9993 12534
rect 9927 12470 9941 12522
rect 9875 12461 9881 12470
rect 9915 12461 9953 12470
rect 9987 12461 9993 12470
rect 9875 12456 9993 12461
rect 9927 12422 9941 12456
rect 9875 12390 9881 12404
rect 9987 12390 9993 12404
rect 9875 12323 9881 12338
rect 9987 12323 9993 12338
rect 9875 12256 9881 12271
rect 9987 12256 9993 12271
rect 9875 11380 9881 12204
rect 9987 11380 9993 12204
rect 9875 10724 9993 11380
rect 9927 10672 9941 10724
rect 9875 10658 9993 10672
rect 9927 10606 9941 10658
rect 9875 10592 9993 10606
rect 9927 10540 9941 10592
rect 9875 10534 9881 10540
rect 9915 10534 9953 10540
rect 9987 10534 9993 10540
rect 9875 10526 9993 10534
rect 9927 10474 9941 10526
rect 9875 10461 9881 10474
rect 9915 10461 9953 10474
rect 9987 10461 9993 10474
rect 9875 10460 9993 10461
rect 9927 10422 9941 10460
rect 9875 10394 9881 10408
rect 9987 10394 9993 10408
rect 9875 10327 9881 10342
rect 9987 10327 9993 10342
rect 9875 10260 9881 10275
rect 9987 10260 9993 10275
rect 9875 9380 9881 10208
rect 9987 9380 9993 10208
rect 9875 8720 9993 9380
rect 9927 8668 9941 8720
rect 9875 8654 9993 8668
rect 9927 8602 9941 8654
rect 9875 8588 9993 8602
rect 9927 8536 9941 8588
rect 9875 8534 9881 8536
rect 9915 8534 9953 8536
rect 9987 8534 9993 8536
rect 9875 8522 9993 8534
rect 9927 8470 9941 8522
rect 9875 8461 9881 8470
rect 9915 8461 9953 8470
rect 9987 8461 9993 8470
rect 9875 8456 9993 8461
rect 9927 8422 9941 8456
rect 9875 8390 9881 8404
rect 9987 8390 9993 8404
rect 9875 8323 9881 8338
rect 9987 8323 9993 8338
rect 9875 8256 9881 8271
rect 9987 8256 9993 8271
rect 9875 7380 9881 8204
rect 9987 7380 9993 8204
rect 9875 6724 9993 7380
rect 9927 6672 9941 6724
rect 9875 6658 9993 6672
rect 9927 6606 9941 6658
rect 9875 6592 9993 6606
rect 9927 6540 9941 6592
rect 9875 6534 9881 6540
rect 9915 6534 9953 6540
rect 9987 6534 9993 6540
rect 9875 6526 9993 6534
rect 9927 6474 9941 6526
rect 9875 6461 9881 6474
rect 9915 6461 9953 6474
rect 9987 6461 9993 6474
rect 9875 6460 9993 6461
rect 9927 6422 9941 6460
rect 9875 6394 9881 6408
rect 9987 6394 9993 6408
rect 9875 6327 9881 6342
rect 9987 6327 9993 6342
rect 9875 6260 9881 6275
rect 9987 6260 9993 6275
rect 9875 5380 9881 6208
rect 9987 5380 9993 6208
tri 9439 5265 9445 5271 sw
tri 9869 5265 9875 5271 se
rect 9875 5265 9993 5380
rect 10152 14345 10270 14357
rect 10152 14311 10158 14345
rect 10192 14311 10230 14345
rect 10264 14311 10270 14345
rect 10152 14267 10270 14311
rect 10152 14233 10158 14267
rect 10192 14233 10230 14267
rect 10264 14233 10270 14267
rect 10152 14189 10270 14233
rect 10152 14155 10158 14189
rect 10192 14155 10230 14189
rect 10264 14155 10270 14189
rect 10152 14111 10270 14155
rect 10152 14077 10158 14111
rect 10192 14077 10230 14111
rect 10264 14077 10270 14111
rect 10152 14033 10270 14077
rect 10152 13999 10158 14033
rect 10192 13999 10230 14033
rect 10264 13999 10270 14033
rect 10152 13955 10270 13999
rect 10152 13921 10158 13955
rect 10192 13921 10230 13955
rect 10264 13921 10270 13955
rect 10152 13892 10270 13921
rect 10204 13840 10218 13892
rect 10152 13826 10270 13840
rect 10204 13774 10218 13826
rect 10152 13765 10158 13774
rect 10192 13765 10230 13774
rect 10264 13765 10270 13774
rect 10152 13760 10270 13765
rect 10204 13708 10218 13760
rect 10152 13694 10158 13708
rect 10192 13694 10230 13708
rect 10264 13694 10270 13708
rect 10204 13642 10218 13694
rect 10152 13628 10158 13642
rect 10192 13628 10230 13642
rect 10264 13628 10270 13642
rect 10204 13576 10218 13628
rect 10152 13568 10270 13576
rect 10152 13562 10158 13568
rect 10192 13562 10230 13568
rect 10264 13562 10270 13568
rect 10204 13510 10218 13562
rect 10152 13495 10270 13510
rect 10204 13443 10218 13495
rect 10152 13428 10270 13443
rect 10204 13376 10218 13428
rect 10152 12714 10270 13376
rect 10152 12680 10158 12714
rect 10192 12680 10230 12714
rect 10264 12680 10270 12714
rect 10152 12641 10270 12680
rect 10152 12607 10158 12641
rect 10192 12607 10230 12641
rect 10264 12607 10270 12641
rect 10152 12568 10270 12607
rect 10152 12534 10158 12568
rect 10192 12534 10230 12568
rect 10264 12534 10270 12568
rect 10152 12495 10270 12534
rect 10152 12461 10158 12495
rect 10192 12461 10230 12495
rect 10264 12461 10270 12495
rect 10152 12422 10270 12461
rect 10152 11892 10158 12422
rect 10264 11892 10270 12422
rect 10152 11826 10158 11840
rect 10264 11826 10270 11840
rect 10152 11760 10158 11774
rect 10264 11760 10270 11774
rect 10152 11694 10158 11708
rect 10264 11694 10270 11708
rect 10152 11628 10158 11642
rect 10264 11628 10270 11642
rect 10152 11562 10158 11576
rect 10264 11562 10270 11576
rect 10152 11495 10158 11510
rect 10264 11495 10270 11510
rect 10152 11428 10158 11443
rect 10264 11428 10270 11443
rect 10204 11376 10218 11380
rect 10152 10714 10270 11376
rect 10152 10680 10158 10714
rect 10192 10680 10230 10714
rect 10264 10680 10270 10714
rect 10152 10641 10270 10680
rect 10152 10607 10158 10641
rect 10192 10607 10230 10641
rect 10264 10607 10270 10641
rect 10152 10568 10270 10607
rect 10152 10534 10158 10568
rect 10192 10534 10230 10568
rect 10264 10534 10270 10568
rect 10152 10495 10270 10534
rect 10152 10461 10158 10495
rect 10192 10461 10230 10495
rect 10264 10461 10270 10495
rect 10152 10422 10270 10461
rect 10152 9896 10158 10422
rect 10264 9896 10270 10422
rect 10152 9830 10158 9844
rect 10264 9830 10270 9844
rect 10152 9764 10158 9778
rect 10264 9764 10270 9778
rect 10152 9698 10158 9712
rect 10264 9698 10270 9712
rect 10152 9632 10158 9646
rect 10264 9632 10270 9646
rect 10152 9566 10158 9580
rect 10264 9566 10270 9580
rect 10152 9499 10158 9514
rect 10264 9499 10270 9514
rect 10152 9432 10158 9447
rect 10264 9432 10270 9447
rect 10152 8714 10270 9380
rect 10152 8680 10158 8714
rect 10192 8680 10230 8714
rect 10264 8680 10270 8714
rect 10152 8641 10270 8680
rect 10152 8607 10158 8641
rect 10192 8607 10230 8641
rect 10264 8607 10270 8641
rect 10152 8568 10270 8607
rect 10152 8534 10158 8568
rect 10192 8534 10230 8568
rect 10264 8534 10270 8568
rect 10152 8495 10270 8534
rect 10152 8461 10158 8495
rect 10192 8461 10230 8495
rect 10264 8461 10270 8495
rect 10152 8422 10270 8461
rect 10152 7892 10158 8422
rect 10264 7892 10270 8422
rect 10152 7826 10158 7840
rect 10264 7826 10270 7840
rect 10152 7760 10158 7774
rect 10264 7760 10270 7774
rect 10152 7694 10158 7708
rect 10264 7694 10270 7708
rect 10152 7628 10158 7642
rect 10264 7628 10270 7642
rect 10152 7562 10158 7576
rect 10264 7562 10270 7576
rect 10152 7495 10158 7510
rect 10264 7495 10270 7510
rect 10152 7428 10158 7443
rect 10264 7428 10270 7443
rect 10204 7376 10218 7380
rect 10152 6714 10270 7376
rect 10152 6680 10158 6714
rect 10192 6680 10230 6714
rect 10264 6680 10270 6714
rect 10152 6641 10270 6680
rect 10152 6607 10158 6641
rect 10192 6607 10230 6641
rect 10264 6607 10270 6641
rect 10152 6568 10270 6607
rect 10152 6534 10158 6568
rect 10192 6534 10230 6568
rect 10264 6534 10270 6568
rect 10152 6495 10270 6534
rect 10152 6461 10158 6495
rect 10192 6461 10230 6495
rect 10264 6461 10270 6495
rect 10152 6422 10270 6461
rect 10152 5896 10158 6422
rect 10264 5896 10270 6422
rect 10152 5830 10158 5844
rect 10264 5830 10270 5844
rect 10152 5764 10158 5778
rect 10264 5764 10270 5778
rect 10152 5698 10158 5712
rect 10264 5698 10270 5712
rect 10152 5632 10158 5646
rect 10264 5632 10270 5646
rect 10152 5566 10158 5580
rect 10264 5566 10270 5580
rect 10152 5499 10158 5514
rect 10264 5499 10270 5514
rect 10152 5432 10158 5447
rect 10264 5432 10270 5447
rect 10152 5368 10270 5380
rect 10481 14338 10495 14390
rect 10983 14720 11101 14726
rect 11035 14668 11049 14720
rect 10983 14654 11101 14668
rect 11035 14602 11049 14654
rect 10983 14588 11101 14602
rect 11035 14536 11049 14588
rect 10983 14522 11101 14536
rect 11035 14470 11049 14522
rect 10983 14456 11101 14470
rect 11035 14404 11049 14456
rect 10983 14390 11101 14404
rect 10429 14323 10435 14338
rect 10469 14323 10507 14338
rect 10541 14323 10547 14338
rect 10481 14271 10495 14323
rect 10429 14267 10547 14271
rect 10429 14256 10435 14267
rect 10469 14256 10507 14267
rect 10541 14256 10547 14267
rect 10481 14204 10495 14256
rect 10429 14189 10547 14204
rect 10429 14155 10435 14189
rect 10469 14155 10507 14189
rect 10541 14155 10547 14189
rect 10429 14111 10547 14155
rect 10429 14077 10435 14111
rect 10469 14077 10507 14111
rect 10541 14077 10547 14111
rect 10429 14033 10547 14077
rect 10429 13999 10435 14033
rect 10469 13999 10507 14033
rect 10541 13999 10547 14033
rect 10429 13955 10547 13999
rect 10429 13921 10435 13955
rect 10469 13921 10507 13955
rect 10541 13921 10547 13955
rect 10429 13877 10547 13921
rect 10429 13843 10435 13877
rect 10469 13843 10507 13877
rect 10541 13843 10547 13877
rect 10429 13799 10547 13843
rect 10429 13765 10435 13799
rect 10469 13765 10507 13799
rect 10541 13765 10547 13799
rect 10429 13722 10547 13765
rect 10429 13688 10435 13722
rect 10469 13688 10507 13722
rect 10541 13688 10547 13722
rect 10429 13645 10547 13688
rect 10429 13611 10435 13645
rect 10469 13611 10507 13645
rect 10541 13611 10547 13645
rect 10429 13568 10547 13611
rect 10429 13534 10435 13568
rect 10469 13534 10507 13568
rect 10541 13534 10547 13568
rect 10429 13491 10547 13534
rect 10429 13457 10435 13491
rect 10469 13457 10507 13491
rect 10541 13457 10547 13491
rect 10429 13414 10547 13457
rect 10429 13380 10435 13414
rect 10469 13380 10507 13414
rect 10541 13380 10547 13414
rect 10429 12720 10547 13380
rect 10481 12668 10495 12720
rect 10429 12654 10547 12668
rect 10481 12602 10495 12654
rect 10429 12588 10547 12602
rect 10481 12536 10495 12588
rect 10429 12534 10435 12536
rect 10469 12534 10507 12536
rect 10541 12534 10547 12536
rect 10429 12522 10547 12534
rect 10481 12470 10495 12522
rect 10429 12461 10435 12470
rect 10469 12461 10507 12470
rect 10541 12461 10547 12470
rect 10429 12456 10547 12461
rect 10481 12422 10495 12456
rect 10429 12390 10435 12404
rect 10541 12390 10547 12404
rect 10429 12323 10435 12338
rect 10541 12323 10547 12338
rect 10429 12256 10435 12271
rect 10541 12256 10547 12271
rect 10429 11380 10435 12204
rect 10541 11380 10547 12204
rect 10429 10724 10547 11380
rect 10481 10672 10495 10724
rect 10429 10658 10547 10672
rect 10481 10606 10495 10658
rect 10429 10592 10547 10606
rect 10481 10540 10495 10592
rect 10429 10534 10435 10540
rect 10469 10534 10507 10540
rect 10541 10534 10547 10540
rect 10429 10526 10547 10534
rect 10481 10474 10495 10526
rect 10429 10461 10435 10474
rect 10469 10461 10507 10474
rect 10541 10461 10547 10474
rect 10429 10460 10547 10461
rect 10481 10422 10495 10460
rect 10429 10394 10435 10408
rect 10541 10394 10547 10408
rect 10429 10327 10435 10342
rect 10541 10327 10547 10342
rect 10429 10260 10435 10275
rect 10541 10260 10547 10275
rect 10429 9380 10435 10208
rect 10541 9380 10547 10208
rect 10429 8720 10547 9380
rect 10481 8668 10495 8720
rect 10429 8654 10547 8668
rect 10481 8602 10495 8654
rect 10429 8588 10547 8602
rect 10481 8536 10495 8588
rect 10429 8534 10435 8536
rect 10469 8534 10507 8536
rect 10541 8534 10547 8536
rect 10429 8522 10547 8534
rect 10481 8470 10495 8522
rect 10429 8461 10435 8470
rect 10469 8461 10507 8470
rect 10541 8461 10547 8470
rect 10429 8456 10547 8461
rect 10481 8422 10495 8456
rect 10429 8390 10435 8404
rect 10541 8390 10547 8404
rect 10429 8323 10435 8338
rect 10541 8323 10547 8338
rect 10429 8256 10435 8271
rect 10541 8256 10547 8271
rect 10429 7380 10435 8204
rect 10541 7380 10547 8204
rect 10429 6724 10547 7380
rect 10481 6672 10495 6724
rect 10429 6658 10547 6672
rect 10481 6606 10495 6658
rect 10429 6592 10547 6606
rect 10481 6540 10495 6592
rect 10429 6534 10435 6540
rect 10469 6534 10507 6540
rect 10541 6534 10547 6540
rect 10429 6526 10547 6534
rect 10481 6474 10495 6526
rect 10429 6461 10435 6474
rect 10469 6461 10507 6474
rect 10541 6461 10547 6474
rect 10429 6460 10547 6461
rect 10481 6422 10495 6460
rect 10429 6394 10435 6408
rect 10541 6394 10547 6408
rect 10429 6327 10435 6342
rect 10541 6327 10547 6342
rect 10429 6260 10435 6275
rect 10541 6260 10547 6275
rect 10429 5380 10435 6208
rect 10541 5380 10547 6208
tri 9993 5265 9999 5271 sw
tri 10423 5265 10429 5271 se
rect 10429 5265 10547 5380
rect 10706 14345 10824 14357
rect 10706 14311 10712 14345
rect 10746 14311 10784 14345
rect 10818 14311 10824 14345
rect 10706 14267 10824 14311
rect 10706 14233 10712 14267
rect 10746 14233 10784 14267
rect 10818 14233 10824 14267
rect 10706 14189 10824 14233
rect 10706 14155 10712 14189
rect 10746 14155 10784 14189
rect 10818 14155 10824 14189
rect 10706 14111 10824 14155
rect 10706 14077 10712 14111
rect 10746 14077 10784 14111
rect 10818 14077 10824 14111
rect 10706 14033 10824 14077
rect 10706 13999 10712 14033
rect 10746 13999 10784 14033
rect 10818 13999 10824 14033
rect 10706 13955 10824 13999
rect 10706 13921 10712 13955
rect 10746 13921 10784 13955
rect 10818 13921 10824 13955
rect 10706 13892 10824 13921
rect 10758 13840 10772 13892
rect 10706 13826 10824 13840
rect 10758 13774 10772 13826
rect 10706 13765 10712 13774
rect 10746 13765 10784 13774
rect 10818 13765 10824 13774
rect 10706 13760 10824 13765
rect 10758 13708 10772 13760
rect 10706 13694 10712 13708
rect 10746 13694 10784 13708
rect 10818 13694 10824 13708
rect 10758 13642 10772 13694
rect 10706 13628 10712 13642
rect 10746 13628 10784 13642
rect 10818 13628 10824 13642
rect 10758 13576 10772 13628
rect 10706 13568 10824 13576
rect 10706 13562 10712 13568
rect 10746 13562 10784 13568
rect 10818 13562 10824 13568
rect 10758 13510 10772 13562
rect 10706 13495 10824 13510
rect 10758 13443 10772 13495
rect 10706 13428 10824 13443
rect 10758 13376 10772 13428
rect 10706 12714 10824 13376
rect 10706 12680 10712 12714
rect 10746 12680 10784 12714
rect 10818 12680 10824 12714
rect 10706 12641 10824 12680
rect 10706 12607 10712 12641
rect 10746 12607 10784 12641
rect 10818 12607 10824 12641
rect 10706 12568 10824 12607
rect 10706 12534 10712 12568
rect 10746 12534 10784 12568
rect 10818 12534 10824 12568
rect 10706 12495 10824 12534
rect 10706 12461 10712 12495
rect 10746 12461 10784 12495
rect 10818 12461 10824 12495
rect 10706 12422 10824 12461
rect 10706 11892 10712 12422
rect 10818 11892 10824 12422
rect 10706 11826 10712 11840
rect 10818 11826 10824 11840
rect 10706 11760 10712 11774
rect 10818 11760 10824 11774
rect 10706 11694 10712 11708
rect 10818 11694 10824 11708
rect 10706 11628 10712 11642
rect 10818 11628 10824 11642
rect 10706 11562 10712 11576
rect 10818 11562 10824 11576
rect 10706 11495 10712 11510
rect 10818 11495 10824 11510
rect 10706 11428 10712 11443
rect 10818 11428 10824 11443
rect 10758 11376 10772 11380
rect 10706 10714 10824 11376
rect 10706 10680 10712 10714
rect 10746 10680 10784 10714
rect 10818 10680 10824 10714
rect 10706 10641 10824 10680
rect 10706 10607 10712 10641
rect 10746 10607 10784 10641
rect 10818 10607 10824 10641
rect 10706 10568 10824 10607
rect 10706 10534 10712 10568
rect 10746 10534 10784 10568
rect 10818 10534 10824 10568
rect 10706 10495 10824 10534
rect 10706 10461 10712 10495
rect 10746 10461 10784 10495
rect 10818 10461 10824 10495
rect 10706 10422 10824 10461
rect 10706 9896 10712 10422
rect 10818 9896 10824 10422
rect 10706 9830 10712 9844
rect 10818 9830 10824 9844
rect 10706 9764 10712 9778
rect 10818 9764 10824 9778
rect 10706 9698 10712 9712
rect 10818 9698 10824 9712
rect 10706 9632 10712 9646
rect 10818 9632 10824 9646
rect 10706 9566 10712 9580
rect 10818 9566 10824 9580
rect 10706 9499 10712 9514
rect 10818 9499 10824 9514
rect 10706 9432 10712 9447
rect 10818 9432 10824 9447
rect 10706 8714 10824 9380
rect 10706 8680 10712 8714
rect 10746 8680 10784 8714
rect 10818 8680 10824 8714
rect 10706 8641 10824 8680
rect 10706 8607 10712 8641
rect 10746 8607 10784 8641
rect 10818 8607 10824 8641
rect 10706 8568 10824 8607
rect 10706 8534 10712 8568
rect 10746 8534 10784 8568
rect 10818 8534 10824 8568
rect 10706 8495 10824 8534
rect 10706 8461 10712 8495
rect 10746 8461 10784 8495
rect 10818 8461 10824 8495
rect 10706 8422 10824 8461
rect 10706 7892 10712 8422
rect 10818 7892 10824 8422
rect 10706 7826 10712 7840
rect 10818 7826 10824 7840
rect 10706 7760 10712 7774
rect 10818 7760 10824 7774
rect 10706 7694 10712 7708
rect 10818 7694 10824 7708
rect 10706 7628 10712 7642
rect 10818 7628 10824 7642
rect 10706 7562 10712 7576
rect 10818 7562 10824 7576
rect 10706 7495 10712 7510
rect 10818 7495 10824 7510
rect 10706 7428 10712 7443
rect 10818 7428 10824 7443
rect 10758 7376 10772 7380
rect 10706 6714 10824 7376
rect 10706 6680 10712 6714
rect 10746 6680 10784 6714
rect 10818 6680 10824 6714
rect 10706 6641 10824 6680
rect 10706 6607 10712 6641
rect 10746 6607 10784 6641
rect 10818 6607 10824 6641
rect 10706 6568 10824 6607
rect 10706 6534 10712 6568
rect 10746 6534 10784 6568
rect 10818 6534 10824 6568
rect 10706 6495 10824 6534
rect 10706 6461 10712 6495
rect 10746 6461 10784 6495
rect 10818 6461 10824 6495
rect 10706 6422 10824 6461
rect 10706 5896 10712 6422
rect 10818 5896 10824 6422
rect 10706 5830 10712 5844
rect 10818 5830 10824 5844
rect 10706 5764 10712 5778
rect 10818 5764 10824 5778
rect 10706 5698 10712 5712
rect 10818 5698 10824 5712
rect 10706 5632 10712 5646
rect 10818 5632 10824 5646
rect 10706 5566 10712 5580
rect 10818 5566 10824 5580
rect 10706 5499 10712 5514
rect 10818 5499 10824 5514
rect 10706 5432 10712 5447
rect 10818 5432 10824 5447
rect 10706 5368 10824 5380
rect 11035 14338 11049 14390
rect 11537 14720 11655 14726
rect 11589 14668 11603 14720
rect 11537 14654 11655 14668
rect 11589 14602 11603 14654
rect 11537 14588 11655 14602
rect 11589 14536 11603 14588
rect 11537 14522 11655 14536
rect 11589 14470 11603 14522
rect 11537 14456 11655 14470
rect 11589 14404 11603 14456
rect 11537 14390 11655 14404
rect 10983 14323 10989 14338
rect 11023 14323 11061 14338
rect 11095 14323 11101 14338
rect 11035 14271 11049 14323
rect 10983 14267 11101 14271
rect 10983 14256 10989 14267
rect 11023 14256 11061 14267
rect 11095 14256 11101 14267
rect 11035 14204 11049 14256
rect 10983 14189 11101 14204
rect 10983 14155 10989 14189
rect 11023 14155 11061 14189
rect 11095 14155 11101 14189
rect 10983 14111 11101 14155
rect 10983 14077 10989 14111
rect 11023 14077 11061 14111
rect 11095 14077 11101 14111
rect 10983 14033 11101 14077
rect 10983 13999 10989 14033
rect 11023 13999 11061 14033
rect 11095 13999 11101 14033
rect 10983 13955 11101 13999
rect 10983 13921 10989 13955
rect 11023 13921 11061 13955
rect 11095 13921 11101 13955
rect 10983 13877 11101 13921
rect 10983 13843 10989 13877
rect 11023 13843 11061 13877
rect 11095 13843 11101 13877
rect 10983 13799 11101 13843
rect 10983 13765 10989 13799
rect 11023 13765 11061 13799
rect 11095 13765 11101 13799
rect 10983 13722 11101 13765
rect 10983 13688 10989 13722
rect 11023 13688 11061 13722
rect 11095 13688 11101 13722
rect 10983 13645 11101 13688
rect 10983 13611 10989 13645
rect 11023 13611 11061 13645
rect 11095 13611 11101 13645
rect 10983 13568 11101 13611
rect 10983 13534 10989 13568
rect 11023 13534 11061 13568
rect 11095 13534 11101 13568
rect 10983 13491 11101 13534
rect 10983 13457 10989 13491
rect 11023 13457 11061 13491
rect 11095 13457 11101 13491
rect 10983 13414 11101 13457
rect 10983 13380 10989 13414
rect 11023 13380 11061 13414
rect 11095 13380 11101 13414
rect 10983 12720 11101 13380
rect 11035 12668 11049 12720
rect 10983 12654 11101 12668
rect 11035 12602 11049 12654
rect 10983 12588 11101 12602
rect 11035 12536 11049 12588
rect 10983 12534 10989 12536
rect 11023 12534 11061 12536
rect 11095 12534 11101 12536
rect 10983 12522 11101 12534
rect 11035 12470 11049 12522
rect 10983 12461 10989 12470
rect 11023 12461 11061 12470
rect 11095 12461 11101 12470
rect 10983 12456 11101 12461
rect 11035 12422 11049 12456
rect 10983 12390 10989 12404
rect 11095 12390 11101 12404
rect 10983 12323 10989 12338
rect 11095 12323 11101 12338
rect 10983 12256 10989 12271
rect 11095 12256 11101 12271
rect 10983 11380 10989 12204
rect 11095 11380 11101 12204
rect 10983 10724 11101 11380
rect 11035 10672 11049 10724
rect 10983 10658 11101 10672
rect 11035 10606 11049 10658
rect 10983 10592 11101 10606
rect 11035 10540 11049 10592
rect 10983 10534 10989 10540
rect 11023 10534 11061 10540
rect 11095 10534 11101 10540
rect 10983 10526 11101 10534
rect 11035 10474 11049 10526
rect 10983 10461 10989 10474
rect 11023 10461 11061 10474
rect 11095 10461 11101 10474
rect 10983 10460 11101 10461
rect 11035 10422 11049 10460
rect 10983 10394 10989 10408
rect 11095 10394 11101 10408
rect 10983 10327 10989 10342
rect 11095 10327 11101 10342
rect 10983 10260 10989 10275
rect 11095 10260 11101 10275
rect 10983 9380 10989 10208
rect 11095 9380 11101 10208
rect 10983 8720 11101 9380
rect 11035 8668 11049 8720
rect 10983 8654 11101 8668
rect 11035 8602 11049 8654
rect 10983 8588 11101 8602
rect 11035 8536 11049 8588
rect 10983 8534 10989 8536
rect 11023 8534 11061 8536
rect 11095 8534 11101 8536
rect 10983 8522 11101 8534
rect 11035 8470 11049 8522
rect 10983 8461 10989 8470
rect 11023 8461 11061 8470
rect 11095 8461 11101 8470
rect 10983 8456 11101 8461
rect 11035 8422 11049 8456
rect 10983 8390 10989 8404
rect 11095 8390 11101 8404
rect 10983 8323 10989 8338
rect 11095 8323 11101 8338
rect 10983 8256 10989 8271
rect 11095 8256 11101 8271
rect 10983 7380 10989 8204
rect 11095 7380 11101 8204
rect 10983 6724 11101 7380
rect 11035 6672 11049 6724
rect 10983 6658 11101 6672
rect 11035 6606 11049 6658
rect 10983 6592 11101 6606
rect 11035 6540 11049 6592
rect 10983 6534 10989 6540
rect 11023 6534 11061 6540
rect 11095 6534 11101 6540
rect 10983 6526 11101 6534
rect 11035 6474 11049 6526
rect 10983 6461 10989 6474
rect 11023 6461 11061 6474
rect 11095 6461 11101 6474
rect 10983 6460 11101 6461
rect 11035 6422 11049 6460
rect 10983 6394 10989 6408
rect 11095 6394 11101 6408
rect 10983 6327 10989 6342
rect 11095 6327 11101 6342
rect 10983 6260 10989 6275
rect 11095 6260 11101 6275
rect 10983 5380 10989 6208
rect 11095 5380 11101 6208
tri 10547 5265 10553 5271 sw
tri 10977 5265 10983 5271 se
rect 10983 5265 11101 5380
rect 11260 14345 11378 14357
rect 11260 14311 11266 14345
rect 11300 14311 11338 14345
rect 11372 14311 11378 14345
rect 11260 14267 11378 14311
rect 11260 14233 11266 14267
rect 11300 14233 11338 14267
rect 11372 14233 11378 14267
rect 11260 14189 11378 14233
rect 11260 14155 11266 14189
rect 11300 14155 11338 14189
rect 11372 14155 11378 14189
rect 11260 14111 11378 14155
rect 11260 14077 11266 14111
rect 11300 14077 11338 14111
rect 11372 14077 11378 14111
rect 11260 14033 11378 14077
rect 11260 13999 11266 14033
rect 11300 13999 11338 14033
rect 11372 13999 11378 14033
rect 11260 13955 11378 13999
rect 11260 13921 11266 13955
rect 11300 13921 11338 13955
rect 11372 13921 11378 13955
rect 11260 13892 11378 13921
rect 11312 13840 11326 13892
rect 11260 13826 11378 13840
rect 11312 13774 11326 13826
rect 11260 13765 11266 13774
rect 11300 13765 11338 13774
rect 11372 13765 11378 13774
rect 11260 13760 11378 13765
rect 11312 13708 11326 13760
rect 11260 13694 11266 13708
rect 11300 13694 11338 13708
rect 11372 13694 11378 13708
rect 11312 13642 11326 13694
rect 11260 13628 11266 13642
rect 11300 13628 11338 13642
rect 11372 13628 11378 13642
rect 11312 13576 11326 13628
rect 11260 13568 11378 13576
rect 11260 13562 11266 13568
rect 11300 13562 11338 13568
rect 11372 13562 11378 13568
rect 11312 13510 11326 13562
rect 11260 13495 11378 13510
rect 11312 13443 11326 13495
rect 11260 13428 11378 13443
rect 11312 13376 11326 13428
rect 11260 12714 11378 13376
rect 11260 12680 11266 12714
rect 11300 12680 11338 12714
rect 11372 12680 11378 12714
rect 11260 12641 11378 12680
rect 11260 12607 11266 12641
rect 11300 12607 11338 12641
rect 11372 12607 11378 12641
rect 11260 12568 11378 12607
rect 11260 12534 11266 12568
rect 11300 12534 11338 12568
rect 11372 12534 11378 12568
rect 11260 12495 11378 12534
rect 11260 12461 11266 12495
rect 11300 12461 11338 12495
rect 11372 12461 11378 12495
rect 11260 12422 11378 12461
rect 11260 11892 11266 12422
rect 11372 11892 11378 12422
rect 11260 11826 11266 11840
rect 11372 11826 11378 11840
rect 11260 11760 11266 11774
rect 11372 11760 11378 11774
rect 11260 11694 11266 11708
rect 11372 11694 11378 11708
rect 11260 11628 11266 11642
rect 11372 11628 11378 11642
rect 11260 11562 11266 11576
rect 11372 11562 11378 11576
rect 11260 11495 11266 11510
rect 11372 11495 11378 11510
rect 11260 11428 11266 11443
rect 11372 11428 11378 11443
rect 11312 11376 11326 11380
rect 11260 10714 11378 11376
rect 11260 10680 11266 10714
rect 11300 10680 11338 10714
rect 11372 10680 11378 10714
rect 11260 10641 11378 10680
rect 11260 10607 11266 10641
rect 11300 10607 11338 10641
rect 11372 10607 11378 10641
rect 11260 10568 11378 10607
rect 11260 10534 11266 10568
rect 11300 10534 11338 10568
rect 11372 10534 11378 10568
rect 11260 10495 11378 10534
rect 11260 10461 11266 10495
rect 11300 10461 11338 10495
rect 11372 10461 11378 10495
rect 11260 10422 11378 10461
rect 11260 9896 11266 10422
rect 11372 9896 11378 10422
rect 11260 9830 11266 9844
rect 11372 9830 11378 9844
rect 11260 9764 11266 9778
rect 11372 9764 11378 9778
rect 11260 9698 11266 9712
rect 11372 9698 11378 9712
rect 11260 9632 11266 9646
rect 11372 9632 11378 9646
rect 11260 9566 11266 9580
rect 11372 9566 11378 9580
rect 11260 9499 11266 9514
rect 11372 9499 11378 9514
rect 11260 9432 11266 9447
rect 11372 9432 11378 9447
rect 11260 8714 11378 9380
rect 11260 8680 11266 8714
rect 11300 8680 11338 8714
rect 11372 8680 11378 8714
rect 11260 8641 11378 8680
rect 11260 8607 11266 8641
rect 11300 8607 11338 8641
rect 11372 8607 11378 8641
rect 11260 8568 11378 8607
rect 11260 8534 11266 8568
rect 11300 8534 11338 8568
rect 11372 8534 11378 8568
rect 11260 8495 11378 8534
rect 11260 8461 11266 8495
rect 11300 8461 11338 8495
rect 11372 8461 11378 8495
rect 11260 8422 11378 8461
rect 11260 7892 11266 8422
rect 11372 7892 11378 8422
rect 11260 7826 11266 7840
rect 11372 7826 11378 7840
rect 11260 7760 11266 7774
rect 11372 7760 11378 7774
rect 11260 7694 11266 7708
rect 11372 7694 11378 7708
rect 11260 7628 11266 7642
rect 11372 7628 11378 7642
rect 11260 7562 11266 7576
rect 11372 7562 11378 7576
rect 11260 7495 11266 7510
rect 11372 7495 11378 7510
rect 11260 7428 11266 7443
rect 11372 7428 11378 7443
rect 11312 7376 11326 7380
rect 11260 6714 11378 7376
rect 11260 6680 11266 6714
rect 11300 6680 11338 6714
rect 11372 6680 11378 6714
rect 11260 6641 11378 6680
rect 11260 6607 11266 6641
rect 11300 6607 11338 6641
rect 11372 6607 11378 6641
rect 11260 6568 11378 6607
rect 11260 6534 11266 6568
rect 11300 6534 11338 6568
rect 11372 6534 11378 6568
rect 11260 6495 11378 6534
rect 11260 6461 11266 6495
rect 11300 6461 11338 6495
rect 11372 6461 11378 6495
rect 11260 6422 11378 6461
rect 11260 5896 11266 6422
rect 11372 5896 11378 6422
rect 11260 5830 11266 5844
rect 11372 5830 11378 5844
rect 11260 5764 11266 5778
rect 11372 5764 11378 5778
rect 11260 5698 11266 5712
rect 11372 5698 11378 5712
rect 11260 5632 11266 5646
rect 11372 5632 11378 5646
rect 11260 5566 11266 5580
rect 11372 5566 11378 5580
rect 11260 5499 11266 5514
rect 11372 5499 11378 5514
rect 11260 5432 11266 5447
rect 11372 5432 11378 5447
rect 11260 5368 11378 5380
rect 11589 14338 11603 14390
rect 12091 14720 12209 14726
rect 12143 14668 12157 14720
rect 12091 14654 12209 14668
rect 12143 14602 12157 14654
rect 12091 14588 12209 14602
rect 12143 14536 12157 14588
rect 12091 14522 12209 14536
rect 12143 14470 12157 14522
rect 12091 14456 12209 14470
rect 12143 14404 12157 14456
rect 12091 14390 12209 14404
rect 11537 14323 11543 14338
rect 11577 14323 11615 14338
rect 11649 14323 11655 14338
rect 11589 14271 11603 14323
rect 11537 14267 11655 14271
rect 11537 14256 11543 14267
rect 11577 14256 11615 14267
rect 11649 14256 11655 14267
rect 11589 14204 11603 14256
rect 11537 14189 11655 14204
rect 11537 14155 11543 14189
rect 11577 14155 11615 14189
rect 11649 14155 11655 14189
rect 11537 14111 11655 14155
rect 11537 14077 11543 14111
rect 11577 14077 11615 14111
rect 11649 14077 11655 14111
rect 11537 14033 11655 14077
rect 11537 13999 11543 14033
rect 11577 13999 11615 14033
rect 11649 13999 11655 14033
rect 11537 13955 11655 13999
rect 11537 13921 11543 13955
rect 11577 13921 11615 13955
rect 11649 13921 11655 13955
rect 11537 13877 11655 13921
rect 11537 13843 11543 13877
rect 11577 13843 11615 13877
rect 11649 13843 11655 13877
rect 11537 13799 11655 13843
rect 11537 13765 11543 13799
rect 11577 13765 11615 13799
rect 11649 13765 11655 13799
rect 11537 13722 11655 13765
rect 11537 13688 11543 13722
rect 11577 13688 11615 13722
rect 11649 13688 11655 13722
rect 11537 13645 11655 13688
rect 11537 13611 11543 13645
rect 11577 13611 11615 13645
rect 11649 13611 11655 13645
rect 11537 13568 11655 13611
rect 11537 13534 11543 13568
rect 11577 13534 11615 13568
rect 11649 13534 11655 13568
rect 11537 13491 11655 13534
rect 11537 13457 11543 13491
rect 11577 13457 11615 13491
rect 11649 13457 11655 13491
rect 11537 13414 11655 13457
rect 11537 13380 11543 13414
rect 11577 13380 11615 13414
rect 11649 13380 11655 13414
rect 11537 12720 11655 13380
rect 11589 12668 11603 12720
rect 11537 12654 11655 12668
rect 11589 12602 11603 12654
rect 11537 12588 11655 12602
rect 11589 12536 11603 12588
rect 11537 12534 11543 12536
rect 11577 12534 11615 12536
rect 11649 12534 11655 12536
rect 11537 12522 11655 12534
rect 11589 12470 11603 12522
rect 11537 12461 11543 12470
rect 11577 12461 11615 12470
rect 11649 12461 11655 12470
rect 11537 12456 11655 12461
rect 11589 12422 11603 12456
rect 11537 12390 11543 12404
rect 11649 12390 11655 12404
rect 11537 12323 11543 12338
rect 11649 12323 11655 12338
rect 11537 12256 11543 12271
rect 11649 12256 11655 12271
rect 11537 11380 11543 12204
rect 11649 11380 11655 12204
rect 11537 10724 11655 11380
rect 11589 10672 11603 10724
rect 11537 10658 11655 10672
rect 11589 10606 11603 10658
rect 11537 10592 11655 10606
rect 11589 10540 11603 10592
rect 11537 10534 11543 10540
rect 11577 10534 11615 10540
rect 11649 10534 11655 10540
rect 11537 10526 11655 10534
rect 11589 10474 11603 10526
rect 11537 10461 11543 10474
rect 11577 10461 11615 10474
rect 11649 10461 11655 10474
rect 11537 10460 11655 10461
rect 11589 10422 11603 10460
rect 11537 10394 11543 10408
rect 11649 10394 11655 10408
rect 11537 10327 11543 10342
rect 11649 10327 11655 10342
rect 11537 10260 11543 10275
rect 11649 10260 11655 10275
rect 11537 9380 11543 10208
rect 11649 9380 11655 10208
rect 11537 8720 11655 9380
rect 11589 8668 11603 8720
rect 11537 8654 11655 8668
rect 11589 8602 11603 8654
rect 11537 8588 11655 8602
rect 11589 8536 11603 8588
rect 11537 8534 11543 8536
rect 11577 8534 11615 8536
rect 11649 8534 11655 8536
rect 11537 8522 11655 8534
rect 11589 8470 11603 8522
rect 11537 8461 11543 8470
rect 11577 8461 11615 8470
rect 11649 8461 11655 8470
rect 11537 8456 11655 8461
rect 11589 8422 11603 8456
rect 11537 8390 11543 8404
rect 11649 8390 11655 8404
rect 11537 8323 11543 8338
rect 11649 8323 11655 8338
rect 11537 8256 11543 8271
rect 11649 8256 11655 8271
rect 11537 7380 11543 8204
rect 11649 7380 11655 8204
rect 11537 6724 11655 7380
rect 11589 6672 11603 6724
rect 11537 6658 11655 6672
rect 11589 6606 11603 6658
rect 11537 6592 11655 6606
rect 11589 6540 11603 6592
rect 11537 6534 11543 6540
rect 11577 6534 11615 6540
rect 11649 6534 11655 6540
rect 11537 6526 11655 6534
rect 11589 6474 11603 6526
rect 11537 6461 11543 6474
rect 11577 6461 11615 6474
rect 11649 6461 11655 6474
rect 11537 6460 11655 6461
rect 11589 6422 11603 6460
rect 11537 6394 11543 6408
rect 11649 6394 11655 6408
rect 11537 6327 11543 6342
rect 11649 6327 11655 6342
rect 11537 6260 11543 6275
rect 11649 6260 11655 6275
rect 11537 5380 11543 6208
rect 11649 5380 11655 6208
tri 11101 5265 11107 5271 sw
tri 11531 5265 11537 5271 se
rect 11537 5265 11655 5380
rect 11814 14345 11932 14357
rect 11814 14311 11820 14345
rect 11854 14311 11892 14345
rect 11926 14311 11932 14345
rect 11814 14267 11932 14311
rect 11814 14233 11820 14267
rect 11854 14233 11892 14267
rect 11926 14233 11932 14267
rect 11814 14189 11932 14233
rect 11814 14155 11820 14189
rect 11854 14155 11892 14189
rect 11926 14155 11932 14189
rect 11814 14111 11932 14155
rect 11814 14077 11820 14111
rect 11854 14077 11892 14111
rect 11926 14077 11932 14111
rect 11814 14033 11932 14077
rect 11814 13999 11820 14033
rect 11854 13999 11892 14033
rect 11926 13999 11932 14033
rect 11814 13955 11932 13999
rect 11814 13921 11820 13955
rect 11854 13921 11892 13955
rect 11926 13921 11932 13955
rect 11814 13892 11932 13921
rect 11866 13840 11880 13892
rect 11814 13826 11932 13840
rect 11866 13774 11880 13826
rect 11814 13765 11820 13774
rect 11854 13765 11892 13774
rect 11926 13765 11932 13774
rect 11814 13760 11932 13765
rect 11866 13708 11880 13760
rect 11814 13694 11820 13708
rect 11854 13694 11892 13708
rect 11926 13694 11932 13708
rect 11866 13642 11880 13694
rect 11814 13628 11820 13642
rect 11854 13628 11892 13642
rect 11926 13628 11932 13642
rect 11866 13576 11880 13628
rect 11814 13568 11932 13576
rect 11814 13562 11820 13568
rect 11854 13562 11892 13568
rect 11926 13562 11932 13568
rect 11866 13510 11880 13562
rect 11814 13495 11932 13510
rect 11866 13443 11880 13495
rect 11814 13428 11932 13443
rect 11866 13376 11880 13428
rect 11814 12714 11932 13376
rect 11814 12680 11820 12714
rect 11854 12680 11892 12714
rect 11926 12680 11932 12714
rect 11814 12641 11932 12680
rect 11814 12607 11820 12641
rect 11854 12607 11892 12641
rect 11926 12607 11932 12641
rect 11814 12568 11932 12607
rect 11814 12534 11820 12568
rect 11854 12534 11892 12568
rect 11926 12534 11932 12568
rect 11814 12495 11932 12534
rect 11814 12461 11820 12495
rect 11854 12461 11892 12495
rect 11926 12461 11932 12495
rect 11814 12422 11932 12461
rect 11814 11892 11820 12422
rect 11926 11892 11932 12422
rect 11814 11826 11820 11840
rect 11926 11826 11932 11840
rect 11814 11760 11820 11774
rect 11926 11760 11932 11774
rect 11814 11694 11820 11708
rect 11926 11694 11932 11708
rect 11814 11628 11820 11642
rect 11926 11628 11932 11642
rect 11814 11562 11820 11576
rect 11926 11562 11932 11576
rect 11814 11495 11820 11510
rect 11926 11495 11932 11510
rect 11814 11428 11820 11443
rect 11926 11428 11932 11443
rect 11866 11376 11880 11380
rect 11814 10714 11932 11376
rect 11814 10680 11820 10714
rect 11854 10680 11892 10714
rect 11926 10680 11932 10714
rect 11814 10641 11932 10680
rect 11814 10607 11820 10641
rect 11854 10607 11892 10641
rect 11926 10607 11932 10641
rect 11814 10568 11932 10607
rect 11814 10534 11820 10568
rect 11854 10534 11892 10568
rect 11926 10534 11932 10568
rect 11814 10495 11932 10534
rect 11814 10461 11820 10495
rect 11854 10461 11892 10495
rect 11926 10461 11932 10495
rect 11814 10422 11932 10461
rect 11814 9896 11820 10422
rect 11926 9896 11932 10422
rect 11814 9830 11820 9844
rect 11926 9830 11932 9844
rect 11814 9764 11820 9778
rect 11926 9764 11932 9778
rect 11814 9698 11820 9712
rect 11926 9698 11932 9712
rect 11814 9632 11820 9646
rect 11926 9632 11932 9646
rect 11814 9566 11820 9580
rect 11926 9566 11932 9580
rect 11814 9499 11820 9514
rect 11926 9499 11932 9514
rect 11814 9432 11820 9447
rect 11926 9432 11932 9447
rect 11814 8714 11932 9380
rect 11814 8680 11820 8714
rect 11854 8680 11892 8714
rect 11926 8680 11932 8714
rect 11814 8641 11932 8680
rect 11814 8607 11820 8641
rect 11854 8607 11892 8641
rect 11926 8607 11932 8641
rect 11814 8568 11932 8607
rect 11814 8534 11820 8568
rect 11854 8534 11892 8568
rect 11926 8534 11932 8568
rect 11814 8495 11932 8534
rect 11814 8461 11820 8495
rect 11854 8461 11892 8495
rect 11926 8461 11932 8495
rect 11814 8422 11932 8461
rect 11814 7892 11820 8422
rect 11926 7892 11932 8422
rect 11814 7826 11820 7840
rect 11926 7826 11932 7840
rect 11814 7760 11820 7774
rect 11926 7760 11932 7774
rect 11814 7694 11820 7708
rect 11926 7694 11932 7708
rect 11814 7628 11820 7642
rect 11926 7628 11932 7642
rect 11814 7562 11820 7576
rect 11926 7562 11932 7576
rect 11814 7495 11820 7510
rect 11926 7495 11932 7510
rect 11814 7428 11820 7443
rect 11926 7428 11932 7443
rect 11866 7376 11880 7380
rect 11814 6714 11932 7376
rect 11814 6680 11820 6714
rect 11854 6680 11892 6714
rect 11926 6680 11932 6714
rect 11814 6641 11932 6680
rect 11814 6607 11820 6641
rect 11854 6607 11892 6641
rect 11926 6607 11932 6641
rect 11814 6568 11932 6607
rect 11814 6534 11820 6568
rect 11854 6534 11892 6568
rect 11926 6534 11932 6568
rect 11814 6495 11932 6534
rect 11814 6461 11820 6495
rect 11854 6461 11892 6495
rect 11926 6461 11932 6495
rect 11814 6422 11932 6461
rect 11814 5896 11820 6422
rect 11926 5896 11932 6422
rect 11814 5830 11820 5844
rect 11926 5830 11932 5844
rect 11814 5764 11820 5778
rect 11926 5764 11932 5778
rect 11814 5698 11820 5712
rect 11926 5698 11932 5712
rect 11814 5632 11820 5646
rect 11926 5632 11932 5646
rect 11814 5566 11820 5580
rect 11926 5566 11932 5580
rect 11814 5499 11820 5514
rect 11926 5499 11932 5514
rect 11814 5432 11820 5447
rect 11926 5432 11932 5447
rect 11814 5368 11932 5380
rect 12143 14338 12157 14390
rect 12645 14720 12763 14726
rect 12697 14668 12711 14720
rect 12645 14654 12763 14668
rect 12697 14602 12711 14654
rect 12645 14588 12763 14602
rect 12697 14536 12711 14588
rect 12645 14522 12763 14536
rect 12697 14470 12711 14522
rect 12645 14456 12763 14470
rect 12697 14404 12711 14456
rect 12645 14390 12763 14404
rect 12091 14323 12097 14338
rect 12131 14323 12169 14338
rect 12203 14323 12209 14338
rect 12143 14271 12157 14323
rect 12091 14267 12209 14271
rect 12091 14256 12097 14267
rect 12131 14256 12169 14267
rect 12203 14256 12209 14267
rect 12143 14204 12157 14256
rect 12091 14189 12209 14204
rect 12091 14155 12097 14189
rect 12131 14155 12169 14189
rect 12203 14155 12209 14189
rect 12091 14111 12209 14155
rect 12091 14077 12097 14111
rect 12131 14077 12169 14111
rect 12203 14077 12209 14111
rect 12091 14033 12209 14077
rect 12091 13999 12097 14033
rect 12131 13999 12169 14033
rect 12203 13999 12209 14033
rect 12091 13955 12209 13999
rect 12091 13921 12097 13955
rect 12131 13921 12169 13955
rect 12203 13921 12209 13955
rect 12091 13877 12209 13921
rect 12091 13843 12097 13877
rect 12131 13843 12169 13877
rect 12203 13843 12209 13877
rect 12091 13799 12209 13843
rect 12091 13765 12097 13799
rect 12131 13765 12169 13799
rect 12203 13765 12209 13799
rect 12091 13722 12209 13765
rect 12091 13688 12097 13722
rect 12131 13688 12169 13722
rect 12203 13688 12209 13722
rect 12091 13645 12209 13688
rect 12091 13611 12097 13645
rect 12131 13611 12169 13645
rect 12203 13611 12209 13645
rect 12091 13568 12209 13611
rect 12091 13534 12097 13568
rect 12131 13534 12169 13568
rect 12203 13534 12209 13568
rect 12091 13491 12209 13534
rect 12091 13457 12097 13491
rect 12131 13457 12169 13491
rect 12203 13457 12209 13491
rect 12091 13414 12209 13457
rect 12091 13380 12097 13414
rect 12131 13380 12169 13414
rect 12203 13380 12209 13414
rect 12091 12720 12209 13380
rect 12143 12668 12157 12720
rect 12091 12654 12209 12668
rect 12143 12602 12157 12654
rect 12091 12588 12209 12602
rect 12143 12536 12157 12588
rect 12091 12534 12097 12536
rect 12131 12534 12169 12536
rect 12203 12534 12209 12536
rect 12091 12522 12209 12534
rect 12143 12470 12157 12522
rect 12091 12461 12097 12470
rect 12131 12461 12169 12470
rect 12203 12461 12209 12470
rect 12091 12456 12209 12461
rect 12143 12422 12157 12456
rect 12091 12390 12097 12404
rect 12203 12390 12209 12404
rect 12091 12323 12097 12338
rect 12203 12323 12209 12338
rect 12091 12256 12097 12271
rect 12203 12256 12209 12271
rect 12091 11380 12097 12204
rect 12203 11380 12209 12204
rect 12091 10724 12209 11380
rect 12143 10672 12157 10724
rect 12091 10658 12209 10672
rect 12143 10606 12157 10658
rect 12091 10592 12209 10606
rect 12143 10540 12157 10592
rect 12091 10534 12097 10540
rect 12131 10534 12169 10540
rect 12203 10534 12209 10540
rect 12091 10526 12209 10534
rect 12143 10474 12157 10526
rect 12091 10461 12097 10474
rect 12131 10461 12169 10474
rect 12203 10461 12209 10474
rect 12091 10460 12209 10461
rect 12143 10422 12157 10460
rect 12091 10394 12097 10408
rect 12203 10394 12209 10408
rect 12091 10327 12097 10342
rect 12203 10327 12209 10342
rect 12091 10260 12097 10275
rect 12203 10260 12209 10275
rect 12091 9380 12097 10208
rect 12203 9380 12209 10208
rect 12091 8720 12209 9380
rect 12143 8668 12157 8720
rect 12091 8654 12209 8668
rect 12143 8602 12157 8654
rect 12091 8588 12209 8602
rect 12143 8536 12157 8588
rect 12091 8534 12097 8536
rect 12131 8534 12169 8536
rect 12203 8534 12209 8536
rect 12091 8522 12209 8534
rect 12143 8470 12157 8522
rect 12091 8461 12097 8470
rect 12131 8461 12169 8470
rect 12203 8461 12209 8470
rect 12091 8456 12209 8461
rect 12143 8422 12157 8456
rect 12091 8390 12097 8404
rect 12203 8390 12209 8404
rect 12091 8323 12097 8338
rect 12203 8323 12209 8338
rect 12091 8256 12097 8271
rect 12203 8256 12209 8271
rect 12091 7380 12097 8204
rect 12203 7380 12209 8204
rect 12091 6724 12209 7380
rect 12143 6672 12157 6724
rect 12091 6658 12209 6672
rect 12143 6606 12157 6658
rect 12091 6592 12209 6606
rect 12143 6540 12157 6592
rect 12091 6534 12097 6540
rect 12131 6534 12169 6540
rect 12203 6534 12209 6540
rect 12091 6526 12209 6534
rect 12143 6474 12157 6526
rect 12091 6461 12097 6474
rect 12131 6461 12169 6474
rect 12203 6461 12209 6474
rect 12091 6460 12209 6461
rect 12143 6422 12157 6460
rect 12091 6394 12097 6408
rect 12203 6394 12209 6408
rect 12091 6327 12097 6342
rect 12203 6327 12209 6342
rect 12091 6260 12097 6275
rect 12203 6260 12209 6275
rect 12091 5380 12097 6208
rect 12203 5380 12209 6208
tri 11655 5265 11661 5271 sw
tri 12085 5265 12091 5271 se
rect 12091 5265 12209 5380
rect 12368 14345 12486 14357
rect 12368 14311 12374 14345
rect 12408 14311 12446 14345
rect 12480 14311 12486 14345
rect 12368 14267 12486 14311
rect 12368 14233 12374 14267
rect 12408 14233 12446 14267
rect 12480 14233 12486 14267
rect 12368 14189 12486 14233
rect 12368 14155 12374 14189
rect 12408 14155 12446 14189
rect 12480 14155 12486 14189
rect 12368 14111 12486 14155
rect 12368 14077 12374 14111
rect 12408 14077 12446 14111
rect 12480 14077 12486 14111
rect 12368 14033 12486 14077
rect 12368 13999 12374 14033
rect 12408 13999 12446 14033
rect 12480 13999 12486 14033
rect 12368 13955 12486 13999
rect 12368 13921 12374 13955
rect 12408 13921 12446 13955
rect 12480 13921 12486 13955
rect 12368 13892 12486 13921
rect 12420 13840 12434 13892
rect 12368 13826 12486 13840
rect 12420 13774 12434 13826
rect 12368 13765 12374 13774
rect 12408 13765 12446 13774
rect 12480 13765 12486 13774
rect 12368 13760 12486 13765
rect 12420 13708 12434 13760
rect 12368 13694 12374 13708
rect 12408 13694 12446 13708
rect 12480 13694 12486 13708
rect 12420 13642 12434 13694
rect 12368 13628 12374 13642
rect 12408 13628 12446 13642
rect 12480 13628 12486 13642
rect 12420 13576 12434 13628
rect 12368 13568 12486 13576
rect 12368 13562 12374 13568
rect 12408 13562 12446 13568
rect 12480 13562 12486 13568
rect 12420 13510 12434 13562
rect 12368 13495 12486 13510
rect 12420 13443 12434 13495
rect 12368 13428 12486 13443
rect 12420 13376 12434 13428
rect 12368 12714 12486 13376
rect 12368 12680 12374 12714
rect 12408 12680 12446 12714
rect 12480 12680 12486 12714
rect 12368 12641 12486 12680
rect 12368 12607 12374 12641
rect 12408 12607 12446 12641
rect 12480 12607 12486 12641
rect 12368 12568 12486 12607
rect 12368 12534 12374 12568
rect 12408 12534 12446 12568
rect 12480 12534 12486 12568
rect 12368 12495 12486 12534
rect 12368 12461 12374 12495
rect 12408 12461 12446 12495
rect 12480 12461 12486 12495
rect 12368 12422 12486 12461
rect 12368 11892 12374 12422
rect 12480 11892 12486 12422
rect 12368 11826 12374 11840
rect 12480 11826 12486 11840
rect 12368 11760 12374 11774
rect 12480 11760 12486 11774
rect 12368 11694 12374 11708
rect 12480 11694 12486 11708
rect 12368 11628 12374 11642
rect 12480 11628 12486 11642
rect 12368 11562 12374 11576
rect 12480 11562 12486 11576
rect 12368 11495 12374 11510
rect 12480 11495 12486 11510
rect 12368 11428 12374 11443
rect 12480 11428 12486 11443
rect 12420 11376 12434 11380
rect 12368 10714 12486 11376
rect 12368 10680 12374 10714
rect 12408 10680 12446 10714
rect 12480 10680 12486 10714
rect 12368 10641 12486 10680
rect 12368 10607 12374 10641
rect 12408 10607 12446 10641
rect 12480 10607 12486 10641
rect 12368 10568 12486 10607
rect 12368 10534 12374 10568
rect 12408 10534 12446 10568
rect 12480 10534 12486 10568
rect 12368 10495 12486 10534
rect 12368 10461 12374 10495
rect 12408 10461 12446 10495
rect 12480 10461 12486 10495
rect 12368 10422 12486 10461
rect 12368 9896 12374 10422
rect 12480 9896 12486 10422
rect 12368 9830 12374 9844
rect 12480 9830 12486 9844
rect 12368 9764 12374 9778
rect 12480 9764 12486 9778
rect 12368 9698 12374 9712
rect 12480 9698 12486 9712
rect 12368 9632 12374 9646
rect 12480 9632 12486 9646
rect 12368 9566 12374 9580
rect 12480 9566 12486 9580
rect 12368 9499 12374 9514
rect 12480 9499 12486 9514
rect 12368 9432 12374 9447
rect 12480 9432 12486 9447
rect 12368 8714 12486 9380
rect 12368 8680 12374 8714
rect 12408 8680 12446 8714
rect 12480 8680 12486 8714
rect 12368 8641 12486 8680
rect 12368 8607 12374 8641
rect 12408 8607 12446 8641
rect 12480 8607 12486 8641
rect 12368 8568 12486 8607
rect 12368 8534 12374 8568
rect 12408 8534 12446 8568
rect 12480 8534 12486 8568
rect 12368 8495 12486 8534
rect 12368 8461 12374 8495
rect 12408 8461 12446 8495
rect 12480 8461 12486 8495
rect 12368 8422 12486 8461
rect 12368 7891 12374 8422
rect 12480 7891 12486 8422
rect 12368 7825 12374 7839
rect 12480 7825 12486 7839
rect 12368 7759 12374 7773
rect 12480 7759 12486 7773
rect 12368 7693 12374 7707
rect 12480 7693 12486 7707
rect 12368 7627 12374 7641
rect 12480 7627 12486 7641
rect 12368 7561 12374 7575
rect 12480 7561 12486 7575
rect 12368 7494 12374 7509
rect 12480 7494 12486 7509
rect 12368 7427 12374 7442
rect 12480 7427 12486 7442
rect 12420 7375 12434 7380
rect 12368 6714 12486 7375
rect 12368 6680 12374 6714
rect 12408 6680 12446 6714
rect 12480 6680 12486 6714
rect 12368 6641 12486 6680
rect 12368 6607 12374 6641
rect 12408 6607 12446 6641
rect 12480 6607 12486 6641
rect 12368 6568 12486 6607
rect 12368 6534 12374 6568
rect 12408 6534 12446 6568
rect 12480 6534 12486 6568
rect 12368 6495 12486 6534
rect 12368 6461 12374 6495
rect 12408 6461 12446 6495
rect 12480 6461 12486 6495
rect 12368 6422 12486 6461
rect 12368 5894 12374 6422
rect 12480 5894 12486 6422
rect 12368 5828 12374 5842
rect 12480 5828 12486 5842
rect 12368 5762 12374 5776
rect 12480 5762 12486 5776
rect 12368 5696 12374 5710
rect 12480 5696 12486 5710
rect 12368 5630 12374 5644
rect 12480 5630 12486 5644
rect 12368 5564 12374 5578
rect 12480 5564 12486 5578
rect 12368 5497 12374 5512
rect 12480 5497 12486 5512
rect 12368 5430 12374 5445
rect 12480 5430 12486 5445
rect 12420 5378 12434 5380
rect 12368 5368 12486 5378
rect 12697 14338 12711 14390
rect 13199 14714 13490 14726
rect 13596 14714 13602 14726
rect 13199 14662 13200 14714
rect 13252 14662 13270 14714
rect 13322 14662 13340 14714
rect 13392 14662 13410 14714
rect 13462 14662 13480 14714
rect 13199 14650 13490 14662
rect 13596 14650 13602 14662
rect 13199 14598 13200 14650
rect 13252 14598 13270 14650
rect 13322 14598 13340 14650
rect 13392 14598 13410 14650
rect 13462 14598 13480 14650
rect 13199 14586 13490 14598
rect 13596 14586 13602 14598
rect 13199 14534 13200 14586
rect 13252 14534 13270 14586
rect 13322 14534 13340 14586
rect 13392 14534 13410 14586
rect 13462 14534 13480 14586
rect 13199 14522 13490 14534
rect 13596 14522 13602 14534
rect 13199 14470 13200 14522
rect 13252 14470 13270 14522
rect 13322 14470 13340 14522
rect 13392 14470 13410 14522
rect 13462 14470 13480 14522
rect 13199 14458 13490 14470
rect 13596 14458 13602 14470
rect 13199 14406 13200 14458
rect 13252 14406 13270 14458
rect 13322 14406 13340 14458
rect 13392 14406 13410 14458
rect 13462 14406 13480 14458
rect 13199 14394 13490 14406
rect 13596 14394 13602 14406
rect 12645 14323 12651 14338
rect 12685 14323 12723 14338
rect 12757 14323 12763 14338
rect 12697 14271 12711 14323
rect 12645 14267 12763 14271
rect 12645 14256 12651 14267
rect 12685 14256 12723 14267
rect 12757 14256 12763 14267
rect 12697 14204 12711 14256
rect 12645 14189 12763 14204
rect 12645 14155 12651 14189
rect 12685 14155 12723 14189
rect 12757 14155 12763 14189
rect 12645 14111 12763 14155
rect 12645 14077 12651 14111
rect 12685 14077 12723 14111
rect 12757 14077 12763 14111
rect 12645 14033 12763 14077
rect 12645 13999 12651 14033
rect 12685 13999 12723 14033
rect 12757 13999 12763 14033
rect 12645 13955 12763 13999
rect 12645 13921 12651 13955
rect 12685 13921 12723 13955
rect 12757 13921 12763 13955
rect 12645 13877 12763 13921
rect 12645 13843 12651 13877
rect 12685 13843 12723 13877
rect 12757 13843 12763 13877
rect 12645 13799 12763 13843
rect 12645 13765 12651 13799
rect 12685 13765 12723 13799
rect 12757 13765 12763 13799
rect 12645 13722 12763 13765
rect 12645 13688 12651 13722
rect 12685 13688 12723 13722
rect 12757 13688 12763 13722
rect 12645 13645 12763 13688
rect 12645 13611 12651 13645
rect 12685 13611 12723 13645
rect 12757 13611 12763 13645
rect 12645 13568 12763 13611
rect 12645 13534 12651 13568
rect 12685 13534 12723 13568
rect 12757 13534 12763 13568
rect 12645 13491 12763 13534
rect 12645 13457 12651 13491
rect 12685 13457 12723 13491
rect 12757 13457 12763 13491
rect 12645 13414 12763 13457
rect 12645 13380 12651 13414
rect 12685 13380 12723 13414
rect 12757 13380 12763 13414
rect 12645 12720 12763 13380
rect 12697 12668 12711 12720
rect 12645 12654 12763 12668
rect 12697 12602 12711 12654
rect 12645 12588 12763 12602
rect 12697 12536 12711 12588
rect 12645 12534 12651 12536
rect 12685 12534 12723 12536
rect 12757 12534 12763 12536
rect 12645 12522 12763 12534
rect 12697 12470 12711 12522
rect 12645 12461 12651 12470
rect 12685 12461 12723 12470
rect 12757 12461 12763 12470
rect 12645 12456 12763 12461
rect 12697 12422 12711 12456
rect 12645 12390 12651 12404
rect 12757 12390 12763 12404
rect 12645 12323 12651 12338
rect 12757 12323 12763 12338
rect 12645 12256 12651 12271
rect 12757 12256 12763 12271
rect 12645 11380 12651 12204
rect 12757 11380 12763 12204
rect 12645 10724 12763 11380
rect 12697 10672 12711 10724
rect 12645 10658 12763 10672
rect 12697 10606 12711 10658
rect 12645 10592 12763 10606
rect 12697 10540 12711 10592
rect 12645 10534 12651 10540
rect 12685 10534 12723 10540
rect 12757 10534 12763 10540
rect 12645 10526 12763 10534
rect 12697 10474 12711 10526
rect 12645 10461 12651 10474
rect 12685 10461 12723 10474
rect 12757 10461 12763 10474
rect 12645 10460 12763 10461
rect 12697 10422 12711 10460
rect 12645 10394 12651 10408
rect 12757 10394 12763 10408
rect 12645 10327 12651 10342
rect 12757 10327 12763 10342
rect 12645 10260 12651 10275
rect 12757 10260 12763 10275
rect 12645 9380 12651 10208
rect 12757 9380 12763 10208
rect 12645 8720 12763 9380
rect 12697 8668 12711 8720
rect 12645 8654 12763 8668
rect 12697 8602 12711 8654
rect 12645 8588 12763 8602
rect 12697 8536 12711 8588
rect 12645 8534 12651 8536
rect 12685 8534 12723 8536
rect 12757 8534 12763 8536
rect 12645 8522 12763 8534
rect 12697 8470 12711 8522
rect 12645 8461 12651 8470
rect 12685 8461 12723 8470
rect 12757 8461 12763 8470
rect 12645 8456 12763 8461
rect 12697 8422 12711 8456
rect 12645 8390 12651 8404
rect 12757 8390 12763 8404
rect 12645 8323 12651 8338
rect 12757 8323 12763 8338
rect 12645 8256 12651 8271
rect 12757 8256 12763 8271
rect 12645 7380 12651 8204
rect 12757 7380 12763 8204
rect 12645 6724 12763 7380
rect 12697 6672 12711 6724
rect 12645 6658 12763 6672
rect 12697 6606 12711 6658
rect 12645 6592 12763 6606
rect 12697 6540 12711 6592
rect 12645 6534 12651 6540
rect 12685 6534 12723 6540
rect 12757 6534 12763 6540
rect 12645 6526 12763 6534
rect 12697 6474 12711 6526
rect 12645 6461 12651 6474
rect 12685 6461 12723 6474
rect 12757 6461 12763 6474
rect 12645 6460 12763 6461
rect 12697 6422 12711 6460
rect 12645 6394 12651 6408
rect 12757 6394 12763 6408
rect 12645 6327 12651 6342
rect 12757 6327 12763 6342
rect 12645 6260 12651 6275
rect 12757 6260 12763 6275
rect 12645 5380 12651 6208
rect 12757 5380 12763 6208
tri 12209 5265 12215 5271 sw
tri 12639 5265 12645 5271 se
rect 12645 5265 12763 5380
rect 12922 14345 13040 14357
rect 12922 14311 12928 14345
rect 12962 14311 13000 14345
rect 13034 14311 13040 14345
rect 12922 14267 13040 14311
rect 12922 14233 12928 14267
rect 12962 14233 13000 14267
rect 13034 14233 13040 14267
rect 12922 14189 13040 14233
rect 12922 14155 12928 14189
rect 12962 14155 13000 14189
rect 13034 14155 13040 14189
rect 12922 14111 13040 14155
rect 12922 14077 12928 14111
rect 12962 14077 13000 14111
rect 13034 14077 13040 14111
rect 12922 14033 13040 14077
rect 12922 13999 12928 14033
rect 12962 13999 13000 14033
rect 13034 13999 13040 14033
rect 12922 13955 13040 13999
rect 12922 13921 12928 13955
rect 12962 13921 13000 13955
rect 13034 13921 13040 13955
rect 12922 13892 13040 13921
rect 12974 13840 12988 13892
rect 12922 13826 13040 13840
rect 12974 13774 12988 13826
rect 12922 13765 12928 13774
rect 12962 13765 13000 13774
rect 13034 13765 13040 13774
rect 12922 13760 13040 13765
rect 12974 13708 12988 13760
rect 12922 13694 12928 13708
rect 12962 13694 13000 13708
rect 13034 13694 13040 13708
rect 12974 13642 12988 13694
rect 12922 13628 12928 13642
rect 12962 13628 13000 13642
rect 13034 13628 13040 13642
rect 12974 13576 12988 13628
rect 12922 13568 13040 13576
rect 12922 13562 12928 13568
rect 12962 13562 13000 13568
rect 13034 13562 13040 13568
rect 12974 13510 12988 13562
rect 12922 13495 13040 13510
rect 12974 13443 12988 13495
rect 12922 13428 13040 13443
rect 12974 13376 12988 13428
rect 12922 12714 13040 13376
rect 12922 12680 12928 12714
rect 12962 12680 13000 12714
rect 13034 12680 13040 12714
rect 12922 12641 13040 12680
rect 12922 12607 12928 12641
rect 12962 12607 13000 12641
rect 13034 12607 13040 12641
rect 12922 12568 13040 12607
rect 12922 12534 12928 12568
rect 12962 12534 13000 12568
rect 13034 12534 13040 12568
rect 12922 12495 13040 12534
rect 12922 12461 12928 12495
rect 12962 12461 13000 12495
rect 13034 12461 13040 12495
rect 12922 12422 13040 12461
rect 12922 11892 12928 12422
rect 13034 11892 13040 12422
rect 12922 11826 12928 11840
rect 13034 11826 13040 11840
rect 12922 11760 12928 11774
rect 13034 11760 13040 11774
rect 12922 11694 12928 11708
rect 13034 11694 13040 11708
rect 12922 11628 12928 11642
rect 13034 11628 13040 11642
rect 12922 11562 12928 11576
rect 13034 11562 13040 11576
rect 12922 11495 12928 11510
rect 13034 11495 13040 11510
rect 12922 11428 12928 11443
rect 13034 11428 13040 11443
rect 12974 11376 12988 11380
rect 12922 10714 13040 11376
rect 12922 10680 12928 10714
rect 12962 10680 13000 10714
rect 13034 10680 13040 10714
rect 12922 10641 13040 10680
rect 12922 10607 12928 10641
rect 12962 10607 13000 10641
rect 13034 10607 13040 10641
rect 12922 10568 13040 10607
rect 12922 10534 12928 10568
rect 12962 10534 13000 10568
rect 13034 10534 13040 10568
rect 12922 10495 13040 10534
rect 12922 10461 12928 10495
rect 12962 10461 13000 10495
rect 13034 10461 13040 10495
rect 12922 10422 13040 10461
rect 12922 9896 12928 10422
rect 13034 9896 13040 10422
rect 12922 9830 12928 9844
rect 13034 9830 13040 9844
rect 12922 9764 12928 9778
rect 13034 9764 13040 9778
rect 12922 9698 12928 9712
rect 13034 9698 13040 9712
rect 12922 9632 12928 9646
rect 13034 9632 13040 9646
rect 12922 9566 12928 9580
rect 13034 9566 13040 9580
rect 12922 9499 12928 9514
rect 13034 9499 13040 9514
rect 12922 9432 12928 9447
rect 13034 9432 13040 9447
rect 12922 8714 13040 9380
rect 12922 8680 12928 8714
rect 12962 8680 13000 8714
rect 13034 8680 13040 8714
rect 12922 8641 13040 8680
rect 12922 8607 12928 8641
rect 12962 8607 13000 8641
rect 13034 8607 13040 8641
rect 12922 8568 13040 8607
rect 12922 8534 12928 8568
rect 12962 8534 13000 8568
rect 13034 8534 13040 8568
rect 12922 8495 13040 8534
rect 12922 8461 12928 8495
rect 12962 8461 13000 8495
rect 13034 8461 13040 8495
rect 12922 8422 13040 8461
rect 12922 7891 12928 8422
rect 13034 7891 13040 8422
rect 12922 7825 12928 7839
rect 13034 7825 13040 7839
rect 12922 7759 12928 7773
rect 13034 7759 13040 7773
rect 12922 7693 12928 7707
rect 13034 7693 13040 7707
rect 12922 7627 12928 7641
rect 13034 7627 13040 7641
rect 12922 7561 12928 7575
rect 13034 7561 13040 7575
rect 12922 7494 12928 7509
rect 13034 7494 13040 7509
rect 12922 7427 12928 7442
rect 13034 7427 13040 7442
rect 12974 7375 12988 7380
rect 12922 6714 13040 7375
rect 12922 6680 12928 6714
rect 12962 6680 13000 6714
rect 13034 6680 13040 6714
rect 12922 6641 13040 6680
rect 12922 6607 12928 6641
rect 12962 6607 13000 6641
rect 13034 6607 13040 6641
rect 12922 6568 13040 6607
rect 12922 6534 12928 6568
rect 12962 6534 13000 6568
rect 13034 6534 13040 6568
rect 12922 6495 13040 6534
rect 12922 6461 12928 6495
rect 12962 6461 13000 6495
rect 13034 6461 13040 6495
rect 12922 6422 13040 6461
rect 12922 5894 12928 6422
rect 13034 5894 13040 6422
rect 12922 5828 12928 5842
rect 13034 5828 13040 5842
rect 12922 5762 12928 5776
rect 13034 5762 13040 5776
rect 12922 5696 12928 5710
rect 13034 5696 13040 5710
rect 12922 5630 12928 5644
rect 13034 5630 13040 5644
rect 12922 5564 12928 5578
rect 13034 5564 13040 5578
rect 12922 5497 12928 5512
rect 13034 5497 13040 5512
rect 12922 5430 12928 5445
rect 13034 5430 13040 5445
rect 13199 14342 13200 14394
rect 13252 14342 13270 14394
rect 13322 14342 13340 14394
rect 13392 14342 13410 14394
rect 13462 14342 13480 14394
rect 13199 14330 13205 14342
rect 13239 14330 13277 14342
rect 13311 14330 13490 14342
rect 13596 14330 13602 14342
rect 13199 14278 13200 14330
rect 13252 14278 13270 14330
rect 13322 14278 13340 14330
rect 13392 14278 13410 14330
rect 13462 14278 13480 14330
rect 13199 14267 13490 14278
rect 13199 14266 13205 14267
rect 13239 14266 13277 14267
rect 13311 14266 13490 14267
rect 13596 14266 13602 14278
rect 13199 14214 13200 14266
rect 13252 14214 13270 14266
rect 13322 14214 13340 14266
rect 13392 14214 13410 14266
rect 13462 14214 13480 14266
rect 13199 14202 13490 14214
rect 13596 14202 13602 14214
rect 13199 14150 13200 14202
rect 13252 14150 13270 14202
rect 13322 14150 13340 14202
rect 13392 14150 13410 14202
rect 13462 14150 13480 14202
rect 13199 14138 13490 14150
rect 13596 14138 13602 14150
rect 13199 14086 13200 14138
rect 13252 14086 13270 14138
rect 13322 14086 13340 14138
rect 13392 14086 13410 14138
rect 13462 14086 13480 14138
rect 13199 14077 13205 14086
rect 13239 14077 13277 14086
rect 13311 14077 13490 14086
rect 13199 14074 13490 14077
rect 13596 14074 13602 14086
rect 13199 14022 13200 14074
rect 13252 14022 13270 14074
rect 13322 14022 13340 14074
rect 13392 14022 13410 14074
rect 13462 14022 13480 14074
rect 13199 14010 13205 14022
rect 13239 14010 13277 14022
rect 13311 14010 13490 14022
rect 13596 14010 13602 14022
rect 13199 13958 13200 14010
rect 13252 13958 13270 14010
rect 13322 13958 13340 14010
rect 13392 13958 13410 14010
rect 13462 13958 13480 14010
rect 13199 13955 13490 13958
rect 13199 13946 13205 13955
rect 13239 13946 13277 13955
rect 13311 13946 13490 13955
rect 13596 13946 13602 13958
rect 13199 13894 13200 13946
rect 13252 13894 13270 13946
rect 13322 13894 13340 13946
rect 13392 13894 13410 13946
rect 13462 13894 13480 13946
rect 13199 13882 13490 13894
rect 13596 13882 13602 13894
rect 13199 13830 13200 13882
rect 13252 13830 13270 13882
rect 13322 13830 13340 13882
rect 13392 13830 13410 13882
rect 13462 13830 13480 13882
rect 13199 13818 13490 13830
rect 13596 13818 13602 13830
rect 13199 13766 13200 13818
rect 13252 13766 13270 13818
rect 13322 13766 13340 13818
rect 13392 13766 13410 13818
rect 13462 13766 13480 13818
rect 13199 13765 13205 13766
rect 13239 13765 13277 13766
rect 13311 13765 13490 13766
rect 13199 13754 13490 13765
rect 13596 13754 13602 13766
rect 13199 13702 13200 13754
rect 13252 13702 13270 13754
rect 13322 13702 13340 13754
rect 13392 13702 13410 13754
rect 13462 13702 13480 13754
rect 13199 13690 13205 13702
rect 13239 13690 13277 13702
rect 13311 13690 13490 13702
rect 13596 13690 13602 13702
rect 13199 13638 13200 13690
rect 13252 13638 13270 13690
rect 13322 13638 13340 13690
rect 13392 13638 13410 13690
rect 13462 13638 13480 13690
rect 13199 13626 13205 13638
rect 13239 13626 13277 13638
rect 13311 13626 13490 13638
rect 13596 13626 13602 13638
rect 13199 13574 13200 13626
rect 13252 13574 13270 13626
rect 13322 13574 13340 13626
rect 13392 13574 13410 13626
rect 13462 13574 13480 13626
rect 13199 13568 13490 13574
rect 13199 13562 13205 13568
rect 13239 13562 13277 13568
rect 13311 13562 13490 13568
rect 13596 13562 13602 13574
rect 13199 13510 13200 13562
rect 13252 13510 13270 13562
rect 13322 13510 13340 13562
rect 13392 13510 13410 13562
rect 13462 13510 13480 13562
rect 13199 13498 13490 13510
rect 13596 13498 13602 13510
rect 13199 13446 13200 13498
rect 13252 13446 13270 13498
rect 13322 13446 13340 13498
rect 13392 13446 13410 13498
rect 13462 13446 13480 13498
rect 13199 13434 13490 13446
rect 13596 13434 13602 13446
rect 13199 13382 13200 13434
rect 13252 13382 13270 13434
rect 13322 13382 13340 13434
rect 13392 13382 13410 13434
rect 13462 13382 13480 13434
rect 13199 13380 13205 13382
rect 13239 13380 13277 13382
rect 13311 13380 13490 13382
rect 13199 13370 13490 13380
rect 13596 13370 13602 13382
rect 13199 13318 13200 13370
rect 13252 13318 13270 13370
rect 13322 13318 13340 13370
rect 13392 13318 13410 13370
rect 13462 13318 13480 13370
rect 13199 13306 13490 13318
rect 13596 13306 13602 13318
rect 13199 13254 13200 13306
rect 13252 13254 13270 13306
rect 13322 13254 13340 13306
rect 13392 13254 13410 13306
rect 13462 13254 13480 13306
rect 13199 13242 13490 13254
rect 13596 13242 13602 13254
rect 13199 13190 13200 13242
rect 13252 13190 13270 13242
rect 13322 13190 13340 13242
rect 13392 13190 13410 13242
rect 13462 13190 13480 13242
rect 13199 13178 13490 13190
rect 13596 13178 13602 13190
rect 13199 13126 13200 13178
rect 13252 13126 13270 13178
rect 13322 13126 13340 13178
rect 13392 13126 13410 13178
rect 13462 13126 13480 13178
rect 13199 13114 13490 13126
rect 13596 13114 13602 13126
rect 13199 13062 13200 13114
rect 13252 13062 13270 13114
rect 13322 13062 13340 13114
rect 13392 13062 13410 13114
rect 13462 13062 13480 13114
rect 13199 13050 13490 13062
rect 13596 13050 13602 13062
rect 13199 12998 13200 13050
rect 13252 12998 13270 13050
rect 13322 12998 13340 13050
rect 13392 12998 13410 13050
rect 13462 12998 13480 13050
rect 13199 12986 13490 12998
rect 13596 12986 13602 12998
rect 13199 12934 13200 12986
rect 13252 12934 13270 12986
rect 13322 12934 13340 12986
rect 13392 12934 13410 12986
rect 13462 12934 13480 12986
rect 13199 12922 13490 12934
rect 13596 12922 13602 12934
rect 13199 12870 13200 12922
rect 13252 12870 13270 12922
rect 13322 12870 13340 12922
rect 13392 12870 13410 12922
rect 13462 12870 13480 12922
rect 13199 12858 13490 12870
rect 13596 12858 13602 12870
rect 13199 12806 13200 12858
rect 13252 12806 13270 12858
rect 13322 12806 13340 12858
rect 13392 12806 13410 12858
rect 13462 12806 13480 12858
rect 13199 12794 13490 12806
rect 13596 12794 13602 12806
rect 13199 12742 13200 12794
rect 13252 12742 13270 12794
rect 13322 12742 13340 12794
rect 13392 12742 13410 12794
rect 13462 12742 13480 12794
rect 13199 12730 13490 12742
rect 13596 12730 13602 12742
rect 13199 12678 13200 12730
rect 13252 12678 13270 12730
rect 13322 12678 13340 12730
rect 13392 12678 13410 12730
rect 13462 12678 13480 12730
rect 13199 12666 13490 12678
rect 13596 12666 13602 12678
rect 13199 12614 13200 12666
rect 13252 12614 13270 12666
rect 13322 12614 13340 12666
rect 13392 12614 13410 12666
rect 13462 12614 13480 12666
rect 13199 12607 13205 12614
rect 13239 12607 13277 12614
rect 13311 12607 13490 12614
rect 13199 12602 13490 12607
rect 13596 12602 13602 12614
rect 13199 12550 13200 12602
rect 13252 12550 13270 12602
rect 13322 12550 13340 12602
rect 13392 12550 13410 12602
rect 13462 12550 13480 12602
rect 13199 12538 13205 12550
rect 13239 12538 13277 12550
rect 13311 12538 13490 12550
rect 13596 12538 13602 12550
rect 13199 12486 13200 12538
rect 13252 12486 13270 12538
rect 13322 12486 13340 12538
rect 13392 12486 13410 12538
rect 13462 12486 13480 12538
rect 13199 12474 13205 12486
rect 13239 12474 13277 12486
rect 13311 12474 13490 12486
rect 13596 12474 13602 12486
rect 13199 12422 13200 12474
rect 13252 12422 13270 12474
rect 13322 12422 13340 12474
rect 13392 12422 13410 12474
rect 13462 12422 13480 12474
rect 13199 12410 13205 12422
rect 13311 12410 13490 12422
rect 13596 12410 13602 12422
rect 13199 12358 13200 12410
rect 13322 12358 13340 12410
rect 13392 12358 13410 12410
rect 13462 12358 13480 12410
rect 13199 12346 13205 12358
rect 13311 12346 13490 12358
rect 13596 12346 13602 12358
rect 13199 12294 13200 12346
rect 13322 12294 13340 12346
rect 13392 12294 13410 12346
rect 13462 12294 13480 12346
rect 13199 12282 13205 12294
rect 13311 12282 13490 12294
rect 13596 12282 13602 12294
rect 13199 12230 13200 12282
rect 13322 12230 13340 12282
rect 13392 12230 13410 12282
rect 13462 12230 13480 12282
rect 13199 12218 13205 12230
rect 13311 12218 13490 12230
rect 13596 12218 13602 12230
rect 13199 12166 13200 12218
rect 13322 12166 13340 12218
rect 13392 12166 13410 12218
rect 13462 12166 13480 12218
rect 13199 12154 13205 12166
rect 13311 12154 13490 12166
rect 13596 12154 13602 12166
rect 13199 12102 13200 12154
rect 13322 12102 13340 12154
rect 13392 12102 13410 12154
rect 13462 12102 13480 12154
rect 13199 12090 13205 12102
rect 13311 12090 13490 12102
rect 13596 12090 13602 12102
rect 13199 12038 13200 12090
rect 13322 12038 13340 12090
rect 13392 12038 13410 12090
rect 13462 12038 13480 12090
rect 13199 12026 13205 12038
rect 13311 12026 13490 12038
rect 13596 12026 13602 12038
rect 13199 11974 13200 12026
rect 13322 11974 13340 12026
rect 13392 11974 13410 12026
rect 13462 11974 13480 12026
rect 13199 11962 13205 11974
rect 13311 11962 13490 11974
rect 13596 11962 13602 11974
rect 13199 11910 13200 11962
rect 13322 11910 13340 11962
rect 13392 11910 13410 11962
rect 13462 11910 13480 11962
rect 13199 11898 13205 11910
rect 13311 11898 13490 11910
rect 13596 11898 13602 11910
rect 13199 11846 13200 11898
rect 13322 11846 13340 11898
rect 13392 11846 13410 11898
rect 13462 11846 13480 11898
rect 13199 11834 13205 11846
rect 13311 11834 13490 11846
rect 13596 11834 13602 11846
rect 13199 11782 13200 11834
rect 13322 11782 13340 11834
rect 13392 11782 13410 11834
rect 13462 11782 13480 11834
rect 13199 11770 13205 11782
rect 13311 11770 13490 11782
rect 13596 11770 13602 11782
rect 13199 11718 13200 11770
rect 13322 11718 13340 11770
rect 13392 11718 13410 11770
rect 13462 11718 13480 11770
rect 13199 11706 13205 11718
rect 13311 11706 13490 11718
rect 13596 11706 13602 11718
rect 13199 11654 13200 11706
rect 13322 11654 13340 11706
rect 13392 11654 13410 11706
rect 13462 11654 13480 11706
rect 13199 11642 13205 11654
rect 13311 11642 13490 11654
rect 13596 11642 13602 11654
rect 13199 11590 13200 11642
rect 13322 11590 13340 11642
rect 13392 11590 13410 11642
rect 13462 11590 13480 11642
rect 13199 11578 13205 11590
rect 13311 11578 13490 11590
rect 13596 11578 13602 11590
rect 13199 11526 13200 11578
rect 13322 11526 13340 11578
rect 13392 11526 13410 11578
rect 13462 11526 13480 11578
rect 13199 11514 13205 11526
rect 13311 11514 13490 11526
rect 13596 11514 13602 11526
rect 13199 11462 13200 11514
rect 13322 11462 13340 11514
rect 13392 11462 13410 11514
rect 13462 11462 13480 11514
rect 13199 11450 13205 11462
rect 13311 11450 13490 11462
rect 13596 11450 13602 11462
rect 13199 11398 13200 11450
rect 13322 11398 13340 11450
rect 13392 11398 13410 11450
rect 13462 11398 13480 11450
rect 13199 11386 13205 11398
rect 13311 11386 13490 11398
rect 13596 11386 13602 11398
rect 13199 11334 13200 11386
rect 13252 11334 13270 11380
rect 13322 11334 13340 11386
rect 13392 11334 13410 11386
rect 13462 11334 13480 11386
rect 13199 11322 13490 11334
rect 13596 11322 13602 11334
rect 13199 11270 13200 11322
rect 13252 11270 13270 11322
rect 13322 11270 13340 11322
rect 13392 11270 13410 11322
rect 13462 11270 13480 11322
rect 13199 11258 13490 11270
rect 13596 11258 13602 11270
rect 13199 11206 13200 11258
rect 13252 11206 13270 11258
rect 13322 11206 13340 11258
rect 13392 11206 13410 11258
rect 13462 11206 13480 11258
rect 13199 11194 13490 11206
rect 13596 11194 13602 11206
rect 13199 11142 13200 11194
rect 13252 11142 13270 11194
rect 13322 11142 13340 11194
rect 13392 11142 13410 11194
rect 13462 11142 13480 11194
rect 13199 11130 13490 11142
rect 13596 11130 13602 11142
rect 13199 11078 13200 11130
rect 13252 11078 13270 11130
rect 13322 11078 13340 11130
rect 13392 11078 13410 11130
rect 13462 11078 13480 11130
rect 13199 11066 13490 11078
rect 13596 11066 13602 11078
rect 13199 11014 13200 11066
rect 13252 11014 13270 11066
rect 13322 11014 13340 11066
rect 13392 11014 13410 11066
rect 13462 11014 13480 11066
rect 13199 11002 13490 11014
rect 13596 11002 13602 11014
rect 13199 10950 13200 11002
rect 13252 10950 13270 11002
rect 13322 10950 13340 11002
rect 13392 10950 13410 11002
rect 13462 10950 13480 11002
rect 13199 10938 13490 10950
rect 13596 10938 13602 10950
rect 13199 10886 13200 10938
rect 13252 10886 13270 10938
rect 13322 10886 13340 10938
rect 13392 10886 13410 10938
rect 13462 10886 13480 10938
rect 13199 10874 13490 10886
rect 13596 10874 13602 10886
rect 13199 10822 13200 10874
rect 13252 10822 13270 10874
rect 13322 10822 13340 10874
rect 13392 10822 13410 10874
rect 13462 10822 13480 10874
rect 13199 10810 13490 10822
rect 13596 10810 13602 10822
rect 13199 10758 13200 10810
rect 13252 10758 13270 10810
rect 13322 10758 13340 10810
rect 13392 10758 13410 10810
rect 13462 10758 13480 10810
rect 13199 10746 13490 10758
rect 13596 10746 13602 10758
rect 13199 10694 13200 10746
rect 13252 10694 13270 10746
rect 13322 10694 13340 10746
rect 13392 10694 13410 10746
rect 13462 10694 13480 10746
rect 13199 10682 13205 10694
rect 13239 10682 13277 10694
rect 13311 10682 13490 10694
rect 13596 10682 13602 10694
rect 13199 10630 13200 10682
rect 13252 10630 13270 10682
rect 13322 10630 13340 10682
rect 13392 10630 13410 10682
rect 13462 10630 13480 10682
rect 13199 10618 13205 10630
rect 13239 10618 13277 10630
rect 13311 10618 13490 10630
rect 13596 10618 13602 10630
rect 13199 10566 13200 10618
rect 13252 10566 13270 10618
rect 13322 10566 13340 10618
rect 13392 10566 13410 10618
rect 13462 10566 13480 10618
rect 13199 10554 13205 10566
rect 13239 10554 13277 10566
rect 13311 10554 13490 10566
rect 13596 10554 13602 10566
rect 13199 10502 13200 10554
rect 13252 10502 13270 10554
rect 13322 10502 13340 10554
rect 13392 10502 13410 10554
rect 13462 10502 13480 10554
rect 13199 10495 13490 10502
rect 13199 10490 13205 10495
rect 13239 10490 13277 10495
rect 13311 10490 13490 10495
rect 13596 10490 13602 10502
rect 13199 10438 13200 10490
rect 13252 10438 13270 10490
rect 13322 10438 13340 10490
rect 13392 10438 13410 10490
rect 13462 10438 13480 10490
rect 13199 10426 13490 10438
rect 13596 10426 13602 10438
rect 13199 10374 13200 10426
rect 13252 10422 13270 10426
rect 13322 10374 13340 10426
rect 13392 10374 13410 10426
rect 13462 10374 13480 10426
rect 13199 10362 13205 10374
rect 13311 10362 13490 10374
rect 13596 10362 13602 10374
rect 13199 10310 13200 10362
rect 13322 10310 13340 10362
rect 13392 10310 13410 10362
rect 13462 10310 13480 10362
rect 13199 10298 13205 10310
rect 13311 10298 13490 10310
rect 13596 10298 13602 10310
rect 13199 10246 13200 10298
rect 13322 10246 13340 10298
rect 13392 10246 13410 10298
rect 13462 10246 13480 10298
rect 13199 10234 13205 10246
rect 13311 10234 13490 10246
rect 13596 10234 13602 10246
rect 13199 10182 13200 10234
rect 13322 10182 13340 10234
rect 13392 10182 13410 10234
rect 13462 10182 13480 10234
rect 13199 10170 13205 10182
rect 13311 10170 13490 10182
rect 13596 10170 13602 10182
rect 13199 10118 13200 10170
rect 13322 10118 13340 10170
rect 13392 10118 13410 10170
rect 13462 10118 13480 10170
rect 13199 10106 13205 10118
rect 13311 10106 13490 10118
rect 13596 10106 13602 10118
rect 13199 10054 13200 10106
rect 13322 10054 13340 10106
rect 13392 10054 13410 10106
rect 13462 10054 13480 10106
rect 13199 10042 13205 10054
rect 13311 10042 13490 10054
rect 13596 10042 13602 10054
rect 13199 9990 13200 10042
rect 13322 9990 13340 10042
rect 13392 9990 13410 10042
rect 13462 9990 13480 10042
rect 13199 9978 13205 9990
rect 13311 9978 13490 9990
rect 13596 9978 13602 9990
rect 13199 9926 13200 9978
rect 13322 9926 13340 9978
rect 13392 9926 13410 9978
rect 13462 9926 13480 9978
rect 13199 9914 13205 9926
rect 13311 9914 13490 9926
rect 13596 9914 13602 9926
rect 13199 9862 13200 9914
rect 13322 9862 13340 9914
rect 13392 9862 13410 9914
rect 13462 9862 13480 9914
rect 13199 9850 13205 9862
rect 13311 9850 13490 9862
rect 13596 9850 13602 9862
rect 13199 9798 13200 9850
rect 13322 9798 13340 9850
rect 13392 9798 13410 9850
rect 13462 9798 13480 9850
rect 13199 9786 13205 9798
rect 13311 9786 13490 9798
rect 13596 9786 13602 9798
rect 13199 9734 13200 9786
rect 13322 9734 13340 9786
rect 13392 9734 13410 9786
rect 13462 9734 13480 9786
rect 13199 9722 13205 9734
rect 13311 9722 13490 9734
rect 13596 9722 13602 9734
rect 13199 9670 13200 9722
rect 13322 9670 13340 9722
rect 13392 9670 13410 9722
rect 13462 9670 13480 9722
rect 13199 9658 13205 9670
rect 13311 9658 13490 9670
rect 13596 9658 13602 9670
rect 13199 9606 13200 9658
rect 13322 9606 13340 9658
rect 13392 9606 13410 9658
rect 13462 9606 13480 9658
rect 13199 9594 13205 9606
rect 13311 9594 13490 9606
rect 13596 9594 13602 9606
rect 13199 9542 13200 9594
rect 13322 9542 13340 9594
rect 13392 9542 13410 9594
rect 13462 9542 13480 9594
rect 13199 9530 13205 9542
rect 13311 9530 13490 9542
rect 13596 9530 13602 9542
rect 13199 9478 13200 9530
rect 13322 9478 13340 9530
rect 13392 9478 13410 9530
rect 13462 9478 13480 9530
rect 13199 9466 13205 9478
rect 13311 9466 13490 9478
rect 13596 9466 13602 9478
rect 13199 9414 13200 9466
rect 13322 9414 13340 9466
rect 13392 9414 13410 9466
rect 13462 9414 13480 9466
rect 13199 9402 13205 9414
rect 13311 9402 13490 9414
rect 13596 9402 13602 9414
rect 13199 9350 13200 9402
rect 13252 9350 13270 9380
rect 13322 9350 13340 9402
rect 13392 9350 13410 9402
rect 13462 9350 13480 9402
rect 13199 9338 13490 9350
rect 13596 9338 13602 9350
rect 13199 9286 13200 9338
rect 13252 9286 13270 9338
rect 13322 9286 13340 9338
rect 13392 9286 13410 9338
rect 13462 9286 13480 9338
rect 13199 9274 13490 9286
rect 13596 9274 13602 9286
rect 13199 9222 13200 9274
rect 13252 9222 13270 9274
rect 13322 9222 13340 9274
rect 13392 9222 13410 9274
rect 13462 9222 13480 9274
rect 13199 9210 13490 9222
rect 13596 9210 13602 9222
rect 13199 9158 13200 9210
rect 13252 9158 13270 9210
rect 13322 9158 13340 9210
rect 13392 9158 13410 9210
rect 13462 9158 13480 9210
rect 13199 9146 13490 9158
rect 13596 9146 13602 9158
rect 13199 9094 13200 9146
rect 13252 9094 13270 9146
rect 13322 9094 13340 9146
rect 13392 9094 13410 9146
rect 13462 9094 13480 9146
rect 13199 9082 13490 9094
rect 13596 9082 13602 9094
rect 13199 9030 13200 9082
rect 13252 9030 13270 9082
rect 13322 9030 13340 9082
rect 13392 9030 13410 9082
rect 13462 9030 13480 9082
rect 13199 9018 13490 9030
rect 13596 9018 13602 9030
rect 13199 8966 13200 9018
rect 13252 8966 13270 9018
rect 13322 8966 13340 9018
rect 13392 8966 13410 9018
rect 13462 8966 13480 9018
rect 13199 8954 13490 8966
rect 13596 8954 13602 8966
rect 13199 8902 13200 8954
rect 13252 8902 13270 8954
rect 13322 8902 13340 8954
rect 13392 8902 13410 8954
rect 13462 8902 13480 8954
rect 13199 8890 13490 8902
rect 13596 8890 13602 8902
rect 13199 8838 13200 8890
rect 13252 8838 13270 8890
rect 13322 8838 13340 8890
rect 13392 8838 13410 8890
rect 13462 8838 13480 8890
rect 13199 8826 13490 8838
rect 13596 8826 13602 8838
rect 13199 8774 13200 8826
rect 13252 8774 13270 8826
rect 13322 8774 13340 8826
rect 13392 8774 13410 8826
rect 13462 8774 13480 8826
rect 13199 8762 13490 8774
rect 13596 8762 13602 8774
rect 13199 8710 13200 8762
rect 13252 8710 13270 8762
rect 13322 8710 13340 8762
rect 13392 8710 13410 8762
rect 13462 8710 13480 8762
rect 13199 8698 13205 8710
rect 13239 8698 13277 8710
rect 13311 8698 13490 8710
rect 13596 8698 13602 8710
rect 13199 8646 13200 8698
rect 13252 8646 13270 8698
rect 13322 8646 13340 8698
rect 13392 8646 13410 8698
rect 13462 8646 13480 8698
rect 13199 8641 13490 8646
rect 13199 8634 13205 8641
rect 13239 8634 13277 8641
rect 13311 8634 13490 8641
rect 13596 8634 13602 8646
rect 13199 8582 13200 8634
rect 13252 8582 13270 8634
rect 13322 8582 13340 8634
rect 13392 8582 13410 8634
rect 13462 8582 13480 8634
rect 13199 8570 13490 8582
rect 13596 8570 13602 8582
rect 13199 8518 13200 8570
rect 13252 8518 13270 8570
rect 13322 8518 13340 8570
rect 13392 8518 13410 8570
rect 13462 8518 13480 8570
rect 13199 8506 13490 8518
rect 13596 8506 13602 8518
rect 13199 8454 13200 8506
rect 13252 8454 13270 8506
rect 13322 8454 13340 8506
rect 13392 8454 13410 8506
rect 13462 8454 13480 8506
rect 13199 8442 13490 8454
rect 13596 8442 13602 8454
rect 13199 8390 13200 8442
rect 13252 8422 13270 8442
rect 13322 8390 13340 8442
rect 13392 8390 13410 8442
rect 13462 8390 13480 8442
rect 13199 8378 13205 8390
rect 13311 8378 13490 8390
rect 13596 8378 13602 8390
rect 13199 8326 13200 8378
rect 13322 8326 13340 8378
rect 13392 8326 13410 8378
rect 13462 8326 13480 8378
rect 13199 8314 13205 8326
rect 13311 8314 13490 8326
rect 13596 8314 13602 8326
rect 13199 8262 13200 8314
rect 13322 8262 13340 8314
rect 13392 8262 13410 8314
rect 13462 8262 13480 8314
rect 13199 8250 13205 8262
rect 13311 8250 13490 8262
rect 13596 8250 13602 8262
rect 13199 8198 13200 8250
rect 13322 8198 13340 8250
rect 13392 8198 13410 8250
rect 13462 8198 13480 8250
rect 13199 8186 13205 8198
rect 13311 8186 13490 8198
rect 13596 8186 13602 8198
rect 13199 8134 13200 8186
rect 13322 8134 13340 8186
rect 13392 8134 13410 8186
rect 13462 8134 13480 8186
rect 13199 8122 13205 8134
rect 13311 8122 13490 8134
rect 13596 8122 13602 8134
rect 13199 8070 13200 8122
rect 13322 8070 13340 8122
rect 13392 8070 13410 8122
rect 13462 8070 13480 8122
rect 13199 8058 13205 8070
rect 13311 8058 13490 8070
rect 13596 8058 13602 8070
rect 13199 8006 13200 8058
rect 13322 8006 13340 8058
rect 13392 8006 13410 8058
rect 13462 8006 13480 8058
rect 13199 7994 13205 8006
rect 13311 7994 13490 8006
rect 13596 7994 13602 8006
rect 13199 7942 13200 7994
rect 13322 7942 13340 7994
rect 13392 7942 13410 7994
rect 13462 7942 13480 7994
rect 13199 7930 13205 7942
rect 13311 7930 13490 7942
rect 13596 7930 13602 7942
rect 13199 7878 13200 7930
rect 13322 7878 13340 7930
rect 13392 7878 13410 7930
rect 13462 7878 13480 7930
rect 13199 7866 13205 7878
rect 13311 7866 13490 7878
rect 13596 7866 13602 7878
rect 13199 7814 13200 7866
rect 13322 7814 13340 7866
rect 13392 7814 13410 7866
rect 13462 7814 13480 7866
rect 13199 7802 13205 7814
rect 13311 7802 13490 7814
rect 13596 7802 13602 7814
rect 13199 7750 13200 7802
rect 13322 7750 13340 7802
rect 13392 7750 13410 7802
rect 13462 7750 13480 7802
rect 13199 7738 13205 7750
rect 13311 7738 13490 7750
rect 13596 7738 13602 7750
rect 13199 7686 13200 7738
rect 13322 7686 13340 7738
rect 13392 7686 13410 7738
rect 13462 7686 13480 7738
rect 13199 7674 13205 7686
rect 13311 7674 13490 7686
rect 13596 7674 13602 7686
rect 13199 7622 13200 7674
rect 13322 7622 13340 7674
rect 13392 7622 13410 7674
rect 13462 7622 13480 7674
rect 13199 7610 13205 7622
rect 13311 7610 13490 7622
rect 13596 7610 13602 7622
rect 13199 7558 13200 7610
rect 13322 7558 13340 7610
rect 13392 7558 13410 7610
rect 13462 7558 13480 7610
rect 13199 7546 13205 7558
rect 13311 7546 13490 7558
rect 13596 7546 13602 7558
rect 13199 7494 13200 7546
rect 13322 7494 13340 7546
rect 13392 7494 13410 7546
rect 13462 7494 13480 7546
rect 13199 7482 13205 7494
rect 13311 7482 13490 7494
rect 13596 7482 13602 7494
rect 13199 7430 13200 7482
rect 13322 7430 13340 7482
rect 13392 7430 13410 7482
rect 13462 7430 13480 7482
rect 13199 7418 13205 7430
rect 13311 7418 13490 7430
rect 13596 7418 13602 7430
rect 13199 7366 13200 7418
rect 13252 7366 13270 7380
rect 13322 7366 13340 7418
rect 13392 7366 13410 7418
rect 13462 7366 13480 7418
rect 13199 7354 13490 7366
rect 13596 7354 13602 7366
rect 13199 7302 13200 7354
rect 13252 7302 13270 7354
rect 13322 7302 13340 7354
rect 13392 7302 13410 7354
rect 13462 7302 13480 7354
rect 13199 7290 13490 7302
rect 13596 7290 13602 7302
rect 13199 7238 13200 7290
rect 13252 7238 13270 7290
rect 13322 7238 13340 7290
rect 13392 7238 13410 7290
rect 13462 7238 13480 7290
rect 13199 7226 13490 7238
rect 13596 7226 13602 7238
rect 13199 7174 13200 7226
rect 13252 7174 13270 7226
rect 13322 7174 13340 7226
rect 13392 7174 13410 7226
rect 13462 7174 13480 7226
rect 13199 7162 13490 7174
rect 13596 7162 13602 7174
rect 13199 7110 13200 7162
rect 13252 7110 13270 7162
rect 13322 7110 13340 7162
rect 13392 7110 13410 7162
rect 13462 7110 13480 7162
tri 13799 7117 13832 7150 se
rect 13832 7117 13838 21329
rect 13199 7098 13490 7110
rect 13596 7098 13602 7110
rect 13199 7046 13200 7098
rect 13252 7046 13270 7098
rect 13322 7046 13340 7098
rect 13392 7046 13410 7098
rect 13462 7046 13480 7098
rect 13780 7071 13838 7117
rect 13199 7034 13490 7046
rect 13596 7034 13602 7046
tri 13799 7038 13832 7071 ne
rect 13199 6982 13200 7034
rect 13252 6982 13270 7034
rect 13322 6982 13340 7034
rect 13392 6982 13410 7034
rect 13462 6982 13480 7034
rect 13199 6970 13490 6982
rect 13596 6970 13602 6982
rect 13199 6918 13200 6970
rect 13252 6918 13270 6970
rect 13322 6918 13340 6970
rect 13392 6918 13410 6970
rect 13462 6918 13480 6970
rect 13199 6906 13490 6918
rect 13596 6906 13602 6918
rect 13199 6854 13200 6906
rect 13252 6854 13270 6906
rect 13322 6854 13340 6906
rect 13392 6854 13410 6906
rect 13462 6854 13480 6906
rect 13199 6842 13490 6854
rect 13596 6842 13602 6854
rect 13199 6790 13200 6842
rect 13252 6790 13270 6842
rect 13322 6790 13340 6842
rect 13392 6790 13410 6842
rect 13462 6790 13480 6842
rect 13199 6778 13490 6790
rect 13596 6778 13602 6790
rect 13199 6726 13200 6778
rect 13252 6726 13270 6778
rect 13322 6726 13340 6778
rect 13392 6726 13410 6778
rect 13462 6726 13480 6778
rect 13199 6714 13490 6726
rect 13596 6714 13602 6726
rect 13199 6662 13200 6714
rect 13252 6662 13270 6714
rect 13322 6662 13340 6714
rect 13392 6662 13410 6714
rect 13462 6662 13480 6714
rect 13199 6650 13490 6662
rect 13596 6650 13602 6662
rect 13199 6598 13200 6650
rect 13252 6598 13270 6650
rect 13322 6598 13340 6650
rect 13392 6598 13410 6650
rect 13462 6598 13480 6650
rect 13199 6586 13490 6598
rect 13596 6586 13602 6598
rect 13199 6534 13200 6586
rect 13252 6534 13270 6586
rect 13322 6534 13340 6586
rect 13392 6534 13410 6586
rect 13462 6534 13480 6586
rect 13199 6522 13490 6534
rect 13596 6522 13602 6534
rect 13199 6470 13200 6522
rect 13252 6470 13270 6522
rect 13322 6470 13340 6522
rect 13392 6470 13410 6522
rect 13462 6470 13480 6522
rect 13199 6461 13205 6470
rect 13239 6461 13277 6470
rect 13311 6461 13490 6470
rect 13199 6458 13490 6461
rect 13596 6458 13602 6470
rect 13199 6406 13200 6458
rect 13252 6422 13270 6458
rect 13322 6406 13340 6458
rect 13392 6406 13410 6458
rect 13462 6406 13480 6458
rect 13199 6394 13205 6406
rect 13311 6394 13490 6406
rect 13596 6394 13602 6406
rect 13199 6342 13200 6394
rect 13322 6342 13340 6394
rect 13392 6342 13410 6394
rect 13462 6342 13480 6394
rect 13199 6330 13205 6342
rect 13311 6330 13490 6342
rect 13596 6330 13602 6342
rect 13199 6278 13200 6330
rect 13322 6278 13340 6330
rect 13392 6278 13410 6330
rect 13462 6278 13480 6330
rect 13199 6266 13205 6278
rect 13311 6266 13490 6278
rect 13596 6266 13602 6278
rect 13199 6214 13200 6266
rect 13322 6214 13340 6266
rect 13392 6214 13410 6266
rect 13462 6214 13480 6266
rect 13199 6202 13205 6214
rect 13311 6202 13490 6214
rect 13596 6202 13602 6214
rect 13199 6150 13200 6202
rect 13322 6150 13340 6202
rect 13392 6150 13410 6202
rect 13462 6150 13480 6202
rect 13199 6138 13205 6150
rect 13311 6138 13490 6150
rect 13596 6138 13602 6150
rect 13199 6086 13200 6138
rect 13322 6086 13340 6138
rect 13392 6086 13410 6138
rect 13462 6086 13480 6138
rect 13199 6074 13205 6086
rect 13311 6074 13490 6086
rect 13596 6074 13602 6086
rect 13199 6022 13200 6074
rect 13322 6022 13340 6074
rect 13392 6022 13410 6074
rect 13462 6022 13480 6074
rect 13199 6010 13205 6022
rect 13311 6010 13490 6022
rect 13596 6010 13602 6022
rect 13199 5958 13200 6010
rect 13322 5958 13340 6010
rect 13392 5958 13410 6010
rect 13462 5958 13480 6010
rect 13199 5946 13205 5958
rect 13311 5946 13490 5958
rect 13596 5946 13602 5958
rect 13199 5894 13200 5946
rect 13322 5894 13340 5946
rect 13392 5894 13410 5946
rect 13462 5894 13480 5946
rect 13199 5882 13205 5894
rect 13311 5882 13490 5894
rect 13596 5882 13602 5894
rect 13199 5830 13200 5882
rect 13322 5830 13340 5882
rect 13392 5830 13410 5882
rect 13462 5830 13480 5882
rect 13199 5818 13205 5830
rect 13311 5818 13490 5830
rect 13596 5818 13602 5830
rect 13199 5766 13200 5818
rect 13322 5766 13340 5818
rect 13392 5766 13410 5818
rect 13462 5766 13480 5818
rect 13532 5766 13550 5815
rect 13199 5754 13205 5766
rect 13311 5754 13490 5766
rect 13524 5754 13562 5766
rect 13596 5754 13602 5766
rect 13199 5702 13200 5754
rect 13322 5702 13340 5754
rect 13392 5702 13410 5754
rect 13462 5702 13480 5754
rect 13532 5702 13550 5754
rect 13199 5690 13205 5702
rect 13311 5690 13490 5702
rect 13524 5690 13562 5702
rect 13596 5690 13602 5702
rect 13199 5638 13200 5690
rect 13322 5638 13340 5690
rect 13392 5638 13410 5690
rect 13462 5638 13480 5690
rect 13532 5638 13550 5690
rect 13199 5626 13205 5638
rect 13311 5630 13602 5638
rect 13311 5626 13490 5630
rect 13524 5626 13562 5630
rect 13596 5626 13602 5630
rect 13199 5574 13200 5626
rect 13322 5574 13340 5626
rect 13392 5574 13410 5626
rect 13462 5574 13480 5626
rect 13532 5574 13550 5626
rect 13199 5562 13205 5574
rect 13311 5562 13602 5574
rect 13199 5510 13200 5562
rect 13322 5510 13340 5562
rect 13392 5510 13410 5562
rect 13462 5510 13480 5562
rect 13532 5510 13550 5562
rect 13199 5498 13205 5510
rect 13311 5498 13602 5510
rect 13199 5446 13200 5498
rect 13322 5446 13340 5498
rect 13392 5446 13410 5498
rect 13462 5446 13480 5498
rect 13532 5446 13550 5498
rect 13199 5434 13205 5446
rect 13311 5434 13602 5446
tri 13162 5380 13199 5417 se
rect 13199 5382 13200 5434
rect 13322 5382 13340 5434
rect 13392 5382 13410 5434
rect 13462 5382 13480 5434
rect 13532 5382 13550 5434
rect 13199 5380 13205 5382
rect 13311 5380 13490 5382
rect 12974 5378 12988 5380
rect 12922 5368 13040 5378
tri 13159 5377 13162 5380 se
rect 13162 5377 13490 5380
rect 13524 5377 13562 5382
rect 13596 5377 13602 5382
tri 13154 5372 13159 5377 se
rect 13159 5372 13602 5377
tri 13150 5368 13154 5372 se
rect 13154 5370 13602 5372
rect 13154 5368 13200 5370
tri 13144 5362 13150 5368 se
rect 13150 5362 13200 5368
tri 13120 5338 13144 5362 se
rect 13144 5338 13200 5362
tri 13086 5304 13120 5338 se
rect 13120 5318 13200 5338
rect 13252 5318 13270 5370
rect 13322 5318 13340 5370
rect 13392 5318 13410 5370
rect 13462 5318 13480 5370
rect 13532 5318 13550 5370
rect 13120 5306 13490 5318
rect 13524 5306 13562 5318
rect 13596 5306 13602 5318
rect 13120 5304 13200 5306
tri 13071 5289 13086 5304 se
rect 13086 5289 13200 5304
tri 13053 5271 13071 5289 se
rect 13071 5271 13200 5289
tri 12763 5265 12769 5271 sw
tri 13047 5265 13053 5271 se
rect 13053 5265 13200 5271
rect 2361 5240 2973 5265
rect 2249 5237 2973 5240
tri 2973 5237 3001 5265 sw
tri 3193 5237 3221 5265 se
rect 3221 5237 3351 5265
tri 3351 5237 3379 5265 sw
tri 3747 5237 3775 5265 se
rect 3775 5237 3905 5265
tri 3905 5237 3933 5265 sw
tri 4301 5237 4329 5265 se
rect 4329 5237 4459 5265
tri 4459 5237 4487 5265 sw
tri 4855 5237 4883 5265 se
rect 4883 5237 5013 5265
tri 5013 5237 5041 5265 sw
tri 5409 5237 5437 5265 se
rect 5437 5237 5567 5265
tri 5567 5237 5595 5265 sw
tri 5963 5237 5991 5265 se
rect 5991 5237 6121 5265
tri 6121 5237 6149 5265 sw
tri 6517 5237 6545 5265 se
rect 6545 5237 6675 5265
tri 6675 5237 6703 5265 sw
tri 7071 5237 7099 5265 se
rect 7099 5237 7229 5265
tri 7229 5237 7257 5265 sw
tri 7625 5237 7653 5265 se
rect 7653 5237 7783 5265
tri 7783 5237 7811 5265 sw
tri 8179 5237 8207 5265 se
rect 8207 5237 8337 5265
tri 8337 5237 8365 5265 sw
tri 8733 5237 8761 5265 se
rect 8761 5237 8891 5265
tri 8891 5237 8919 5265 sw
tri 9287 5237 9315 5265 se
rect 9315 5237 9445 5265
tri 9445 5237 9473 5265 sw
tri 9841 5237 9869 5265 se
rect 9869 5237 9999 5265
tri 9999 5237 10027 5265 sw
tri 10395 5237 10423 5265 se
rect 10423 5237 10553 5265
tri 10553 5237 10581 5265 sw
tri 10949 5237 10977 5265 se
rect 10977 5237 11107 5265
tri 11107 5237 11135 5265 sw
tri 11503 5237 11531 5265 se
rect 11531 5237 11661 5265
tri 11661 5237 11689 5265 sw
tri 12057 5237 12085 5265 se
rect 12085 5237 12215 5265
tri 12215 5237 12243 5265 sw
tri 12611 5237 12639 5265 se
rect 12639 5237 12769 5265
tri 12769 5237 12797 5265 sw
tri 13019 5237 13047 5265 se
rect 13047 5254 13200 5265
rect 13252 5254 13270 5306
rect 13322 5254 13340 5306
rect 13392 5254 13410 5306
rect 13462 5254 13480 5306
rect 13532 5254 13550 5306
rect 13047 5242 13490 5254
rect 13524 5242 13562 5254
rect 13596 5242 13602 5254
rect 13047 5237 13200 5242
rect 2249 5197 13200 5237
rect 13252 5197 13270 5242
rect 13322 5197 13340 5242
rect 13392 5197 13410 5242
rect 2249 5163 2287 5197
rect 2321 5163 2360 5197
rect 2394 5163 2433 5197
rect 2467 5163 2506 5197
rect 2540 5163 2579 5197
rect 2613 5163 2652 5197
rect 2686 5163 2725 5197
rect 2759 5163 2798 5197
rect 2832 5163 2871 5197
rect 2905 5163 2944 5197
rect 2978 5163 3017 5197
rect 3051 5163 3090 5197
rect 3124 5163 3163 5197
rect 3197 5163 3236 5197
rect 3270 5163 3309 5197
rect 3343 5163 3382 5197
rect 3416 5163 3455 5197
rect 3489 5163 3528 5197
rect 3562 5163 3601 5197
rect 3635 5163 3674 5197
rect 3708 5163 3747 5197
rect 3781 5163 3820 5197
rect 3854 5163 3893 5197
rect 3927 5163 3966 5197
rect 4000 5163 4039 5197
rect 4073 5163 4112 5197
rect 4146 5163 4185 5197
rect 4219 5163 4258 5197
rect 4292 5163 4331 5197
rect 4365 5163 4404 5197
rect 4438 5163 4477 5197
rect 4511 5163 4550 5197
rect 4584 5163 4623 5197
rect 4657 5163 4696 5197
rect 4730 5163 4769 5197
rect 4803 5163 4842 5197
rect 4876 5163 4915 5197
rect 4949 5163 4988 5197
rect 5022 5163 5061 5197
rect 5095 5163 5134 5197
rect 5168 5163 5207 5197
rect 5241 5163 5280 5197
rect 5314 5163 5353 5197
rect 5387 5163 5426 5197
rect 13462 5190 13480 5242
rect 13532 5190 13550 5242
rect 13452 5178 13490 5190
rect 13524 5178 13562 5190
rect 13596 5178 13602 5190
rect 2249 5125 5426 5163
rect 13462 5126 13480 5178
rect 13532 5126 13550 5178
rect 2249 5091 2287 5125
rect 2321 5091 2360 5125
rect 2394 5091 2433 5125
rect 2467 5091 2506 5125
rect 2540 5091 2579 5125
rect 2613 5091 2652 5125
rect 2686 5091 2725 5125
rect 2759 5091 2798 5125
rect 2832 5091 2871 5125
rect 2905 5091 2944 5125
rect 2978 5091 3017 5125
rect 3051 5091 3090 5125
rect 3124 5091 3163 5125
rect 3197 5091 3236 5125
rect 3270 5091 3309 5125
rect 3343 5091 3382 5125
rect 3416 5091 3455 5125
rect 3489 5091 3528 5125
rect 3562 5091 3601 5125
rect 3635 5091 3674 5125
rect 3708 5091 3747 5125
rect 3781 5091 3820 5125
rect 3854 5091 3893 5125
rect 3927 5091 3966 5125
rect 4000 5091 4039 5125
rect 4073 5091 4112 5125
rect 4146 5091 4185 5125
rect 4219 5091 4258 5125
rect 4292 5091 4331 5125
rect 4365 5091 4404 5125
rect 4438 5091 4477 5125
rect 4511 5091 4550 5125
rect 4584 5091 4623 5125
rect 4657 5091 4696 5125
rect 4730 5091 4769 5125
rect 4803 5091 4842 5125
rect 4876 5091 4915 5125
rect 4949 5091 4988 5125
rect 5022 5091 5061 5125
rect 5095 5091 5134 5125
rect 5168 5091 5207 5125
rect 5241 5091 5280 5125
rect 5314 5091 5353 5125
rect 5387 5091 5426 5125
rect 13452 5119 13602 5126
rect 13452 5114 13490 5119
rect 13524 5114 13562 5119
rect 13596 5114 13602 5119
rect 2249 5053 5426 5091
rect 13462 5062 13480 5114
rect 13532 5062 13550 5114
rect 2249 5019 2287 5053
rect 2321 5019 2360 5053
rect 2394 5019 2433 5053
rect 2467 5019 2506 5053
rect 2540 5019 2579 5053
rect 2613 5019 2652 5053
rect 2686 5019 2725 5053
rect 2759 5019 2798 5053
rect 2832 5019 2871 5053
rect 2905 5019 2944 5053
rect 2978 5019 3017 5053
rect 3051 5019 3090 5053
rect 3124 5019 3163 5053
rect 3197 5019 3236 5053
rect 3270 5019 3309 5053
rect 3343 5019 3382 5053
rect 3416 5019 3455 5053
rect 3489 5019 3528 5053
rect 3562 5019 3601 5053
rect 3635 5019 3674 5053
rect 3708 5019 3747 5053
rect 3781 5019 3820 5053
rect 3854 5019 3893 5053
rect 3927 5019 3966 5053
rect 4000 5019 4039 5053
rect 4073 5019 4112 5053
rect 4146 5019 4185 5053
rect 4219 5019 4258 5053
rect 4292 5019 4331 5053
rect 4365 5019 4404 5053
rect 4438 5019 4477 5053
rect 4511 5019 4550 5053
rect 4584 5019 4623 5053
rect 4657 5019 4696 5053
rect 4730 5019 4769 5053
rect 4803 5019 4842 5053
rect 4876 5019 4915 5053
rect 4949 5019 4988 5053
rect 5022 5019 5061 5053
rect 5095 5019 5134 5053
rect 5168 5019 5207 5053
rect 5241 5019 5280 5053
rect 5314 5019 5353 5053
rect 5387 5019 5426 5053
rect 13452 5049 13602 5062
rect 2249 4997 13200 5019
rect 13252 4997 13270 5019
rect 13322 4997 13340 5019
rect 13392 4997 13410 5019
rect 13462 4997 13480 5049
rect 13532 4997 13550 5049
rect 2249 4991 13602 4997
rect 13832 6895 13838 7071
rect 13944 6895 13950 21329
rect 13832 6856 13950 6895
rect 13832 6822 13838 6856
rect 13872 6822 13910 6856
rect 13944 6822 13950 6856
rect 13832 6783 13950 6822
rect 13832 6749 13838 6783
rect 13872 6749 13910 6783
rect 13944 6749 13950 6783
rect 13832 6710 13950 6749
rect 13832 6676 13838 6710
rect 13872 6676 13910 6710
rect 13944 6676 13950 6710
rect 13832 6637 13950 6676
rect 13832 6603 13838 6637
rect 13872 6603 13910 6637
rect 13944 6603 13950 6637
rect 13832 6564 13950 6603
rect 13832 6530 13838 6564
rect 13872 6530 13910 6564
rect 13944 6530 13950 6564
rect 13832 6491 13950 6530
rect 13832 6457 13838 6491
rect 13872 6457 13910 6491
rect 13944 6457 13950 6491
rect 13832 6418 13950 6457
rect 13832 6384 13838 6418
rect 13872 6384 13910 6418
rect 13944 6384 13950 6418
rect 13832 6345 13950 6384
rect 13832 6311 13838 6345
rect 13872 6311 13910 6345
rect 13944 6311 13950 6345
rect 13832 6272 13950 6311
rect 13832 6238 13838 6272
rect 13872 6238 13910 6272
rect 13944 6238 13950 6272
rect 13832 6199 13950 6238
rect 13832 6165 13838 6199
rect 13872 6165 13910 6199
rect 13944 6165 13950 6199
rect 13832 6126 13950 6165
rect 13832 6092 13838 6126
rect 13872 6092 13910 6126
rect 13944 6092 13950 6126
rect 13832 6053 13950 6092
rect 13832 6019 13838 6053
rect 13872 6019 13910 6053
rect 13944 6019 13950 6053
rect 13832 5980 13950 6019
rect 13832 5946 13838 5980
rect 13872 5946 13910 5980
rect 13944 5946 13950 5980
rect 13832 5907 13950 5946
rect 13832 5873 13838 5907
rect 13872 5873 13910 5907
rect 13944 5873 13950 5907
rect 13832 5834 13950 5873
rect 13832 5800 13838 5834
rect 13872 5800 13910 5834
rect 13944 5800 13950 5834
rect 13832 5761 13950 5800
rect 13832 5727 13838 5761
rect 13872 5727 13910 5761
rect 13944 5727 13950 5761
rect 13832 5688 13950 5727
rect 13832 5654 13838 5688
rect 13872 5654 13910 5688
rect 13944 5654 13950 5688
rect 13832 5615 13950 5654
rect 13832 5581 13838 5615
rect 13872 5581 13910 5615
rect 13944 5581 13950 5615
rect 13832 5542 13950 5581
rect 13832 5508 13838 5542
rect 13872 5508 13910 5542
rect 13944 5508 13950 5542
rect 13832 5469 13950 5508
rect 13832 5435 13838 5469
rect 13872 5435 13910 5469
rect 13944 5435 13950 5469
rect 13832 5396 13950 5435
rect 13832 5362 13838 5396
rect 13872 5362 13910 5396
rect 13944 5362 13950 5396
rect 13832 5323 13950 5362
rect 13832 5289 13838 5323
rect 13872 5289 13910 5323
rect 13944 5289 13950 5323
rect 13832 5250 13950 5289
rect 13832 5216 13838 5250
rect 13872 5216 13910 5250
rect 13944 5216 13950 5250
rect 13832 5177 13950 5216
rect 13832 5143 13838 5177
rect 13872 5143 13910 5177
rect 13944 5143 13950 5177
rect 13832 5104 13950 5143
rect 13832 5070 13838 5104
rect 13872 5070 13910 5104
rect 13944 5070 13950 5104
rect 13832 5031 13950 5070
rect 13832 4997 13838 5031
rect 13872 4997 13910 5031
rect 13944 4997 13950 5031
rect 1938 4943 2056 4983
rect 1938 4909 1944 4943
rect 1978 4909 2016 4943
rect 2050 4909 2056 4943
rect 13832 4958 13950 4997
rect 13832 4924 13838 4958
rect 13872 4924 13910 4958
rect 13944 4924 13950 4958
rect 1938 4885 2056 4909
tri 13824 4902 13832 4910 se
rect 13832 4902 13950 4924
tri 2056 4885 2073 4902 sw
tri 13807 4885 13824 4902 se
rect 13824 4885 13950 4902
rect 1938 4877 2073 4885
tri 2073 4877 2081 4885 sw
tri 13799 4877 13807 4885 se
rect 13807 4877 13838 4885
rect 1938 4871 4968 4877
rect 5020 4871 5085 4877
rect 5137 4871 5202 4877
rect 5254 4871 13838 4877
tri 1687 4837 1710 4860 sw
rect 1938 4837 1950 4871
rect 1984 4837 2023 4871
rect 2057 4837 2096 4871
rect 2130 4837 2169 4871
rect 2203 4837 2242 4871
rect 2276 4837 2315 4871
rect 2349 4837 2388 4871
rect 2422 4837 2461 4871
rect 2495 4837 2534 4871
rect 2568 4837 2607 4871
rect 2641 4837 2680 4871
rect 2714 4837 2753 4871
rect 2787 4837 2826 4871
rect 2860 4837 2899 4871
rect 2933 4837 2972 4871
rect 3006 4837 3045 4871
rect 3079 4837 3118 4871
rect 3152 4837 3191 4871
rect 3225 4837 3264 4871
rect 3298 4837 3337 4871
rect 3371 4837 3410 4871
rect 3444 4837 3483 4871
rect 3517 4837 3556 4871
rect 3590 4837 3629 4871
rect 3663 4837 3702 4871
rect 3736 4837 3775 4871
rect 3809 4837 3848 4871
rect 3882 4837 3921 4871
rect 3955 4837 3994 4871
rect 4028 4837 4067 4871
rect 4101 4837 4140 4871
rect 4174 4837 4213 4871
rect 4247 4837 4286 4871
rect 4320 4837 4359 4871
rect 4393 4837 4432 4871
rect 4466 4837 4505 4871
rect 4539 4837 4578 4871
rect 4612 4837 4651 4871
rect 4685 4837 4724 4871
rect 4758 4837 4797 4871
rect 4831 4837 4870 4871
rect 4904 4837 4943 4871
rect 5050 4837 5085 4871
rect 5137 4837 5162 4871
rect 5196 4837 5202 4871
rect 1487 4799 1710 4837
tri 1710 4799 1748 4837 sw
rect 1938 4825 4968 4837
rect 5020 4825 5085 4837
rect 5137 4825 5202 4837
rect 13765 4851 13838 4871
rect 13872 4851 13910 4885
rect 13944 4851 13950 4885
rect 1938 4811 5235 4825
rect 13765 4812 13950 4851
rect 1938 4799 4968 4811
rect 5020 4799 5085 4811
rect 5137 4799 5202 4811
rect 1487 4765 1748 4799
tri 1748 4765 1782 4799 sw
rect 1938 4765 1950 4799
rect 1984 4765 2023 4799
rect 2057 4765 2096 4799
rect 2130 4765 2169 4799
rect 2203 4765 2242 4799
rect 2276 4765 2315 4799
rect 2349 4765 2388 4799
rect 2422 4765 2461 4799
rect 2495 4765 2534 4799
rect 2568 4765 2607 4799
rect 2641 4765 2680 4799
rect 2714 4765 2753 4799
rect 2787 4765 2826 4799
rect 2860 4765 2899 4799
rect 2933 4765 2972 4799
rect 3006 4765 3045 4799
rect 3079 4765 3118 4799
rect 3152 4765 3191 4799
rect 3225 4765 3264 4799
rect 3298 4765 3337 4799
rect 3371 4765 3410 4799
rect 3444 4765 3483 4799
rect 3517 4765 3556 4799
rect 3590 4765 3629 4799
rect 3663 4765 3702 4799
rect 3736 4765 3775 4799
rect 3809 4765 3848 4799
rect 3882 4765 3921 4799
rect 3955 4765 3994 4799
rect 4028 4765 4067 4799
rect 4101 4765 4140 4799
rect 4174 4765 4213 4799
rect 4247 4765 4286 4799
rect 4320 4765 4359 4799
rect 4393 4765 4432 4799
rect 4466 4765 4505 4799
rect 4539 4765 4578 4799
rect 4612 4765 4651 4799
rect 4685 4765 4724 4799
rect 4758 4765 4797 4799
rect 4831 4765 4870 4799
rect 4904 4765 4943 4799
rect 5050 4765 5085 4799
rect 5137 4765 5162 4799
rect 5196 4765 5202 4799
rect 13765 4778 13838 4812
rect 13872 4778 13910 4812
rect 13944 4778 13950 4812
rect 13765 4766 13950 4778
rect 13765 4765 13943 4766
rect 1487 4759 1782 4765
tri 1782 4759 1788 4765 sw
rect 1938 4759 4968 4765
rect 5020 4759 5085 4765
rect 5137 4759 5202 4765
rect 5254 4759 13943 4765
tri 13943 4759 13950 4766 nw
rect 13982 39418 14957 39522
rect 13982 39384 14775 39418
rect 14809 39384 14917 39418
rect 14951 39384 14957 39418
rect 13982 39372 14957 39384
rect 1487 4650 1788 4759
tri 1788 4650 1897 4759 sw
tri 13956 4727 13982 4753 se
rect 13982 4727 14182 39372
tri 14182 39338 14216 39372 nw
rect 10369 4721 14182 4727
rect 10421 4669 10445 4721
rect 10497 4669 14182 4721
rect 1487 4618 9036 4650
tri 9036 4618 9068 4650 sw
rect 10369 4635 14182 4669
rect 1487 4608 9068 4618
tri 9068 4608 9078 4618 sw
rect 1487 4458 9078 4608
tri 8958 4452 8964 4458 ne
rect 8964 4452 9078 4458
tri 9078 4452 9234 4608 sw
rect 10421 4583 10445 4635
rect 10497 4583 14182 4635
rect 10369 4577 14182 4583
tri 13404 4464 13517 4577 ne
tri 8964 4445 8971 4452 ne
rect 8971 4445 9234 4452
tri 1417 4416 1446 4445 sw
tri 8971 4416 9000 4445 ne
rect 9000 4416 9234 4445
rect 1287 4373 8928 4416
tri 8928 4373 8971 4416 sw
tri 9000 4373 9043 4416 ne
rect 9043 4373 9234 4416
rect 1287 4370 8971 4373
tri 8908 4360 8918 4370 ne
rect 8918 4360 8971 4370
tri 914 4332 942 4360 sw
tri 8918 4332 8946 4360 ne
rect 8946 4348 8971 4360
tri 8971 4348 8996 4373 sw
tri 9043 4348 9068 4373 ne
rect 9068 4348 9234 4373
tri 9234 4348 9338 4452 sw
rect 8946 4332 8996 4348
rect 814 4307 6923 4332
tri 6923 4307 6948 4332 sw
tri 8946 4307 8971 4332 ne
rect 8971 4307 8996 4332
tri 8996 4307 9037 4348 sw
tri 9068 4307 9109 4348 ne
rect 9109 4307 13246 4348
rect 814 4302 6948 4307
tri 814 4278 838 4302 ne
rect 838 4278 6948 4302
tri 6948 4278 6977 4307 sw
tri 8971 4278 9000 4307 ne
rect 9000 4278 9037 4307
tri 838 4252 864 4278 ne
rect 864 4252 6977 4278
tri 6889 4221 6920 4252 ne
rect 6920 4241 6977 4252
tri 6977 4241 7014 4278 sw
tri 9000 4241 9037 4278 ne
tri 9037 4241 9103 4307 sw
tri 9109 4241 9175 4307 ne
rect 9175 4241 13246 4307
rect 6920 4221 7014 4241
tri 7014 4221 7034 4241 sw
tri 9037 4221 9057 4241 ne
rect 9057 4221 9103 4241
tri 1251 4175 1297 4221 se
rect 1297 4220 5948 4221
rect 1297 4175 5209 4220
tri 1185 4109 1251 4175 se
rect 1251 4168 5209 4175
rect 5261 4168 5278 4220
rect 5330 4168 5346 4220
rect 5398 4168 5414 4220
rect 5466 4168 5482 4220
rect 5534 4168 5550 4220
rect 5602 4168 5618 4220
rect 5670 4168 5686 4220
rect 5738 4168 5754 4220
rect 5806 4168 5822 4220
rect 5874 4168 5890 4220
rect 5942 4168 5948 4220
rect 1251 4109 5948 4168
tri 6920 4164 6977 4221 ne
rect 6977 4175 7034 4221
tri 7034 4175 7080 4221 sw
tri 9057 4175 9103 4221 ne
tri 9103 4175 9169 4241 sw
tri 9175 4175 9241 4241 ne
rect 9241 4175 13246 4241
rect 6977 4164 7080 4175
tri 7080 4164 7091 4175 sw
tri 9103 4164 9114 4175 ne
rect 9114 4171 9169 4175
tri 9169 4171 9173 4175 sw
tri 9241 4171 9245 4175 ne
rect 9245 4171 13246 4175
rect 9114 4164 9173 4171
tri 447 3950 481 3984 se
rect 481 3950 760 3984
tri 419 3922 447 3950 se
rect 447 3922 760 3950
tri 416 3919 419 3922 se
rect 419 3919 760 3922
tri 142 3888 173 3919 se
rect 173 3888 760 3919
tri 90 3836 142 3888 se
rect 142 3836 760 3888
tri 56 3802 90 3836 se
rect 90 3805 760 3836
rect 90 3802 757 3805
tri 757 3802 760 3805 nw
tri 1148 4072 1185 4109 se
rect 1185 4096 5948 4109
rect 1185 4072 5209 4096
rect 1148 4044 5209 4072
rect 5261 4044 5278 4096
rect 5330 4044 5346 4096
rect 5398 4044 5414 4096
rect 5466 4044 5482 4096
rect 5534 4044 5550 4096
rect 5602 4044 5618 4096
rect 5670 4044 5686 4096
rect 5738 4044 5754 4096
rect 5806 4044 5822 4096
rect 5874 4044 5890 4096
rect 5942 4044 5948 4096
tri 6977 4050 7091 4164 ne
tri 7091 4109 7146 4164 sw
tri 9114 4109 9169 4164 ne
rect 9169 4109 9173 4164
tri 9173 4109 9235 4171 sw
tri 12951 4109 13013 4171 ne
rect 13013 4109 13246 4171
rect 7091 4072 7146 4109
tri 7146 4072 7183 4109 sw
tri 9169 4072 9206 4109 ne
rect 9206 4072 12824 4109
tri 12824 4072 12861 4109 sw
tri 13013 4072 13050 4109 ne
rect 13050 4072 13246 4109
rect 7091 4050 7183 4072
tri 7183 4050 7205 4072 sw
tri 9206 4050 9228 4072 ne
rect 9228 4058 12861 4072
tri 12861 4058 12875 4072 sw
tri 13050 4058 13064 4072 ne
rect 9228 4050 12875 4058
tri 7091 4044 7097 4050 ne
rect 7097 4044 7205 4050
tri 7205 4044 7211 4050 sw
tri 9228 4044 9234 4050 ne
rect 9234 4044 12875 4050
rect 1148 4029 1590 4044
tri 1590 4029 1605 4044 nw
tri 7097 4029 7112 4044 ne
rect 7112 4029 7211 4044
tri 7211 4029 7226 4044 sw
tri 9234 4029 9249 4044 ne
rect 9249 4029 12875 4044
rect 1148 4012 1573 4029
tri 1573 4012 1590 4029 nw
tri 7112 4012 7129 4029 ne
rect 7129 4012 7226 4029
tri 7226 4012 7243 4029 sw
tri 12790 4012 12807 4029 ne
rect 12807 4012 12875 4029
rect 1148 3984 1545 4012
tri 1545 3984 1573 4012 nw
tri 1615 3984 1643 4012 se
rect 1643 3984 1886 4012
rect 1148 3974 1535 3984
tri 1535 3974 1545 3984 nw
tri 1605 3974 1615 3984 se
rect 1615 3974 1668 3984
rect 1148 3958 1519 3974
tri 1519 3958 1535 3974 nw
tri 1589 3958 1605 3974 se
rect 1605 3958 1668 3974
rect 1148 3950 1511 3958
tri 1511 3950 1519 3958 nw
tri 1581 3950 1589 3958 se
rect 1589 3950 1668 3958
rect 1702 3950 1753 3984
rect 1787 3950 1838 3984
rect 1872 3950 1886 3984
rect 1148 3924 1485 3950
tri 1485 3924 1511 3950 nw
tri 1555 3924 1581 3950 se
rect 1581 3932 1886 3950
tri 7129 3936 7205 4012 ne
rect 7205 3958 7243 4012
tri 7243 3958 7297 4012 sw
tri 12807 3958 12861 4012 ne
rect 12861 3958 12875 4012
tri 12875 3958 12975 4058 sw
rect 7205 3936 7297 3958
tri 7297 3936 7319 3958 sw
tri 12861 3936 12883 3958 ne
rect 12883 3936 12975 3958
tri 7205 3932 7209 3936 ne
rect 7209 3932 11514 3936
rect 1581 3924 1669 3932
tri 1669 3924 1677 3932 nw
tri 7209 3924 7217 3932 ne
rect 7217 3924 11514 3932
tri 12883 3924 12895 3936 ne
rect 1148 3922 1483 3924
tri 1483 3922 1485 3924 nw
tri 1553 3922 1555 3924 se
rect 1555 3922 1667 3924
tri 1667 3922 1669 3924 nw
tri 7217 3922 7219 3924 ne
rect 7219 3922 11514 3924
rect 1148 3898 1459 3922
tri 1459 3898 1483 3922 nw
tri 1529 3898 1553 3922 se
rect 1553 3898 1643 3922
tri 1643 3898 1667 3922 nw
tri 7219 3898 7243 3922 ne
rect 7243 3898 11514 3922
rect 1148 3888 1449 3898
tri 1449 3888 1459 3898 nw
tri 1519 3888 1529 3898 se
rect 1529 3888 1633 3898
tri 1633 3888 1643 3898 nw
tri 7243 3888 7253 3898 ne
rect 7253 3888 11514 3898
tri 42 3788 56 3802 se
rect 56 3788 743 3802
tri 743 3788 757 3802 nw
tri 24 3770 42 3788 se
rect 42 3770 725 3788
tri 725 3770 743 3788 nw
tri 1130 3770 1148 3788 se
rect 1148 3770 1428 3888
tri 1428 3867 1449 3888 nw
tri 1498 3867 1519 3888 se
rect 1519 3867 1612 3888
tri 1612 3867 1633 3888 nw
tri 7253 3867 7274 3888 ne
rect 7274 3867 11514 3888
rect 24 3739 694 3770
tri 694 3739 725 3770 nw
tri 1099 3739 1130 3770 se
rect 1130 3739 1428 3770
rect 24 3705 660 3739
tri 660 3705 694 3739 nw
tri 1065 3705 1099 3739 se
rect 1099 3705 1428 3739
rect 24 3680 635 3705
tri 635 3680 660 3705 nw
tri 1040 3680 1065 3705 se
rect 1065 3680 1428 3705
rect 24 3664 352 3680
tri 352 3664 368 3680 nw
tri 1024 3664 1040 3680 se
rect 1040 3664 1428 3680
rect 24 3630 318 3664
tri 318 3630 352 3664 nw
tri 990 3630 1024 3664 se
rect 1024 3630 1428 3664
rect 24 3626 314 3630
tri 314 3626 318 3630 nw
tri 986 3626 990 3630 se
rect 990 3626 1428 3630
rect 24 3595 283 3626
tri 283 3595 314 3626 nw
tri 955 3595 986 3626 se
rect 986 3595 1428 3626
rect 24 3592 280 3595
tri 280 3592 283 3595 nw
tri 353 3592 356 3595 se
rect 356 3592 1428 3595
rect 24 3589 277 3592
tri 277 3589 280 3592 nw
tri 350 3589 353 3592 se
rect 353 3589 1428 3592
rect 24 3555 243 3589
tri 243 3555 277 3589 nw
tri 316 3555 350 3589 se
rect 350 3555 368 3589
rect 402 3555 467 3589
rect 501 3555 565 3589
rect 599 3555 1428 3589
rect 24 690 224 3555
tri 224 3536 243 3555 nw
tri 297 3536 316 3555 se
rect 316 3536 1428 3555
tri 283 3522 297 3536 se
rect 297 3522 1428 3536
tri 281 3520 283 3522 se
rect 283 3520 1428 3522
tri 278 3517 281 3520 se
rect 281 3517 1428 3520
tri 264 3503 278 3517 se
rect 278 3503 368 3517
rect 264 3483 368 3503
rect 402 3483 467 3517
rect 501 3483 565 3517
rect 599 3483 1428 3517
rect 264 3442 1428 3483
rect 264 3408 345 3442
rect 379 3408 420 3442
rect 454 3408 494 3442
rect 528 3408 568 3442
rect 602 3408 642 3442
rect 676 3408 716 3442
rect 750 3408 791 3442
rect 825 3408 866 3442
rect 900 3408 941 3442
rect 975 3408 1016 3442
rect 1050 3408 1091 3442
rect 1125 3408 1166 3442
rect 1200 3408 1241 3442
rect 1275 3408 1316 3442
rect 1350 3408 1428 3442
rect 264 3370 1428 3408
rect 264 3336 270 3370
rect 304 3336 1388 3370
rect 1422 3336 1428 3370
rect 264 3322 1428 3336
rect 264 3297 369 3322
rect 264 3263 270 3297
rect 304 3288 369 3297
rect 403 3288 553 3322
rect 587 3288 737 3322
rect 771 3288 921 3322
rect 955 3288 1105 3322
rect 1139 3288 1289 3322
rect 1323 3298 1428 3322
rect 1323 3288 1388 3298
rect 304 3264 1388 3288
rect 1422 3264 1428 3298
rect 304 3263 1428 3264
rect 264 3248 1428 3263
rect 264 3224 369 3248
rect 264 3190 270 3224
rect 304 3214 369 3224
rect 403 3214 553 3248
rect 587 3214 737 3248
rect 771 3214 921 3248
rect 955 3214 1105 3248
rect 1139 3214 1289 3248
rect 1323 3226 1428 3248
rect 1323 3214 1388 3226
rect 304 3192 1388 3214
rect 1422 3192 1428 3226
rect 304 3190 1428 3192
rect 264 3174 1428 3190
rect 264 3151 369 3174
rect 264 3117 270 3151
rect 304 3140 369 3151
rect 403 3164 553 3174
rect 403 3140 419 3164
tri 419 3140 443 3164 nw
tri 513 3140 537 3164 ne
rect 537 3140 553 3164
rect 587 3164 737 3174
rect 587 3140 603 3164
tri 603 3140 627 3164 nw
tri 697 3140 721 3164 ne
rect 721 3140 737 3164
rect 771 3164 921 3174
rect 771 3140 787 3164
tri 787 3140 811 3164 nw
tri 881 3140 905 3164 ne
rect 905 3140 921 3164
rect 955 3164 1105 3174
rect 955 3140 971 3164
tri 971 3140 995 3164 nw
tri 1065 3140 1089 3164 ne
rect 1089 3140 1105 3164
rect 1139 3164 1289 3174
rect 1139 3140 1155 3164
tri 1155 3140 1179 3164 nw
tri 1249 3140 1273 3164 ne
rect 1273 3140 1289 3164
rect 1323 3154 1428 3174
rect 1323 3140 1388 3154
rect 304 3117 409 3140
tri 409 3130 419 3140 nw
tri 537 3130 547 3140 ne
rect 264 3100 409 3117
rect 547 3100 593 3140
tri 593 3130 603 3140 nw
tri 721 3130 731 3140 ne
rect 731 3100 777 3140
tri 777 3130 787 3140 nw
tri 905 3130 915 3140 ne
rect 915 3100 961 3140
tri 961 3130 971 3140 nw
tri 1089 3130 1099 3140 ne
rect 1099 3100 1145 3140
tri 1145 3130 1155 3140 nw
tri 1273 3130 1283 3140 ne
rect 1283 3120 1388 3140
rect 1422 3120 1428 3154
rect 1283 3100 1428 3120
rect 264 3078 369 3100
rect 264 3044 270 3078
rect 304 3066 369 3078
rect 403 3066 409 3100
rect 304 3044 409 3066
rect 264 3026 409 3044
rect 264 3005 369 3026
rect 264 2971 270 3005
rect 304 2992 369 3005
rect 403 2992 409 3026
rect 304 2971 409 2992
rect 264 2951 409 2971
rect 264 2932 369 2951
rect 264 2898 270 2932
rect 304 2917 369 2932
rect 403 2917 409 2951
rect 304 2898 409 2917
rect 264 2876 409 2898
rect 264 2859 369 2876
rect 264 2825 270 2859
rect 304 2842 369 2859
rect 403 2842 409 2876
rect 304 2825 409 2842
rect 264 2801 409 2825
rect 264 2786 369 2801
rect 264 2752 270 2786
rect 304 2767 369 2786
rect 403 2767 409 2801
rect 304 2752 409 2767
rect 264 2726 409 2752
rect 264 2713 369 2726
rect 264 2679 270 2713
rect 304 2692 369 2713
rect 403 2692 409 2726
rect 304 2679 409 2692
rect 264 2651 409 2679
rect 264 2640 369 2651
rect 264 2606 270 2640
rect 304 2617 369 2640
rect 403 2617 409 2651
rect 304 2606 409 2617
rect 264 2576 409 2606
rect 264 2567 369 2576
rect 264 2533 270 2567
rect 304 2542 369 2567
rect 403 2542 409 2576
rect 304 2533 409 2542
rect 264 2501 409 2533
rect 264 2494 369 2501
rect 264 2460 270 2494
rect 304 2467 369 2494
rect 403 2467 409 2501
rect 304 2460 409 2467
rect 264 2426 409 2460
rect 264 2421 369 2426
rect 264 2387 270 2421
rect 304 2392 369 2421
rect 403 2392 409 2426
rect 304 2387 409 2392
rect 264 2351 409 2387
rect 264 2348 369 2351
rect 264 2314 270 2348
rect 304 2317 369 2348
rect 403 2317 409 2351
rect 304 2314 409 2317
rect 264 2276 409 2314
rect 264 2242 270 2276
rect 304 2242 369 2276
rect 403 2242 409 2276
rect 264 2204 409 2242
rect 264 2170 270 2204
rect 304 2201 409 2204
rect 304 2170 369 2201
rect 264 2167 369 2170
rect 403 2167 409 2201
rect 264 2132 409 2167
rect 264 2098 270 2132
rect 304 2126 409 2132
rect 304 2098 369 2126
rect 264 2092 369 2098
rect 403 2092 409 2126
rect 264 2060 409 2092
rect 264 2026 270 2060
rect 304 2051 409 2060
rect 304 2026 369 2051
rect 264 2017 369 2026
rect 403 2017 409 2051
rect 264 1988 409 2017
rect 264 1954 270 1988
rect 304 1976 409 1988
rect 304 1954 369 1976
rect 264 1942 369 1954
rect 403 1942 409 1976
rect 264 1916 409 1942
rect 264 1882 270 1916
rect 304 1882 409 1916
rect 264 1844 409 1882
rect 264 1810 270 1844
rect 304 1810 409 1844
rect 264 1792 409 1810
rect 264 1772 369 1792
rect 264 1738 270 1772
rect 304 1758 369 1772
rect 403 1758 409 1792
rect 304 1738 409 1758
rect 264 1718 409 1738
rect 264 1700 369 1718
rect 264 1666 270 1700
rect 304 1684 369 1700
rect 403 1684 409 1718
rect 304 1666 409 1684
rect 264 1644 409 1666
rect 264 1628 369 1644
rect 264 1594 270 1628
rect 304 1610 369 1628
rect 403 1610 409 1644
rect 304 1594 409 1610
rect 264 1570 409 1594
rect 264 1556 369 1570
rect 264 1522 270 1556
rect 304 1536 369 1556
rect 403 1536 409 1570
rect 304 1522 409 1536
rect 264 1496 409 1522
rect 264 1484 369 1496
rect 264 1450 270 1484
rect 304 1462 369 1484
rect 403 1462 409 1496
rect 304 1450 409 1462
rect 264 1422 409 1450
rect 264 1412 369 1422
rect 264 1378 270 1412
rect 304 1388 369 1412
rect 403 1388 409 1422
rect 304 1378 409 1388
rect 264 1348 409 1378
rect 264 1340 369 1348
rect 264 1306 270 1340
rect 304 1314 369 1340
rect 403 1314 409 1348
rect 304 1306 409 1314
rect 264 1274 409 1306
rect 264 1268 369 1274
rect 264 1234 270 1268
rect 304 1240 369 1268
rect 403 1240 409 1274
rect 304 1234 409 1240
rect 264 1200 409 1234
rect 264 1196 369 1200
rect 264 1162 270 1196
rect 304 1166 369 1196
rect 403 1166 409 1200
rect 304 1162 409 1166
rect 264 1126 409 1162
rect 264 1124 369 1126
rect 264 1090 270 1124
rect 304 1092 369 1124
rect 403 1092 409 1126
rect 304 1090 409 1092
rect 264 1052 409 1090
rect 264 1018 270 1052
rect 304 1018 369 1052
rect 403 1018 409 1052
rect 264 980 409 1018
rect 264 946 270 980
rect 304 978 409 980
rect 304 946 369 978
rect 264 944 369 946
rect 403 944 409 978
rect 264 908 409 944
rect 264 874 270 908
rect 304 903 409 908
rect 304 874 369 903
rect 264 869 369 874
rect 403 869 409 903
rect 264 862 409 869
tri 329 836 355 862 ne
rect 355 836 409 862
tri 355 830 361 836 ne
rect 361 830 409 836
tri 361 828 363 830 ne
rect 363 828 409 830
rect 363 794 369 828
rect 403 794 409 828
rect 363 753 409 794
rect 363 719 369 753
rect 403 719 409 753
tri 224 690 234 700 sw
rect 24 682 234 690
tri 234 682 242 690 sw
rect 24 678 242 682
tri 242 678 246 682 sw
rect 363 678 409 719
rect 24 644 246 678
tri 246 644 280 678 sw
rect 363 644 369 678
rect 403 644 409 678
rect 24 637 280 644
tri 280 637 287 644 sw
rect 24 632 287 637
tri 287 632 292 637 sw
rect 363 632 409 644
rect 455 3088 501 3100
rect 455 3054 461 3088
rect 495 3054 501 3088
rect 455 3015 501 3054
rect 455 2981 461 3015
rect 495 2981 501 3015
rect 455 2942 501 2981
rect 455 2908 461 2942
rect 495 2908 501 2942
rect 455 2869 501 2908
rect 455 2835 461 2869
rect 495 2835 501 2869
rect 455 2796 501 2835
rect 455 2762 461 2796
rect 495 2762 501 2796
rect 455 2723 501 2762
rect 455 2689 461 2723
rect 495 2689 501 2723
rect 455 2650 501 2689
rect 455 2616 461 2650
rect 495 2616 501 2650
rect 455 2577 501 2616
rect 455 2543 461 2577
rect 495 2543 501 2577
rect 455 2504 501 2543
rect 455 2470 461 2504
rect 495 2470 501 2504
rect 455 2431 501 2470
rect 455 2397 461 2431
rect 495 2397 501 2431
rect 455 2358 501 2397
rect 455 2324 461 2358
rect 495 2324 501 2358
rect 455 2284 501 2324
rect 455 2250 461 2284
rect 495 2250 501 2284
rect 455 2210 501 2250
rect 455 2176 461 2210
rect 495 2176 501 2210
rect 455 2136 501 2176
rect 455 2102 461 2136
rect 495 2102 501 2136
rect 455 2062 501 2102
rect 455 2028 461 2062
rect 495 2028 501 2062
rect 455 1792 501 2028
rect 455 1758 461 1792
rect 495 1758 501 1792
rect 455 1718 501 1758
rect 455 1684 461 1718
rect 495 1684 501 1718
rect 455 1644 501 1684
rect 455 1610 461 1644
rect 495 1610 501 1644
rect 455 1570 501 1610
rect 455 1536 461 1570
rect 495 1536 501 1570
rect 455 1496 501 1536
rect 455 1462 461 1496
rect 495 1462 501 1496
rect 455 1422 501 1462
rect 455 1388 461 1422
rect 495 1388 501 1422
rect 455 1348 501 1388
rect 455 1314 461 1348
rect 495 1314 501 1348
rect 455 1274 501 1314
rect 455 1240 461 1274
rect 495 1240 501 1274
rect 455 1200 501 1240
rect 455 1166 461 1200
rect 495 1166 501 1200
rect 455 1126 501 1166
rect 455 1092 461 1126
rect 495 1092 501 1126
rect 455 1052 501 1092
rect 455 1018 461 1052
rect 495 1018 501 1052
rect 455 978 501 1018
rect 455 944 461 978
rect 495 944 501 978
rect 455 904 501 944
rect 455 870 461 904
rect 495 870 501 904
rect 455 830 501 870
rect 455 796 461 830
rect 495 796 501 830
rect 455 756 501 796
rect 455 722 461 756
rect 495 722 501 756
rect 455 682 501 722
rect 455 648 461 682
rect 495 648 501 682
tri 453 632 455 634 se
rect 455 632 501 648
rect 547 3066 553 3100
rect 587 3066 593 3100
rect 547 3026 593 3066
rect 547 2992 553 3026
rect 587 2992 593 3026
rect 547 2951 593 2992
rect 547 2917 553 2951
rect 587 2917 593 2951
rect 547 2876 593 2917
rect 547 2842 553 2876
rect 587 2842 593 2876
rect 547 2801 593 2842
rect 547 2767 553 2801
rect 587 2767 593 2801
rect 547 2726 593 2767
rect 547 2692 553 2726
rect 587 2692 593 2726
rect 547 2651 593 2692
rect 547 2617 553 2651
rect 587 2617 593 2651
rect 547 2576 593 2617
rect 547 2542 553 2576
rect 587 2542 593 2576
rect 547 2501 593 2542
rect 547 2467 553 2501
rect 587 2467 593 2501
rect 547 2426 593 2467
rect 547 2392 553 2426
rect 587 2392 593 2426
rect 547 2351 593 2392
rect 547 2317 553 2351
rect 587 2317 593 2351
rect 547 2276 593 2317
rect 547 2242 553 2276
rect 587 2242 593 2276
rect 547 2201 593 2242
rect 547 2167 553 2201
rect 587 2167 593 2201
rect 547 2126 593 2167
rect 547 2092 553 2126
rect 587 2092 593 2126
rect 547 2051 593 2092
rect 547 2017 553 2051
rect 587 2017 593 2051
rect 547 1976 593 2017
rect 547 1942 553 1976
rect 587 1942 593 1976
rect 547 1792 593 1942
rect 547 1758 553 1792
rect 587 1758 593 1792
rect 547 1718 593 1758
rect 547 1684 553 1718
rect 587 1684 593 1718
rect 547 1644 593 1684
rect 547 1610 553 1644
rect 587 1610 593 1644
rect 547 1570 593 1610
rect 547 1536 553 1570
rect 587 1536 593 1570
rect 547 1496 593 1536
rect 547 1462 553 1496
rect 587 1462 593 1496
rect 547 1422 593 1462
rect 547 1388 553 1422
rect 587 1388 593 1422
rect 547 1348 593 1388
rect 547 1314 553 1348
rect 587 1314 593 1348
rect 547 1274 593 1314
rect 547 1240 553 1274
rect 587 1240 593 1274
rect 547 1200 593 1240
rect 547 1166 553 1200
rect 587 1166 593 1200
rect 547 1126 593 1166
rect 547 1092 553 1126
rect 587 1092 593 1126
rect 547 1052 593 1092
rect 547 1018 553 1052
rect 587 1018 593 1052
rect 547 978 593 1018
rect 547 944 553 978
rect 587 944 593 978
rect 547 903 593 944
rect 547 869 553 903
rect 587 869 593 903
rect 547 828 593 869
rect 547 794 553 828
rect 587 794 593 828
rect 547 753 593 794
rect 547 719 553 753
rect 587 719 593 753
rect 547 678 593 719
rect 547 644 553 678
rect 587 644 593 678
tri 501 632 503 634 sw
rect 547 632 593 644
rect 639 3088 685 3100
rect 639 3054 645 3088
rect 679 3054 685 3088
rect 639 3015 685 3054
rect 639 2981 645 3015
rect 679 2981 685 3015
rect 639 2942 685 2981
rect 639 2908 645 2942
rect 679 2908 685 2942
rect 639 2869 685 2908
rect 639 2835 645 2869
rect 679 2835 685 2869
rect 639 2796 685 2835
rect 639 2762 645 2796
rect 679 2762 685 2796
rect 639 2723 685 2762
rect 639 2689 645 2723
rect 679 2689 685 2723
rect 639 2650 685 2689
rect 639 2616 645 2650
rect 679 2616 685 2650
rect 639 2577 685 2616
rect 639 2543 645 2577
rect 679 2543 685 2577
rect 639 2504 685 2543
rect 639 2470 645 2504
rect 679 2470 685 2504
rect 639 2431 685 2470
rect 639 2397 645 2431
rect 679 2397 685 2431
rect 639 2358 685 2397
rect 639 2324 645 2358
rect 679 2324 685 2358
rect 639 2284 685 2324
rect 639 2250 645 2284
rect 679 2250 685 2284
rect 639 2210 685 2250
rect 639 2176 645 2210
rect 679 2176 685 2210
rect 639 2136 685 2176
rect 639 2102 645 2136
rect 679 2102 685 2136
rect 639 2062 685 2102
rect 639 2028 645 2062
rect 679 2028 685 2062
rect 639 1792 685 2028
rect 639 1758 645 1792
rect 679 1758 685 1792
rect 639 1718 685 1758
rect 639 1684 645 1718
rect 679 1684 685 1718
rect 639 1644 685 1684
rect 639 1610 645 1644
rect 679 1610 685 1644
rect 639 1570 685 1610
rect 639 1536 645 1570
rect 679 1536 685 1570
rect 639 1496 685 1536
rect 639 1462 645 1496
rect 679 1462 685 1496
rect 639 1422 685 1462
rect 639 1388 645 1422
rect 679 1388 685 1422
rect 639 1348 685 1388
rect 639 1314 645 1348
rect 679 1314 685 1348
rect 639 1274 685 1314
rect 639 1240 645 1274
rect 679 1240 685 1274
rect 639 1200 685 1240
rect 639 1166 645 1200
rect 679 1166 685 1200
rect 639 1126 685 1166
rect 639 1092 645 1126
rect 679 1092 685 1126
rect 639 1052 685 1092
rect 639 1018 645 1052
rect 679 1018 685 1052
rect 639 978 685 1018
rect 639 944 645 978
rect 679 944 685 978
rect 639 904 685 944
rect 639 870 645 904
rect 679 870 685 904
rect 639 830 685 870
rect 639 796 645 830
rect 679 796 685 830
rect 639 756 685 796
rect 639 722 645 756
rect 679 722 685 756
rect 639 682 685 722
rect 639 648 645 682
rect 679 648 685 682
tri 637 632 639 634 se
rect 639 632 685 648
rect 731 3066 737 3100
rect 771 3066 777 3100
rect 731 3026 777 3066
rect 731 2992 737 3026
rect 771 2992 777 3026
rect 731 2951 777 2992
rect 731 2917 737 2951
rect 771 2917 777 2951
rect 731 2876 777 2917
rect 731 2842 737 2876
rect 771 2842 777 2876
rect 731 2801 777 2842
rect 731 2767 737 2801
rect 771 2767 777 2801
rect 731 2726 777 2767
rect 731 2692 737 2726
rect 771 2692 777 2726
rect 731 2651 777 2692
rect 731 2617 737 2651
rect 771 2617 777 2651
rect 731 2576 777 2617
rect 731 2542 737 2576
rect 771 2542 777 2576
rect 731 2501 777 2542
rect 731 2467 737 2501
rect 771 2467 777 2501
rect 731 2426 777 2467
rect 731 2392 737 2426
rect 771 2392 777 2426
rect 731 2351 777 2392
rect 731 2317 737 2351
rect 771 2317 777 2351
rect 731 2276 777 2317
rect 731 2242 737 2276
rect 771 2242 777 2276
rect 731 2201 777 2242
rect 731 2167 737 2201
rect 771 2167 777 2201
rect 731 2126 777 2167
rect 731 2092 737 2126
rect 771 2092 777 2126
rect 731 2051 777 2092
rect 731 2017 737 2051
rect 771 2017 777 2051
rect 731 1976 777 2017
rect 731 1942 737 1976
rect 771 1942 777 1976
rect 731 1792 777 1942
rect 731 1758 737 1792
rect 771 1758 777 1792
rect 731 1718 777 1758
rect 731 1684 737 1718
rect 771 1684 777 1718
rect 731 1644 777 1684
rect 731 1610 737 1644
rect 771 1610 777 1644
rect 731 1570 777 1610
rect 731 1536 737 1570
rect 771 1536 777 1570
rect 731 1496 777 1536
rect 731 1462 737 1496
rect 771 1462 777 1496
rect 731 1422 777 1462
rect 731 1388 737 1422
rect 771 1388 777 1422
rect 731 1348 777 1388
rect 731 1314 737 1348
rect 771 1314 777 1348
rect 731 1274 777 1314
rect 731 1240 737 1274
rect 771 1240 777 1274
rect 731 1200 777 1240
rect 731 1166 737 1200
rect 771 1166 777 1200
rect 731 1126 777 1166
rect 731 1092 737 1126
rect 771 1092 777 1126
rect 731 1052 777 1092
rect 731 1018 737 1052
rect 771 1018 777 1052
rect 731 978 777 1018
rect 731 944 737 978
rect 771 944 777 978
rect 731 903 777 944
rect 731 869 737 903
rect 771 869 777 903
rect 731 828 777 869
rect 731 794 737 828
rect 771 794 777 828
rect 731 753 777 794
rect 731 719 737 753
rect 771 719 777 753
rect 731 678 777 719
rect 731 644 737 678
rect 771 644 777 678
tri 685 632 687 634 sw
rect 731 632 777 644
rect 823 3088 869 3100
rect 823 3054 829 3088
rect 863 3054 869 3088
rect 823 3015 869 3054
rect 823 2981 829 3015
rect 863 2981 869 3015
rect 823 2942 869 2981
rect 823 2908 829 2942
rect 863 2908 869 2942
rect 823 2869 869 2908
rect 823 2835 829 2869
rect 863 2835 869 2869
rect 823 2796 869 2835
rect 823 2762 829 2796
rect 863 2762 869 2796
rect 823 2723 869 2762
rect 823 2689 829 2723
rect 863 2689 869 2723
rect 823 2650 869 2689
rect 823 2616 829 2650
rect 863 2616 869 2650
rect 823 2577 869 2616
rect 823 2543 829 2577
rect 863 2543 869 2577
rect 823 2504 869 2543
rect 823 2470 829 2504
rect 863 2470 869 2504
rect 823 2431 869 2470
rect 823 2397 829 2431
rect 863 2397 869 2431
rect 823 2358 869 2397
rect 823 2324 829 2358
rect 863 2324 869 2358
rect 823 2284 869 2324
rect 823 2250 829 2284
rect 863 2250 869 2284
rect 823 2210 869 2250
rect 823 2176 829 2210
rect 863 2176 869 2210
rect 823 2136 869 2176
rect 823 2102 829 2136
rect 863 2102 869 2136
rect 823 2062 869 2102
rect 823 2028 829 2062
rect 863 2028 869 2062
rect 823 1792 869 2028
rect 823 1758 829 1792
rect 863 1758 869 1792
rect 823 1718 869 1758
rect 823 1684 829 1718
rect 863 1684 869 1718
rect 823 1644 869 1684
rect 823 1610 829 1644
rect 863 1610 869 1644
rect 823 1570 869 1610
rect 823 1536 829 1570
rect 863 1536 869 1570
rect 823 1496 869 1536
rect 823 1462 829 1496
rect 863 1462 869 1496
rect 823 1422 869 1462
rect 823 1388 829 1422
rect 863 1388 869 1422
rect 823 1348 869 1388
rect 823 1314 829 1348
rect 863 1314 869 1348
rect 823 1274 869 1314
rect 823 1240 829 1274
rect 863 1240 869 1274
rect 823 1200 869 1240
rect 823 1166 829 1200
rect 863 1166 869 1200
rect 823 1126 869 1166
rect 823 1092 829 1126
rect 863 1092 869 1126
rect 823 1052 869 1092
rect 823 1018 829 1052
rect 863 1018 869 1052
rect 823 978 869 1018
rect 823 944 829 978
rect 863 944 869 978
rect 823 904 869 944
rect 823 870 829 904
rect 863 870 869 904
rect 823 830 869 870
rect 823 796 829 830
rect 863 796 869 830
rect 823 756 869 796
rect 823 722 829 756
rect 863 722 869 756
rect 823 682 869 722
rect 823 648 829 682
rect 863 648 869 682
tri 821 632 823 634 se
rect 823 632 869 648
rect 915 3066 921 3100
rect 955 3066 961 3100
rect 915 3026 961 3066
rect 915 2992 921 3026
rect 955 2992 961 3026
rect 915 2951 961 2992
rect 915 2917 921 2951
rect 955 2917 961 2951
rect 915 2876 961 2917
rect 915 2842 921 2876
rect 955 2842 961 2876
rect 915 2801 961 2842
rect 915 2767 921 2801
rect 955 2767 961 2801
rect 915 2726 961 2767
rect 915 2692 921 2726
rect 955 2692 961 2726
rect 915 2651 961 2692
rect 915 2617 921 2651
rect 955 2617 961 2651
rect 915 2576 961 2617
rect 915 2542 921 2576
rect 955 2542 961 2576
rect 915 2501 961 2542
rect 915 2467 921 2501
rect 955 2467 961 2501
rect 915 2426 961 2467
rect 915 2392 921 2426
rect 955 2392 961 2426
rect 915 2351 961 2392
rect 915 2317 921 2351
rect 955 2317 961 2351
rect 915 2276 961 2317
rect 915 2242 921 2276
rect 955 2242 961 2276
rect 915 2201 961 2242
rect 915 2167 921 2201
rect 955 2167 961 2201
rect 915 2126 961 2167
rect 915 2092 921 2126
rect 955 2092 961 2126
rect 915 2051 961 2092
rect 915 2017 921 2051
rect 955 2017 961 2051
rect 915 1976 961 2017
rect 915 1942 921 1976
rect 955 1942 961 1976
rect 915 1792 961 1942
rect 915 1758 921 1792
rect 955 1758 961 1792
rect 915 1718 961 1758
rect 915 1684 921 1718
rect 955 1684 961 1718
rect 915 1644 961 1684
rect 915 1610 921 1644
rect 955 1610 961 1644
rect 915 1570 961 1610
rect 915 1536 921 1570
rect 955 1536 961 1570
rect 915 1496 961 1536
rect 915 1462 921 1496
rect 955 1462 961 1496
rect 915 1422 961 1462
rect 915 1388 921 1422
rect 955 1388 961 1422
rect 915 1348 961 1388
rect 915 1314 921 1348
rect 955 1314 961 1348
rect 915 1274 961 1314
rect 915 1240 921 1274
rect 955 1240 961 1274
rect 915 1200 961 1240
rect 915 1166 921 1200
rect 955 1166 961 1200
rect 915 1126 961 1166
rect 915 1092 921 1126
rect 955 1092 961 1126
rect 915 1052 961 1092
rect 915 1018 921 1052
rect 955 1018 961 1052
rect 915 978 961 1018
rect 915 944 921 978
rect 955 944 961 978
rect 915 903 961 944
rect 915 869 921 903
rect 955 869 961 903
rect 915 828 961 869
rect 915 794 921 828
rect 955 794 961 828
rect 915 753 961 794
rect 915 719 921 753
rect 955 719 961 753
rect 915 678 961 719
rect 915 644 921 678
rect 955 644 961 678
tri 869 632 871 634 sw
rect 915 632 961 644
rect 1007 3088 1053 3100
rect 1007 3054 1013 3088
rect 1047 3054 1053 3088
rect 1007 3015 1053 3054
rect 1007 2981 1013 3015
rect 1047 2981 1053 3015
rect 1007 2942 1053 2981
rect 1007 2908 1013 2942
rect 1047 2908 1053 2942
rect 1007 2869 1053 2908
rect 1007 2835 1013 2869
rect 1047 2835 1053 2869
rect 1007 2796 1053 2835
rect 1007 2762 1013 2796
rect 1047 2762 1053 2796
rect 1007 2723 1053 2762
rect 1007 2689 1013 2723
rect 1047 2689 1053 2723
rect 1007 2650 1053 2689
rect 1007 2616 1013 2650
rect 1047 2616 1053 2650
rect 1007 2577 1053 2616
rect 1007 2543 1013 2577
rect 1047 2543 1053 2577
rect 1007 2504 1053 2543
rect 1007 2470 1013 2504
rect 1047 2470 1053 2504
rect 1007 2431 1053 2470
rect 1007 2397 1013 2431
rect 1047 2397 1053 2431
rect 1007 2358 1053 2397
rect 1007 2324 1013 2358
rect 1047 2324 1053 2358
rect 1007 2284 1053 2324
rect 1007 2250 1013 2284
rect 1047 2250 1053 2284
rect 1007 2210 1053 2250
rect 1007 2176 1013 2210
rect 1047 2176 1053 2210
rect 1007 2136 1053 2176
rect 1007 2102 1013 2136
rect 1047 2102 1053 2136
rect 1007 2062 1053 2102
rect 1007 2028 1013 2062
rect 1047 2028 1053 2062
rect 1007 1792 1053 2028
rect 1007 1758 1013 1792
rect 1047 1758 1053 1792
rect 1007 1718 1053 1758
rect 1007 1684 1013 1718
rect 1047 1684 1053 1718
rect 1007 1644 1053 1684
rect 1007 1610 1013 1644
rect 1047 1610 1053 1644
rect 1007 1570 1053 1610
rect 1007 1536 1013 1570
rect 1047 1536 1053 1570
rect 1007 1496 1053 1536
rect 1007 1462 1013 1496
rect 1047 1462 1053 1496
rect 1007 1422 1053 1462
rect 1007 1388 1013 1422
rect 1047 1388 1053 1422
rect 1007 1348 1053 1388
rect 1007 1314 1013 1348
rect 1047 1314 1053 1348
rect 1007 1274 1053 1314
rect 1007 1240 1013 1274
rect 1047 1240 1053 1274
rect 1007 1200 1053 1240
rect 1007 1166 1013 1200
rect 1047 1166 1053 1200
rect 1007 1126 1053 1166
rect 1007 1092 1013 1126
rect 1047 1092 1053 1126
rect 1007 1052 1053 1092
rect 1007 1018 1013 1052
rect 1047 1018 1053 1052
rect 1007 978 1053 1018
rect 1007 944 1013 978
rect 1047 944 1053 978
rect 1007 904 1053 944
rect 1007 870 1013 904
rect 1047 870 1053 904
rect 1007 830 1053 870
rect 1007 796 1013 830
rect 1047 796 1053 830
rect 1007 756 1053 796
rect 1007 722 1013 756
rect 1047 722 1053 756
rect 1007 682 1053 722
rect 1007 648 1013 682
rect 1047 648 1053 682
tri 1005 632 1007 634 se
rect 1007 632 1053 648
rect 1099 3066 1105 3100
rect 1139 3066 1145 3100
rect 1099 3026 1145 3066
rect 1099 2992 1105 3026
rect 1139 2992 1145 3026
rect 1099 2951 1145 2992
rect 1099 2917 1105 2951
rect 1139 2917 1145 2951
rect 1099 2876 1145 2917
rect 1099 2842 1105 2876
rect 1139 2842 1145 2876
rect 1099 2801 1145 2842
rect 1099 2767 1105 2801
rect 1139 2767 1145 2801
rect 1099 2726 1145 2767
rect 1099 2692 1105 2726
rect 1139 2692 1145 2726
rect 1099 2651 1145 2692
rect 1099 2617 1105 2651
rect 1139 2617 1145 2651
rect 1099 2576 1145 2617
rect 1099 2542 1105 2576
rect 1139 2542 1145 2576
rect 1099 2501 1145 2542
rect 1099 2467 1105 2501
rect 1139 2467 1145 2501
rect 1099 2426 1145 2467
rect 1099 2392 1105 2426
rect 1139 2392 1145 2426
rect 1099 2351 1145 2392
rect 1099 2317 1105 2351
rect 1139 2317 1145 2351
rect 1099 2276 1145 2317
rect 1099 2242 1105 2276
rect 1139 2242 1145 2276
rect 1099 2201 1145 2242
rect 1099 2167 1105 2201
rect 1139 2167 1145 2201
rect 1099 2126 1145 2167
rect 1099 2092 1105 2126
rect 1139 2092 1145 2126
rect 1099 2051 1145 2092
rect 1099 2017 1105 2051
rect 1139 2017 1145 2051
rect 1099 1976 1145 2017
rect 1099 1942 1105 1976
rect 1139 1942 1145 1976
rect 1099 1792 1145 1942
rect 1099 1758 1105 1792
rect 1139 1758 1145 1792
rect 1099 1718 1145 1758
rect 1099 1684 1105 1718
rect 1139 1684 1145 1718
rect 1099 1644 1145 1684
rect 1099 1610 1105 1644
rect 1139 1610 1145 1644
rect 1099 1570 1145 1610
rect 1099 1536 1105 1570
rect 1139 1536 1145 1570
rect 1099 1496 1145 1536
rect 1099 1462 1105 1496
rect 1139 1462 1145 1496
rect 1099 1422 1145 1462
rect 1099 1388 1105 1422
rect 1139 1388 1145 1422
rect 1099 1348 1145 1388
rect 1099 1314 1105 1348
rect 1139 1314 1145 1348
rect 1099 1274 1145 1314
rect 1099 1240 1105 1274
rect 1139 1240 1145 1274
rect 1099 1200 1145 1240
rect 1099 1166 1105 1200
rect 1139 1166 1145 1200
rect 1099 1126 1145 1166
rect 1099 1092 1105 1126
rect 1139 1092 1145 1126
rect 1099 1052 1145 1092
rect 1099 1018 1105 1052
rect 1139 1018 1145 1052
rect 1099 978 1145 1018
rect 1099 944 1105 978
rect 1139 944 1145 978
rect 1099 903 1145 944
rect 1099 869 1105 903
rect 1139 869 1145 903
rect 1099 828 1145 869
rect 1099 794 1105 828
rect 1139 794 1145 828
rect 1099 753 1145 794
rect 1099 719 1105 753
rect 1139 719 1145 753
rect 1099 678 1145 719
rect 1099 644 1105 678
rect 1139 644 1145 678
tri 1053 632 1055 634 sw
rect 1099 632 1145 644
rect 1191 3088 1237 3100
rect 1191 3054 1197 3088
rect 1231 3054 1237 3088
rect 1191 3015 1237 3054
rect 1191 2981 1197 3015
rect 1231 2981 1237 3015
rect 1191 2942 1237 2981
rect 1191 2908 1197 2942
rect 1231 2908 1237 2942
rect 1191 2869 1237 2908
rect 1191 2835 1197 2869
rect 1231 2835 1237 2869
rect 1191 2796 1237 2835
rect 1191 2762 1197 2796
rect 1231 2762 1237 2796
rect 1191 2723 1237 2762
rect 1191 2689 1197 2723
rect 1231 2689 1237 2723
rect 1191 2650 1237 2689
rect 1191 2616 1197 2650
rect 1231 2616 1237 2650
rect 1191 2577 1237 2616
rect 1191 2543 1197 2577
rect 1231 2543 1237 2577
rect 1191 2504 1237 2543
rect 1191 2470 1197 2504
rect 1231 2470 1237 2504
rect 1191 2431 1237 2470
rect 1191 2397 1197 2431
rect 1231 2397 1237 2431
rect 1191 2358 1237 2397
rect 1191 2324 1197 2358
rect 1231 2324 1237 2358
rect 1191 2284 1237 2324
rect 1191 2250 1197 2284
rect 1231 2250 1237 2284
rect 1191 2210 1237 2250
rect 1191 2176 1197 2210
rect 1231 2176 1237 2210
rect 1191 2136 1237 2176
rect 1191 2102 1197 2136
rect 1231 2102 1237 2136
rect 1191 2062 1237 2102
rect 1191 2028 1197 2062
rect 1231 2028 1237 2062
rect 1191 1792 1237 2028
rect 1191 1758 1197 1792
rect 1231 1758 1237 1792
rect 1191 1718 1237 1758
rect 1191 1684 1197 1718
rect 1231 1684 1237 1718
rect 1191 1644 1237 1684
rect 1191 1610 1197 1644
rect 1231 1610 1237 1644
rect 1191 1570 1237 1610
rect 1191 1536 1197 1570
rect 1231 1536 1237 1570
rect 1191 1496 1237 1536
rect 1191 1462 1197 1496
rect 1231 1462 1237 1496
rect 1191 1422 1237 1462
rect 1191 1388 1197 1422
rect 1231 1388 1237 1422
rect 1191 1348 1237 1388
rect 1191 1314 1197 1348
rect 1231 1314 1237 1348
rect 1191 1274 1237 1314
rect 1191 1240 1197 1274
rect 1231 1240 1237 1274
rect 1191 1200 1237 1240
rect 1191 1166 1197 1200
rect 1231 1166 1237 1200
rect 1191 1126 1237 1166
rect 1191 1092 1197 1126
rect 1231 1092 1237 1126
rect 1191 1052 1237 1092
rect 1191 1018 1197 1052
rect 1231 1018 1237 1052
rect 1191 978 1237 1018
rect 1191 944 1197 978
rect 1231 944 1237 978
rect 1191 904 1237 944
rect 1191 870 1197 904
rect 1231 870 1237 904
rect 1191 830 1237 870
rect 1191 796 1197 830
rect 1231 796 1237 830
rect 1191 756 1237 796
rect 1191 722 1197 756
rect 1231 722 1237 756
rect 1191 682 1237 722
rect 1191 648 1197 682
rect 1231 648 1237 682
tri 1189 632 1191 634 se
rect 1191 632 1237 648
rect 24 615 292 632
tri 292 615 309 632 sw
tri 436 615 453 632 se
rect 453 615 503 632
tri 503 615 520 632 sw
tri 620 615 637 632 se
rect 637 615 687 632
tri 687 615 704 632 sw
tri 804 615 821 632 se
rect 821 615 871 632
tri 871 615 888 632 sw
tri 988 615 1005 632 se
rect 1005 615 1055 632
tri 1055 615 1072 632 sw
tri 1172 615 1189 632 se
rect 1189 615 1237 632
rect 24 613 309 615
tri 309 613 311 615 sw
tri 434 613 436 615 se
rect 436 613 520 615
tri 520 613 522 615 sw
tri 618 613 620 615 se
rect 620 613 704 615
tri 704 613 706 615 sw
tri 802 613 804 615 se
rect 804 613 888 615
tri 888 613 890 615 sw
tri 986 613 988 615 se
rect 988 613 1072 615
tri 1072 613 1074 615 sw
tri 1170 613 1172 615 se
rect 1172 613 1237 615
rect 24 607 311 613
tri 311 607 317 613 sw
tri 428 607 434 613 se
rect 434 607 522 613
tri 522 607 528 613 sw
tri 612 607 618 613 se
rect 618 607 706 613
tri 706 607 712 613 sw
tri 796 607 802 613 se
rect 802 607 890 613
tri 890 607 896 613 sw
tri 980 607 986 613 se
rect 986 607 1074 613
tri 1074 607 1080 613 sw
tri 1164 607 1170 613 se
rect 1170 607 1237 613
rect 24 577 317 607
tri 317 577 347 607 sw
tri 398 577 428 607 se
rect 428 577 461 607
rect 24 573 461 577
rect 495 600 528 607
tri 528 600 535 607 sw
tri 605 600 612 607 se
rect 612 600 645 607
rect 495 573 645 600
rect 679 600 712 607
tri 712 600 719 607 sw
tri 789 600 796 607 se
rect 796 600 829 607
rect 679 573 829 600
rect 863 600 896 607
tri 896 600 903 607 sw
tri 973 600 980 607 se
rect 980 600 1013 607
rect 863 573 1013 600
rect 1047 600 1080 607
tri 1080 600 1087 607 sw
tri 1157 600 1164 607 se
rect 1164 600 1197 607
rect 1047 573 1197 600
rect 1231 573 1237 607
rect 24 532 1237 573
rect 24 498 461 532
rect 495 498 645 532
rect 679 498 829 532
rect 863 498 1013 532
rect 1047 498 1197 532
rect 1231 498 1237 532
rect 24 400 1237 498
rect 1283 3066 1289 3100
rect 1323 3082 1428 3100
rect 1323 3066 1388 3082
rect 1283 3048 1388 3066
rect 1422 3048 1428 3082
rect 1283 3026 1428 3048
rect 1283 2992 1289 3026
rect 1323 3010 1428 3026
rect 1323 2992 1388 3010
rect 1283 2976 1388 2992
rect 1422 2976 1428 3010
rect 1283 2951 1428 2976
rect 1283 2917 1289 2951
rect 1323 2938 1428 2951
rect 1323 2917 1388 2938
rect 1283 2904 1388 2917
rect 1422 2904 1428 2938
rect 1283 2876 1428 2904
rect 1283 2842 1289 2876
rect 1323 2866 1428 2876
rect 1323 2842 1388 2866
rect 1283 2832 1388 2842
rect 1422 2832 1428 2866
rect 1283 2801 1428 2832
rect 1283 2767 1289 2801
rect 1323 2794 1428 2801
rect 1323 2767 1388 2794
rect 1283 2760 1388 2767
rect 1422 2760 1428 2794
rect 1283 2726 1428 2760
rect 1283 2692 1289 2726
rect 1323 2722 1428 2726
rect 1323 2692 1388 2722
rect 1283 2688 1388 2692
rect 1422 2688 1428 2722
rect 1283 2651 1428 2688
rect 1283 2617 1289 2651
rect 1323 2650 1428 2651
rect 1323 2617 1388 2650
rect 1283 2616 1388 2617
rect 1422 2616 1428 2650
rect 1283 2578 1428 2616
rect 1283 2576 1388 2578
rect 1283 2542 1289 2576
rect 1323 2544 1388 2576
rect 1422 2544 1428 2578
rect 1323 2542 1428 2544
rect 1283 2506 1428 2542
rect 1283 2501 1388 2506
rect 1283 2467 1289 2501
rect 1323 2472 1388 2501
rect 1422 2472 1428 2506
rect 1323 2467 1428 2472
rect 1283 2434 1428 2467
rect 1283 2426 1388 2434
rect 1283 2392 1289 2426
rect 1323 2400 1388 2426
rect 1422 2400 1428 2434
rect 1323 2392 1428 2400
rect 1283 2362 1428 2392
rect 1283 2351 1388 2362
rect 1283 2317 1289 2351
rect 1323 2328 1388 2351
rect 1422 2328 1428 2362
rect 1323 2317 1428 2328
rect 1283 2290 1428 2317
rect 1283 2276 1388 2290
rect 1283 2242 1289 2276
rect 1323 2256 1388 2276
rect 1422 2256 1428 2290
rect 1323 2242 1428 2256
rect 1283 2218 1428 2242
rect 1283 2201 1388 2218
rect 1283 2167 1289 2201
rect 1323 2184 1388 2201
rect 1422 2184 1428 2218
rect 1323 2167 1428 2184
rect 1283 2146 1428 2167
rect 1283 2126 1388 2146
rect 1283 2092 1289 2126
rect 1323 2112 1388 2126
rect 1422 2112 1428 2146
rect 1323 2092 1428 2112
rect 1283 2074 1428 2092
rect 1283 2051 1388 2074
rect 1283 2017 1289 2051
rect 1323 2040 1388 2051
rect 1422 2040 1428 2074
rect 1323 2017 1428 2040
rect 1283 2002 1428 2017
rect 1283 1976 1388 2002
rect 1283 1942 1289 1976
rect 1323 1968 1388 1976
rect 1422 1968 1428 2002
rect 1323 1942 1428 1968
rect 1283 1930 1428 1942
rect 1283 1896 1388 1930
rect 1422 1896 1428 1930
rect 1283 1858 1428 1896
rect 1283 1824 1388 1858
rect 1422 1824 1428 1858
rect 1283 1792 1428 1824
rect 1283 1758 1289 1792
rect 1323 1785 1428 1792
rect 1323 1758 1388 1785
rect 1283 1751 1388 1758
rect 1422 1751 1428 1785
rect 1283 1718 1428 1751
rect 1283 1684 1289 1718
rect 1323 1712 1428 1718
rect 1323 1684 1388 1712
rect 1283 1678 1388 1684
rect 1422 1678 1428 1712
rect 1283 1644 1428 1678
rect 1283 1610 1289 1644
rect 1323 1639 1428 1644
rect 1323 1610 1388 1639
rect 1283 1605 1388 1610
rect 1422 1605 1428 1639
rect 1283 1570 1428 1605
rect 1283 1536 1289 1570
rect 1323 1566 1428 1570
rect 1323 1536 1388 1566
rect 1283 1532 1388 1536
rect 1422 1532 1428 1566
rect 1283 1496 1428 1532
rect 1283 1462 1289 1496
rect 1323 1493 1428 1496
rect 1323 1462 1388 1493
rect 1283 1459 1388 1462
rect 1422 1459 1428 1493
rect 1283 1421 1428 1459
rect 1283 1387 1289 1421
rect 1323 1420 1428 1421
rect 1323 1387 1388 1420
rect 1283 1386 1388 1387
rect 1422 1386 1428 1420
rect 1283 1347 1428 1386
rect 1283 1346 1388 1347
rect 1283 1312 1289 1346
rect 1323 1313 1388 1346
rect 1422 1313 1428 1347
rect 1323 1312 1428 1313
rect 1283 1274 1428 1312
rect 1283 1271 1388 1274
rect 1283 1237 1289 1271
rect 1323 1240 1388 1271
rect 1422 1240 1428 1274
rect 1323 1237 1428 1240
rect 1283 1201 1428 1237
rect 1283 1196 1388 1201
rect 1283 1162 1289 1196
rect 1323 1167 1388 1196
rect 1422 1167 1428 1201
rect 1323 1162 1428 1167
rect 1283 1128 1428 1162
rect 1283 1121 1388 1128
rect 1283 1087 1289 1121
rect 1323 1094 1388 1121
rect 1422 1094 1428 1128
rect 1323 1087 1428 1094
rect 1283 1055 1428 1087
rect 1283 1046 1388 1055
rect 1283 1012 1289 1046
rect 1323 1021 1388 1046
rect 1422 1021 1428 1055
rect 1323 1012 1428 1021
rect 1283 982 1428 1012
rect 1283 971 1388 982
rect 1283 937 1289 971
rect 1323 948 1388 971
rect 1422 948 1428 982
rect 1323 937 1428 948
rect 1283 909 1428 937
rect 1283 896 1388 909
rect 1283 862 1289 896
rect 1323 875 1388 896
rect 1422 875 1428 909
rect 1323 862 1428 875
rect 1283 836 1428 862
rect 1283 821 1388 836
rect 1283 787 1289 821
rect 1323 802 1388 821
rect 1422 802 1428 836
rect 1323 787 1428 802
rect 1283 763 1428 787
rect 1283 746 1388 763
rect 1283 712 1289 746
rect 1323 729 1388 746
rect 1422 729 1428 763
rect 1323 712 1428 729
rect 1283 690 1428 712
rect 1283 671 1388 690
rect 1283 637 1289 671
rect 1323 656 1388 671
rect 1422 656 1428 690
rect 1323 644 1428 656
tri 1468 3837 1498 3867 se
rect 1498 3837 1582 3867
tri 1582 3837 1612 3867 nw
tri 7274 3856 7285 3867 ne
rect 7285 3856 11514 3867
tri 11266 3837 11285 3856 ne
rect 11285 3837 11514 3856
rect 1468 3836 1581 3837
tri 1581 3836 1582 3837 nw
tri 11285 3836 11286 3837 ne
rect 11286 3836 11514 3837
rect 1323 637 1334 644
rect 1283 615 1334 637
tri 1334 615 1363 644 nw
rect 1283 613 1332 615
tri 1332 613 1334 615 nw
rect 1283 596 1329 613
tri 1329 610 1332 613 nw
rect 1283 562 1289 596
rect 1323 562 1329 596
rect 1283 521 1329 562
rect 1283 487 1289 521
rect 1323 487 1329 521
rect 1283 446 1329 487
rect 1283 412 1289 446
rect 1323 412 1329 446
tri 1466 433 1468 435 se
rect 1468 433 1548 3836
tri 1548 3803 1581 3836 nw
tri 11286 3803 11319 3836 ne
rect 11319 3803 11514 3836
tri 11319 3802 11320 3803 ne
rect 11320 3802 11514 3803
tri 11320 3739 11383 3802 ne
rect 11383 3739 11514 3802
tri 11383 3738 11384 3739 ne
tri 1463 430 1466 433 se
rect 1466 430 1548 433
rect 1283 400 1329 412
tri 1433 400 1463 430 se
rect 1463 400 1548 430
tri 1429 396 1433 400 se
rect 1433 396 1548 400
tri 1428 395 1429 396 se
rect 1429 395 1548 396
tri 1427 394 1428 395 se
rect 1428 394 1548 395
tri 1395 362 1427 394 se
rect 1427 362 1548 394
rect 411 356 1548 362
rect 411 322 426 356
rect 460 322 500 356
rect 534 322 574 356
rect 608 322 648 356
rect 682 322 721 356
rect 755 322 794 356
rect 828 322 867 356
rect 901 322 940 356
rect 974 322 1013 356
rect 1047 322 1086 356
rect 1120 322 1159 356
rect 1193 322 1232 356
rect 1266 322 1548 356
rect 411 273 1548 322
rect 1671 3666 11313 3670
rect 1671 3664 4820 3666
rect 4872 3664 4885 3666
rect 1671 3630 1749 3664
rect 1783 3630 1822 3664
rect 1856 3630 1895 3664
rect 1929 3630 1968 3664
rect 2002 3630 2041 3664
rect 2075 3630 2113 3664
rect 2147 3630 2185 3664
rect 2219 3630 2257 3664
rect 2291 3630 2329 3664
rect 2363 3630 2401 3664
rect 2435 3630 2473 3664
rect 2507 3630 2545 3664
rect 2579 3630 2617 3664
rect 2651 3630 2689 3664
rect 2723 3630 2761 3664
rect 2795 3630 2833 3664
rect 2867 3630 2905 3664
rect 2939 3630 2977 3664
rect 3011 3630 3049 3664
rect 3083 3630 3121 3664
rect 3155 3630 3193 3664
rect 3227 3630 3265 3664
rect 3299 3630 3432 3664
rect 3466 3630 3505 3664
rect 3539 3630 3578 3664
rect 3612 3630 3651 3664
rect 3685 3630 3724 3664
rect 3758 3630 3797 3664
rect 3831 3630 3870 3664
rect 3904 3630 3942 3664
rect 3976 3630 4014 3664
rect 4048 3630 4086 3664
rect 4120 3630 4158 3664
rect 4192 3630 4230 3664
rect 4264 3630 4302 3664
rect 4336 3630 4374 3664
rect 4408 3630 4446 3664
rect 4480 3630 4518 3664
rect 4552 3630 4590 3664
rect 4624 3630 4662 3664
rect 4696 3630 4734 3664
rect 4768 3630 4806 3664
rect 4872 3630 4878 3664
rect 1671 3614 4820 3630
rect 4872 3614 4885 3630
rect 4937 3614 4950 3666
rect 5002 3614 5015 3666
rect 5067 3614 5080 3666
rect 5132 3614 5145 3666
rect 5197 3664 5210 3666
rect 5262 3664 5275 3666
rect 5327 3664 5340 3666
rect 5392 3664 5405 3666
rect 5457 3664 5470 3666
rect 5522 3664 5535 3666
rect 5587 3664 5600 3666
rect 5200 3630 5210 3664
rect 5272 3630 5275 3664
rect 5522 3630 5526 3664
rect 5587 3630 5598 3664
rect 5197 3614 5210 3630
rect 5262 3614 5275 3630
rect 5327 3614 5340 3630
rect 5392 3614 5405 3630
rect 5457 3614 5470 3630
rect 5522 3614 5535 3630
rect 5587 3614 5600 3630
rect 5652 3614 5665 3666
rect 5717 3614 5730 3666
rect 5782 3614 5795 3666
rect 5847 3664 5860 3666
rect 5912 3664 5925 3666
rect 5977 3664 5990 3666
rect 6042 3664 6055 3666
rect 6107 3664 6120 3666
rect 6172 3664 6185 3666
rect 6237 3664 6250 3666
rect 5848 3630 5860 3664
rect 5920 3630 5925 3664
rect 6172 3630 6174 3664
rect 6237 3630 6246 3664
rect 5847 3614 5860 3630
rect 5912 3614 5925 3630
rect 5977 3614 5990 3630
rect 6042 3614 6055 3630
rect 6107 3614 6120 3630
rect 6172 3614 6185 3630
rect 6237 3614 6250 3630
rect 6302 3614 6315 3666
rect 6367 3614 6380 3666
rect 6432 3614 6445 3666
rect 6497 3614 6510 3666
rect 6562 3664 6575 3666
rect 6627 3664 6640 3666
rect 6692 3664 6705 3666
rect 6757 3664 6770 3666
rect 6822 3664 6835 3666
rect 6887 3664 6900 3666
rect 6568 3630 6575 3664
rect 6887 3630 6894 3664
rect 6562 3614 6575 3630
rect 6627 3614 6640 3630
rect 6692 3614 6705 3630
rect 6757 3614 6770 3630
rect 6822 3614 6835 3630
rect 6887 3614 6900 3630
rect 6952 3614 6965 3666
rect 7017 3614 7030 3666
rect 7082 3614 7095 3666
rect 7147 3614 7160 3666
rect 7212 3664 7225 3666
rect 7216 3630 7225 3664
rect 7212 3614 7225 3630
rect 7277 3614 7290 3666
rect 7342 3614 7355 3666
rect 7407 3614 7419 3666
rect 7471 3614 7483 3666
rect 7535 3614 7547 3666
rect 7599 3664 7611 3666
rect 7663 3664 7675 3666
rect 7727 3664 7739 3666
rect 7791 3664 7803 3666
rect 7855 3664 7867 3666
rect 7608 3630 7611 3664
rect 7855 3630 7862 3664
rect 7599 3614 7611 3630
rect 7663 3614 7675 3630
rect 7727 3614 7739 3630
rect 7791 3614 7803 3630
rect 7855 3614 7867 3630
rect 7919 3614 7931 3666
rect 7983 3614 7995 3666
rect 8047 3614 8059 3666
rect 8111 3664 8123 3666
rect 8175 3664 8187 3666
rect 8239 3664 8251 3666
rect 8303 3664 8315 3666
rect 8367 3664 8379 3666
rect 8431 3664 8443 3666
rect 8112 3630 8123 3664
rect 8184 3630 8187 3664
rect 8431 3630 8438 3664
rect 8111 3614 8123 3630
rect 8175 3614 8187 3630
rect 8239 3614 8251 3630
rect 8303 3614 8315 3630
rect 8367 3614 8379 3630
rect 8431 3614 8443 3630
rect 8495 3614 8507 3666
rect 8559 3614 8571 3666
rect 8623 3614 8635 3666
rect 8687 3664 8699 3666
rect 8751 3664 8763 3666
rect 8815 3664 8827 3666
rect 8879 3664 8891 3666
rect 8943 3664 8955 3666
rect 9007 3664 9019 3666
rect 8688 3630 8699 3664
rect 8760 3630 8763 3664
rect 9007 3630 9014 3664
rect 8687 3614 8699 3630
rect 8751 3614 8763 3630
rect 8815 3614 8827 3630
rect 8879 3614 8891 3630
rect 8943 3614 8955 3630
rect 9007 3614 9019 3630
rect 9071 3614 9083 3666
rect 9135 3614 9147 3666
rect 9199 3614 9211 3666
rect 9263 3664 9275 3666
rect 9327 3664 9339 3666
rect 9391 3664 9403 3666
rect 9455 3664 9467 3666
rect 9519 3664 9531 3666
rect 9583 3664 9595 3666
rect 9264 3630 9275 3664
rect 9336 3630 9339 3664
rect 9583 3630 9590 3664
rect 9263 3614 9275 3630
rect 9327 3614 9339 3630
rect 9391 3614 9403 3630
rect 9455 3614 9467 3630
rect 9519 3614 9531 3630
rect 9583 3614 9595 3630
rect 9647 3614 9659 3666
rect 9711 3614 9723 3666
rect 9775 3614 9787 3666
rect 9839 3664 9851 3666
rect 9903 3664 9915 3666
rect 9967 3664 9979 3666
rect 10031 3664 10043 3666
rect 10095 3664 10107 3666
rect 10159 3664 10171 3666
rect 9840 3630 9851 3664
rect 9912 3630 9915 3664
rect 10159 3630 10166 3664
rect 9839 3614 9851 3630
rect 9903 3614 9915 3630
rect 9967 3614 9979 3630
rect 10031 3614 10043 3630
rect 10095 3614 10107 3630
rect 10159 3614 10171 3630
rect 10223 3614 10235 3666
rect 10287 3614 10299 3666
rect 10351 3614 10363 3666
rect 10415 3664 10427 3666
rect 10479 3664 10491 3666
rect 10543 3664 10555 3666
rect 10607 3664 10619 3666
rect 10671 3664 10683 3666
rect 10735 3664 10747 3666
rect 10416 3630 10427 3664
rect 10488 3630 10491 3664
rect 10735 3630 10742 3664
rect 10415 3614 10427 3630
rect 10479 3614 10491 3630
rect 10543 3614 10555 3630
rect 10607 3614 10619 3630
rect 10671 3614 10683 3630
rect 10735 3614 10747 3630
rect 10799 3614 10811 3666
rect 10863 3664 11313 3666
rect 10863 3630 10886 3664
rect 10920 3630 10958 3664
rect 10992 3630 11030 3664
rect 11064 3630 11102 3664
rect 11136 3630 11174 3664
rect 11208 3630 11313 3664
rect 10863 3614 11313 3630
rect 1671 3592 11313 3614
rect 1671 3558 1677 3592
rect 1711 3578 11313 3592
rect 1711 3558 4820 3578
rect 1671 3556 4820 3558
rect 4872 3556 4885 3578
rect 1671 3522 1785 3556
rect 1819 3522 1859 3556
rect 1893 3522 1933 3556
rect 1967 3522 2007 3556
rect 2041 3522 2081 3556
rect 2115 3522 2155 3556
rect 2189 3522 2229 3556
rect 2263 3522 2303 3556
rect 2337 3522 2377 3556
rect 2411 3522 2451 3556
rect 2485 3522 2525 3556
rect 2559 3522 2599 3556
rect 2633 3522 2673 3556
rect 2707 3522 2747 3556
rect 2781 3522 2821 3556
rect 2855 3522 2895 3556
rect 2929 3522 2969 3556
rect 3003 3522 3043 3556
rect 3077 3522 3117 3556
rect 3151 3522 3191 3556
rect 3225 3522 3265 3556
rect 3299 3542 3432 3556
rect 3299 3522 3331 3542
rect 1671 3520 3331 3522
rect 1671 3486 1677 3520
rect 1711 3486 3331 3520
rect 3400 3522 3432 3542
rect 3466 3522 3505 3556
rect 3539 3522 3578 3556
rect 3612 3522 3651 3556
rect 3685 3522 3724 3556
rect 3758 3522 3797 3556
rect 3831 3522 3870 3556
rect 3904 3522 3942 3556
rect 3976 3522 4014 3556
rect 4048 3522 4086 3556
rect 4120 3522 4158 3556
rect 4192 3522 4230 3556
rect 4264 3522 4302 3556
rect 4336 3522 4374 3556
rect 4408 3522 4446 3556
rect 4480 3522 4518 3556
rect 4552 3522 4590 3556
rect 4624 3522 4662 3556
rect 4696 3522 4734 3556
rect 4768 3522 4806 3556
rect 4872 3526 4878 3556
rect 4937 3526 4950 3578
rect 5002 3526 5015 3578
rect 5067 3526 5080 3578
rect 5132 3526 5145 3578
rect 5197 3556 5210 3578
rect 5262 3556 5275 3578
rect 5327 3556 5340 3578
rect 5392 3556 5405 3578
rect 5457 3556 5470 3578
rect 5522 3556 5535 3578
rect 5587 3556 5600 3578
rect 5200 3526 5210 3556
rect 5272 3526 5275 3556
rect 5522 3526 5526 3556
rect 5587 3526 5598 3556
rect 5652 3526 5665 3578
rect 5717 3526 5730 3578
rect 5782 3526 5795 3578
rect 5847 3556 5860 3578
rect 5912 3556 5925 3578
rect 5977 3556 5990 3578
rect 6042 3556 6055 3578
rect 6107 3556 6120 3578
rect 6172 3556 6185 3578
rect 6237 3556 6250 3578
rect 5848 3526 5860 3556
rect 5920 3526 5925 3556
rect 6172 3526 6174 3556
rect 6237 3526 6246 3556
rect 6302 3526 6315 3578
rect 6367 3526 6380 3578
rect 6432 3526 6445 3578
rect 6497 3526 6510 3578
rect 6562 3556 6575 3578
rect 6627 3556 6640 3578
rect 6692 3556 6705 3578
rect 6757 3556 6770 3578
rect 6822 3556 6835 3578
rect 6887 3556 6900 3578
rect 6568 3526 6575 3556
rect 6887 3526 6894 3556
rect 6952 3526 6965 3578
rect 7017 3526 7030 3578
rect 7082 3526 7095 3578
rect 7147 3526 7160 3578
rect 7212 3556 7225 3578
rect 7216 3526 7225 3556
rect 7277 3526 7290 3578
rect 7342 3526 7355 3578
rect 7407 3526 7419 3578
rect 7471 3526 7483 3578
rect 7535 3526 7547 3578
rect 7599 3556 7611 3578
rect 7663 3556 7675 3578
rect 7727 3556 7739 3578
rect 7791 3556 7803 3578
rect 7855 3556 7867 3578
rect 7608 3526 7611 3556
rect 7855 3526 7862 3556
rect 7919 3526 7931 3578
rect 7983 3526 7995 3578
rect 8047 3526 8059 3578
rect 8111 3556 8123 3578
rect 8175 3556 8187 3578
rect 8239 3556 8251 3578
rect 8303 3556 8315 3578
rect 8367 3556 8379 3578
rect 8431 3556 8443 3578
rect 8112 3526 8123 3556
rect 8184 3526 8187 3556
rect 8431 3526 8438 3556
rect 8495 3526 8507 3578
rect 8559 3526 8571 3578
rect 8623 3526 8635 3578
rect 8687 3556 8699 3578
rect 8751 3556 8763 3578
rect 8815 3556 8827 3578
rect 8879 3556 8891 3578
rect 8943 3556 8955 3578
rect 9007 3556 9019 3578
rect 8688 3526 8699 3556
rect 8760 3526 8763 3556
rect 9007 3526 9014 3556
rect 9071 3526 9083 3578
rect 9135 3526 9147 3578
rect 9199 3526 9211 3578
rect 9263 3556 9275 3578
rect 9327 3556 9339 3578
rect 9391 3556 9403 3578
rect 9455 3556 9467 3578
rect 9519 3556 9531 3578
rect 9583 3556 9595 3578
rect 9264 3526 9275 3556
rect 9336 3526 9339 3556
rect 9583 3526 9590 3556
rect 9647 3526 9659 3578
rect 9711 3526 9723 3578
rect 9775 3526 9787 3578
rect 9839 3556 9851 3578
rect 9903 3556 9915 3578
rect 9967 3556 9979 3578
rect 10031 3556 10043 3578
rect 10095 3556 10107 3578
rect 10159 3556 10171 3578
rect 9840 3526 9851 3556
rect 9912 3526 9915 3556
rect 10159 3526 10166 3556
rect 10223 3526 10235 3578
rect 10287 3526 10299 3578
rect 10351 3526 10363 3578
rect 10415 3556 10427 3578
rect 10479 3556 10491 3578
rect 10543 3556 10555 3578
rect 10607 3556 10619 3578
rect 10671 3556 10683 3578
rect 10735 3556 10747 3578
rect 10416 3526 10427 3556
rect 10488 3526 10491 3556
rect 10735 3526 10742 3556
rect 10799 3526 10811 3578
rect 10863 3556 11313 3578
rect 10863 3526 10886 3556
rect 4840 3522 4878 3526
rect 4912 3522 4950 3526
rect 4984 3522 5022 3526
rect 5056 3522 5094 3526
rect 5128 3522 5166 3526
rect 5200 3522 5238 3526
rect 5272 3522 5310 3526
rect 5344 3522 5382 3526
rect 5416 3522 5454 3526
rect 5488 3522 5526 3526
rect 5560 3522 5598 3526
rect 5632 3522 5670 3526
rect 5704 3522 5742 3526
rect 5776 3522 5814 3526
rect 5848 3522 5886 3526
rect 5920 3522 5958 3526
rect 5992 3522 6030 3526
rect 6064 3522 6102 3526
rect 6136 3522 6174 3526
rect 6208 3522 6246 3526
rect 6280 3522 6318 3526
rect 6352 3522 6390 3526
rect 6424 3522 6462 3526
rect 6496 3522 6534 3526
rect 6568 3522 6606 3526
rect 6640 3522 6678 3526
rect 6712 3522 6750 3526
rect 6784 3522 6822 3526
rect 6856 3522 6894 3526
rect 6928 3522 6966 3526
rect 7000 3522 7038 3526
rect 7072 3522 7110 3526
rect 7144 3522 7182 3526
rect 7216 3522 7428 3526
rect 7462 3522 7501 3526
rect 7535 3522 7574 3526
rect 7608 3522 7646 3526
rect 7680 3522 7718 3526
rect 7752 3522 7790 3526
rect 7824 3522 7862 3526
rect 7896 3522 7934 3526
rect 7968 3522 8006 3526
rect 8040 3522 8078 3526
rect 8112 3522 8150 3526
rect 8184 3522 8222 3526
rect 8256 3522 8294 3526
rect 8328 3522 8366 3526
rect 8400 3522 8438 3526
rect 8472 3522 8510 3526
rect 8544 3522 8582 3526
rect 8616 3522 8654 3526
rect 8688 3522 8726 3526
rect 8760 3522 8798 3526
rect 8832 3522 8870 3526
rect 8904 3522 8942 3526
rect 8976 3522 9014 3526
rect 9048 3522 9086 3526
rect 9120 3522 9158 3526
rect 9192 3522 9230 3526
rect 9264 3522 9302 3526
rect 9336 3522 9374 3526
rect 9408 3522 9446 3526
rect 9480 3522 9518 3526
rect 9552 3522 9590 3526
rect 9624 3522 9662 3526
rect 9696 3522 9734 3526
rect 9768 3522 9806 3526
rect 9840 3522 9878 3526
rect 9912 3522 9950 3526
rect 9984 3522 10022 3526
rect 10056 3522 10094 3526
rect 10128 3522 10166 3526
rect 10200 3522 10238 3526
rect 10272 3522 10310 3526
rect 10344 3522 10382 3526
rect 10416 3522 10454 3526
rect 10488 3522 10526 3526
rect 10560 3522 10598 3526
rect 10632 3522 10670 3526
rect 10704 3522 10742 3526
rect 10776 3522 10814 3526
rect 10848 3522 10886 3526
rect 10920 3522 10958 3556
rect 10992 3522 11030 3556
rect 11064 3522 11102 3556
rect 11136 3522 11174 3556
rect 11208 3542 11313 3556
rect 11208 3522 11240 3542
rect 3400 3516 11240 3522
rect 1671 3484 3331 3486
rect 1671 3450 1785 3484
rect 1819 3461 3331 3484
tri 3413 3466 3463 3516 nw
tri 7185 3482 7219 3516 ne
rect 7219 3482 7233 3516
tri 7219 3468 7233 3482 ne
rect 7411 3482 7425 3516
tri 7425 3482 7459 3516 nw
tri 11197 3482 11231 3516 ne
tri 7411 3468 7425 3482 nw
rect 1819 3450 1892 3461
rect 1671 3448 1892 3450
rect 1671 3414 1677 3448
rect 1711 3427 1892 3448
rect 1926 3427 1967 3461
rect 2001 3427 2042 3461
rect 2076 3427 2117 3461
rect 2151 3427 2192 3461
rect 2226 3427 2266 3461
rect 2300 3427 2340 3461
rect 2374 3427 2414 3461
rect 2448 3427 2488 3461
rect 2522 3427 2562 3461
rect 2596 3427 2636 3461
rect 2670 3427 2710 3461
rect 2744 3427 2784 3461
rect 2818 3427 2858 3461
rect 2892 3427 2932 3461
rect 2966 3427 3006 3461
rect 3040 3427 3080 3461
rect 3114 3427 3154 3461
rect 3188 3427 3228 3461
rect 3262 3427 3331 3461
rect 1711 3414 3331 3427
rect 1671 3412 3331 3414
rect 1671 3378 1785 3412
rect 1819 3389 3331 3412
rect 1819 3378 1892 3389
rect 1671 3376 1892 3378
rect 1671 3342 1677 3376
rect 1711 3355 1892 3376
rect 1926 3355 1967 3389
rect 2001 3355 2042 3389
rect 2076 3355 2117 3389
rect 2151 3355 2192 3389
rect 2226 3355 2266 3389
rect 2300 3355 2340 3389
rect 2374 3355 2414 3389
rect 2448 3355 2488 3389
rect 2522 3355 2562 3389
rect 2596 3355 2636 3389
rect 2670 3355 2710 3389
rect 2744 3355 2784 3389
rect 2818 3355 2858 3389
rect 2892 3355 2932 3389
rect 2966 3355 3006 3389
rect 3040 3355 3080 3389
rect 3114 3355 3154 3389
rect 3188 3355 3228 3389
rect 3262 3355 3331 3389
rect 1711 3342 3331 3355
rect 1671 3340 3331 3342
rect 1671 3306 1785 3340
rect 1819 3317 3331 3340
rect 1819 3306 1892 3317
rect 1671 3304 1892 3306
rect 1671 3270 1677 3304
rect 1711 3283 1892 3304
rect 1926 3283 1967 3317
rect 2001 3283 2042 3317
rect 2076 3283 2117 3317
rect 2151 3283 2192 3317
rect 2226 3283 2266 3317
rect 2300 3283 2340 3317
rect 2374 3283 2414 3317
rect 2448 3283 2488 3317
rect 2522 3283 2562 3317
rect 2596 3283 2636 3317
rect 2670 3283 2710 3317
rect 2744 3283 2784 3317
rect 2818 3283 2858 3317
rect 2892 3283 2932 3317
rect 2966 3283 3006 3317
rect 3040 3283 3080 3317
rect 3114 3283 3154 3317
rect 3188 3283 3228 3317
rect 3262 3283 3331 3317
rect 1711 3270 3331 3283
rect 1671 3268 3331 3270
rect 1671 3234 1785 3268
rect 1819 3245 3331 3268
rect 1819 3234 1892 3245
rect 1671 3232 1892 3234
rect 1671 3198 1677 3232
rect 1711 3211 1892 3232
rect 1926 3211 1967 3245
rect 2001 3211 2042 3245
rect 2076 3211 2117 3245
rect 2151 3211 2192 3245
rect 2226 3211 2266 3245
rect 2300 3211 2340 3245
rect 2374 3211 2414 3245
rect 2448 3211 2488 3245
rect 2522 3211 2562 3245
rect 2596 3211 2636 3245
rect 2670 3211 2710 3245
rect 2744 3211 2784 3245
rect 2818 3211 2858 3245
rect 2892 3211 2932 3245
rect 2966 3211 3006 3245
rect 3040 3211 3080 3245
rect 3114 3211 3154 3245
rect 3188 3211 3228 3245
rect 3262 3211 3331 3245
rect 1711 3198 3331 3211
rect 1671 3196 3331 3198
rect 1671 3162 1785 3196
rect 1819 3173 3331 3196
rect 1819 3162 1892 3173
rect 1671 3160 1892 3162
rect 1671 3126 1677 3160
rect 1711 3139 1892 3160
rect 1926 3139 1967 3173
rect 2001 3139 2042 3173
rect 2076 3139 2117 3173
rect 2151 3139 2192 3173
rect 2226 3139 2266 3173
rect 2300 3139 2340 3173
rect 2374 3139 2414 3173
rect 2448 3139 2488 3173
rect 2522 3139 2562 3173
rect 2596 3139 2636 3173
rect 2670 3139 2710 3173
rect 2744 3139 2784 3173
rect 2818 3139 2858 3173
rect 2892 3139 2932 3173
rect 2966 3139 3006 3173
rect 3040 3139 3080 3173
rect 3114 3139 3154 3173
rect 3188 3139 3228 3173
rect 3262 3139 3331 3173
rect 1711 3133 3331 3139
rect 1711 3129 1891 3133
tri 1891 3129 1895 3133 nw
tri 3274 3129 3278 3133 ne
rect 3278 3129 3331 3133
rect 1711 3126 1874 3129
rect 1671 3124 1874 3126
rect 1671 3090 1785 3124
rect 1819 3112 1874 3124
tri 1874 3112 1891 3129 nw
tri 3278 3112 3295 3129 ne
rect 3295 3112 3331 3129
rect 1819 3090 1852 3112
tri 1852 3090 1874 3112 nw
tri 3295 3090 3317 3112 ne
rect 3317 3090 3331 3112
rect 1671 3088 1825 3090
rect 1671 3054 1677 3088
rect 1711 3054 1825 3088
tri 1825 3063 1852 3090 nw
tri 3317 3076 3331 3090 ne
rect 3937 3410 4237 3416
rect 3937 3358 3938 3410
rect 3990 3358 4020 3410
rect 4072 3358 4102 3410
rect 4154 3358 4184 3410
rect 4236 3358 4237 3410
rect 3937 3344 4237 3358
rect 3937 3292 3938 3344
rect 3990 3292 4020 3344
rect 4072 3292 4102 3344
rect 4154 3292 4184 3344
rect 4236 3292 4237 3344
rect 3937 3278 4237 3292
rect 3937 3226 3938 3278
rect 3990 3226 4020 3278
rect 4072 3226 4102 3278
rect 4154 3226 4184 3278
rect 4236 3226 4237 3278
rect 3937 3212 4237 3226
rect 3937 3160 3938 3212
rect 3990 3160 4020 3212
rect 4072 3160 4102 3212
rect 4154 3160 4184 3212
rect 4236 3160 4237 3212
rect 3937 3146 4237 3160
rect 3937 3094 3938 3146
rect 3990 3094 4020 3146
rect 4072 3094 4102 3146
rect 4154 3094 4184 3146
rect 4236 3094 4237 3146
rect 3937 3079 4237 3094
rect 1671 3052 1825 3054
rect 1671 3018 1785 3052
rect 1819 3018 1825 3052
rect 1671 3016 1825 3018
rect 1671 2982 1677 3016
rect 1711 2982 1825 3016
rect 1671 2980 1825 2982
rect 1671 2946 1785 2980
rect 1819 2946 1825 2980
rect 1671 2944 1825 2946
rect 1671 2910 1677 2944
rect 1711 2910 1825 2944
rect 1671 2908 1825 2910
rect 1671 2874 1785 2908
rect 1819 2874 1825 2908
rect 1671 2872 1825 2874
rect 1671 2838 1677 2872
rect 1711 2838 1825 2872
rect 1671 2836 1825 2838
rect 1671 2802 1785 2836
rect 1819 2802 1825 2836
rect 1671 2800 1825 2802
rect 1671 2766 1677 2800
rect 1711 2766 1825 2800
rect 1671 2764 1825 2766
rect 1671 2730 1785 2764
rect 1819 2730 1825 2764
rect 1671 2728 1825 2730
rect 1671 2694 1677 2728
rect 1711 2694 1825 2728
rect 1671 2692 1825 2694
rect 1671 2658 1785 2692
rect 1819 2658 1825 2692
rect 1671 2656 1825 2658
rect 1671 2622 1677 2656
rect 1711 2622 1825 2656
rect 1671 2620 1825 2622
rect 1671 2586 1785 2620
rect 1819 2586 1825 2620
rect 1671 2584 1825 2586
rect 1671 2550 1677 2584
rect 1711 2550 1825 2584
rect 1671 2547 1825 2550
rect 1671 2513 1785 2547
rect 1819 2513 1825 2547
rect 1671 2511 1825 2513
rect 1671 2477 1677 2511
rect 1711 2477 1825 2511
rect 1671 2474 1825 2477
rect 1671 2440 1785 2474
rect 1819 2440 1825 2474
rect 1671 2438 1825 2440
rect 1671 2404 1677 2438
rect 1711 2404 1825 2438
rect 1671 2401 1825 2404
rect 1671 2367 1785 2401
rect 1819 2367 1825 2401
rect 1671 2365 1825 2367
rect 1671 2331 1677 2365
rect 1711 2331 1825 2365
rect 1671 2328 1825 2331
rect 1671 2294 1785 2328
rect 1819 2294 1825 2328
rect 1671 2292 1825 2294
rect 1671 2258 1677 2292
rect 1711 2258 1825 2292
rect 1671 2255 1825 2258
rect 1671 2221 1785 2255
rect 1819 2221 1825 2255
rect 1671 2219 1825 2221
rect 1671 2185 1677 2219
rect 1711 2185 1825 2219
rect 1671 2182 1825 2185
rect 1671 2148 1785 2182
rect 1819 2148 1825 2182
rect 1671 2146 1825 2148
rect 1671 2112 1677 2146
rect 1711 2112 1825 2146
rect 1671 2109 1825 2112
rect 1671 2075 1785 2109
rect 1819 2075 1825 2109
rect 1671 2073 1825 2075
rect 1671 2039 1677 2073
rect 1711 2039 1825 2073
rect 1671 2036 1825 2039
rect 1671 2002 1785 2036
rect 1819 2002 1825 2036
rect 1671 2000 1825 2002
rect 1671 1966 1677 2000
rect 1711 1966 1825 2000
rect 1671 1963 1825 1966
rect 1671 1929 1785 1963
rect 1819 1929 1825 1963
rect 1671 1927 1825 1929
rect 1671 1893 1677 1927
rect 1711 1893 1825 1927
rect 1671 1890 1825 1893
rect 1671 1856 1785 1890
rect 1819 1856 1825 1890
rect 1671 1854 1825 1856
rect 1671 1820 1677 1854
rect 1711 1820 1825 1854
rect 1671 1817 1825 1820
rect 1671 1783 1785 1817
rect 1819 1783 1825 1817
rect 1671 1781 1825 1783
rect 1671 1747 1677 1781
rect 1711 1747 1825 1781
rect 1671 1744 1825 1747
rect 1671 1710 1785 1744
rect 1819 1710 1825 1744
rect 1671 1708 1825 1710
rect 1671 1674 1677 1708
rect 1711 1674 1825 1708
rect 1671 1671 1825 1674
rect 1671 1637 1785 1671
rect 1819 1637 1825 1671
rect 1671 1635 1825 1637
rect 1671 1601 1677 1635
rect 1711 1601 1825 1635
rect 1671 1598 1825 1601
rect 1671 1564 1785 1598
rect 1819 1564 1825 1598
rect 1671 1562 1825 1564
rect 1671 1528 1677 1562
rect 1711 1528 1825 1562
rect 1671 1525 1825 1528
rect 1671 1491 1785 1525
rect 1819 1491 1825 1525
rect 1671 1489 1825 1491
rect 1671 1455 1677 1489
rect 1711 1455 1825 1489
rect 1671 1452 1825 1455
rect 1671 1418 1785 1452
rect 1819 1418 1825 1452
rect 1671 1416 1825 1418
rect 1671 1382 1677 1416
rect 1711 1382 1825 1416
rect 1671 1379 1825 1382
rect 1671 1345 1785 1379
rect 1819 1345 1825 1379
rect 1671 1343 1825 1345
rect 1671 1309 1677 1343
rect 1711 1309 1825 1343
rect 1671 1306 1825 1309
rect 1671 1272 1785 1306
rect 1819 1272 1825 1306
rect 1671 1270 1825 1272
rect 1671 1236 1677 1270
rect 1711 1236 1825 1270
rect 1671 1233 1825 1236
rect 1671 1199 1785 1233
rect 1819 1199 1825 1233
rect 1671 1197 1825 1199
rect 1671 1163 1677 1197
rect 1711 1163 1825 1197
rect 1671 1160 1825 1163
rect 1671 1126 1785 1160
rect 1819 1126 1825 1160
rect 1671 1124 1825 1126
rect 1671 1090 1677 1124
rect 1711 1090 1825 1124
rect 1671 1087 1825 1090
rect 1671 1053 1785 1087
rect 1819 1053 1825 1087
rect 1671 1051 1825 1053
rect 1671 1017 1677 1051
rect 1711 1017 1825 1051
rect 1671 1014 1825 1017
rect 1671 980 1785 1014
rect 1819 980 1825 1014
rect 1671 978 1825 980
rect 1671 944 1677 978
rect 1711 944 1825 978
rect 1671 941 1825 944
rect 1671 907 1785 941
rect 1819 907 1825 941
rect 1671 905 1825 907
rect 1671 871 1677 905
rect 1711 871 1825 905
rect 1671 868 1825 871
rect 1671 834 1785 868
rect 1819 834 1825 868
rect 1671 832 1825 834
rect 1671 798 1677 832
rect 1711 798 1825 832
rect 1671 795 1825 798
rect 1671 761 1785 795
rect 1819 761 1825 795
rect 1671 759 1825 761
rect 1671 725 1677 759
rect 1711 725 1825 759
rect 1671 722 1825 725
rect 1671 688 1785 722
rect 1819 688 1825 722
rect 1671 686 1825 688
rect 1671 652 1677 686
rect 1711 656 1825 686
rect 1933 2862 1939 3042
rect 2119 2990 2132 3042
rect 2184 2990 2197 3042
rect 2249 2990 2262 3042
rect 2314 2990 2327 3042
rect 2379 2990 2392 3042
rect 2444 2990 2457 3042
rect 2509 2990 2522 3042
rect 2574 2990 2587 3042
rect 2639 2990 2652 3042
rect 2704 2990 2717 3042
rect 2769 2990 2782 3042
rect 2834 2990 2847 3042
rect 2899 2990 2912 3042
rect 2964 2990 2977 3042
rect 3029 2990 3042 3042
rect 3094 2990 3107 3042
rect 3159 2990 3223 3042
rect 2119 2978 3223 2990
rect 2119 2926 2132 2978
rect 2184 2926 2197 2978
rect 2249 2926 2262 2978
rect 2314 2926 2327 2978
rect 2379 2926 2392 2978
rect 2444 2926 2457 2978
rect 2509 2926 2522 2978
rect 2574 2926 2587 2978
rect 2639 2926 2652 2978
rect 2704 2926 2717 2978
rect 2769 2926 2782 2978
rect 2834 2926 2847 2978
rect 2899 2926 2912 2978
rect 2964 2926 2977 2978
rect 3029 2926 3042 2978
rect 3094 2926 3107 2978
rect 2055 2914 3107 2926
rect 2055 2862 2068 2914
rect 2120 2862 2133 2914
rect 2185 2862 2198 2914
rect 2250 2862 2263 2914
rect 2315 2862 2328 2914
rect 2380 2862 2393 2914
rect 2445 2862 2458 2914
rect 2510 2862 2523 2914
rect 2575 2862 2588 2914
rect 2640 2862 2653 2914
rect 2705 2862 2718 2914
rect 2770 2862 2783 2914
rect 2835 2862 2848 2914
rect 2900 2862 2913 2914
rect 2965 2862 2978 2914
rect 3030 2862 3043 2914
rect 1933 2850 3043 2862
rect 1933 2798 1939 2850
rect 1991 2798 2004 2850
rect 2056 2798 2069 2850
rect 2121 2798 2134 2850
rect 2186 2798 2199 2850
rect 2251 2798 2264 2850
rect 2316 2798 2329 2850
rect 2381 2798 2394 2850
rect 2446 2798 2459 2850
rect 2511 2798 2524 2850
rect 2576 2798 2589 2850
rect 2641 2798 2654 2850
rect 2706 2798 2719 2850
rect 2771 2798 2784 2850
rect 2836 2798 2849 2850
rect 2901 2798 2914 2850
rect 2966 2798 2979 2850
rect 1933 2786 2979 2798
rect 1933 2734 1939 2786
rect 1991 2734 2004 2786
rect 2056 2734 2069 2786
rect 2121 2734 2134 2786
rect 2186 2734 2199 2786
rect 2251 2734 2264 2786
rect 2316 2734 2329 2786
rect 2381 2734 2394 2786
rect 2446 2734 2459 2786
rect 2511 2734 2524 2786
rect 2576 2734 2589 2786
rect 2641 2734 2654 2786
rect 2706 2734 2719 2786
rect 2771 2734 2784 2786
rect 2836 2734 2849 2786
rect 2901 2734 2915 2786
rect 1933 2722 2915 2734
rect 1933 2670 1939 2722
rect 1991 2670 2004 2722
rect 2056 2670 2069 2722
rect 2121 2670 2134 2722
rect 2186 2670 2199 2722
rect 2251 2670 2264 2722
rect 2316 2670 2329 2722
rect 2381 2670 2394 2722
rect 2446 2670 2459 2722
rect 2511 2670 2524 2722
rect 2576 2670 2589 2722
rect 2641 2670 2654 2722
rect 2706 2670 2719 2722
rect 2771 2670 2785 2722
rect 2837 2670 2851 2722
rect 1933 2658 2851 2670
rect 1933 2606 1939 2658
rect 1991 2606 2004 2658
rect 2056 2606 2069 2658
rect 2121 2606 2134 2658
rect 2186 2606 2199 2658
rect 2251 2606 2264 2658
rect 2316 2606 2329 2658
rect 2381 2606 2394 2658
rect 2446 2606 2459 2658
rect 2511 2606 2524 2658
rect 2576 2606 2589 2658
rect 2641 2606 2655 2658
rect 2707 2606 2721 2658
rect 2773 2606 2787 2658
rect 1933 2594 2787 2606
rect 1933 2542 1939 2594
rect 1991 2542 2004 2594
rect 2056 2542 2069 2594
rect 2121 2542 2134 2594
rect 2186 2542 2199 2594
rect 2251 2542 2264 2594
rect 2316 2542 2329 2594
rect 2381 2542 2394 2594
rect 2446 2542 2459 2594
rect 2511 2542 2525 2594
rect 2577 2542 2591 2594
rect 2643 2542 2657 2594
rect 2709 2542 2723 2594
rect 1933 2530 2723 2542
rect 1933 2478 1939 2530
rect 1991 2478 2004 2530
rect 2056 2478 2069 2530
rect 2121 2478 2134 2530
rect 2186 2478 2199 2530
rect 2251 2478 2264 2530
rect 2316 2478 2329 2530
rect 2381 2478 2395 2530
rect 2447 2478 2461 2530
rect 2513 2478 2527 2530
rect 2579 2478 2593 2530
rect 2645 2478 2659 2530
rect 1933 2466 2659 2478
rect 1933 2414 1939 2466
rect 1991 2414 2004 2466
rect 2056 2414 2069 2466
rect 2121 2414 2134 2466
rect 2186 2414 2199 2466
rect 2251 2414 2265 2466
rect 2317 2414 2331 2466
rect 2383 2414 2397 2466
rect 2449 2414 2463 2466
rect 2515 2414 2529 2466
rect 2581 2414 2595 2466
rect 2647 2414 2659 2466
rect 1933 2402 2659 2414
rect 1933 2350 1939 2402
rect 1991 2350 2004 2402
rect 2056 2350 2069 2402
rect 2121 2350 2135 2402
rect 2187 2350 2201 2402
rect 2253 2350 2267 2402
rect 2319 2350 2333 2402
rect 2385 2350 2399 2402
rect 2451 2350 2465 2402
rect 2517 2350 2531 2402
rect 2583 2401 2659 2402
rect 2583 2350 2595 2401
rect 1933 2349 2595 2350
rect 2647 2350 2659 2401
rect 2647 2349 2723 2350
rect 1933 2338 2723 2349
rect 1933 2286 1939 2338
rect 1991 2286 2005 2338
rect 2057 2286 2071 2338
rect 2123 2286 2137 2338
rect 2189 2286 2203 2338
rect 2255 2286 2269 2338
rect 2321 2286 2335 2338
rect 2387 2286 2401 2338
rect 2453 2286 2467 2338
rect 2519 2337 2723 2338
rect 2519 2286 2531 2337
rect 1933 2285 2531 2286
rect 2583 2336 2659 2337
rect 2583 2285 2595 2336
rect 1933 2284 2595 2285
rect 2647 2285 2659 2336
rect 2711 2286 2723 2337
rect 2711 2285 2787 2286
rect 2647 2284 2787 2285
rect 1933 2274 2787 2284
rect 1933 2222 1939 2274
rect 1991 2222 2005 2274
rect 2057 2222 2071 2274
rect 2123 2222 2137 2274
rect 2189 2222 2203 2274
rect 2255 2222 2269 2274
rect 2321 2222 2336 2274
rect 2388 2222 2403 2274
rect 2455 2273 2787 2274
rect 2455 2222 2467 2273
rect 1933 2221 2467 2222
rect 2519 2272 2723 2273
rect 2519 2221 2531 2272
rect 1933 2220 2531 2221
rect 2583 2271 2659 2272
rect 2583 2220 2595 2271
rect 1933 2219 2595 2220
rect 2647 2220 2659 2271
rect 2711 2221 2723 2272
rect 2775 2222 2787 2273
rect 2775 2221 2851 2222
rect 2711 2220 2851 2221
rect 2647 2219 2851 2220
rect 1933 2209 2851 2219
rect 1933 2157 2403 2209
rect 2455 2208 2787 2209
rect 2455 2157 2467 2208
rect 1933 2156 2467 2157
rect 2519 2207 2723 2208
rect 2519 2156 2531 2207
rect 1933 2155 2531 2156
rect 2583 2206 2659 2207
rect 2583 2155 2595 2206
rect 1933 2154 2595 2155
rect 2647 2155 2659 2206
rect 2711 2156 2723 2207
rect 2775 2157 2787 2208
rect 2839 2158 2851 2209
rect 2839 2157 2915 2158
rect 2775 2156 2915 2157
rect 2711 2155 2915 2156
rect 2647 2154 2915 2155
rect 1933 2145 2915 2154
rect 1933 2144 2851 2145
rect 1933 2092 2403 2144
rect 2455 2143 2787 2144
rect 2455 2092 2467 2143
rect 1933 2091 2467 2092
rect 2519 2142 2723 2143
rect 2519 2091 2531 2142
rect 1933 2090 2531 2091
rect 2583 2141 2659 2142
rect 2583 2090 2595 2141
rect 1933 2089 2595 2090
rect 2647 2090 2659 2141
rect 2711 2091 2723 2142
rect 2775 2092 2787 2143
rect 2839 2093 2851 2144
rect 2903 2094 2915 2145
rect 2903 2093 2979 2094
rect 2839 2092 2979 2093
rect 2775 2091 2979 2092
rect 2711 2090 2979 2091
rect 2647 2089 2979 2090
rect 1933 2081 2979 2089
rect 1933 2080 2915 2081
rect 1933 2079 2851 2080
rect 1933 2027 2403 2079
rect 2455 2078 2787 2079
rect 2455 2027 2467 2078
rect 1933 2026 2467 2027
rect 2519 2077 2723 2078
rect 2519 2026 2531 2077
rect 1933 2025 2531 2026
rect 2583 2076 2659 2077
rect 2583 2025 2595 2076
rect 1933 2024 2595 2025
rect 2647 2025 2659 2076
rect 2711 2026 2723 2077
rect 2775 2027 2787 2078
rect 2839 2028 2851 2079
rect 2903 2029 2915 2080
rect 2967 2030 2979 2081
rect 2967 2029 3043 2030
rect 2903 2028 3043 2029
rect 2839 2027 3043 2028
rect 2775 2026 3043 2027
rect 2711 2025 3043 2026
rect 2647 2024 3043 2025
rect 1933 2017 3043 2024
rect 1933 2016 2979 2017
rect 1933 2015 2915 2016
rect 1933 2014 2851 2015
rect 1933 1962 2403 2014
rect 2455 2013 2787 2014
rect 2455 1962 2467 2013
rect 1933 1961 2467 1962
rect 2519 2012 2723 2013
rect 2519 1961 2531 2012
rect 1933 1960 2531 1961
rect 2583 2011 2659 2012
rect 2583 1960 2595 2011
rect 1933 1959 2595 1960
rect 2647 1960 2659 2011
rect 2711 1961 2723 2012
rect 2775 1962 2787 2013
rect 2839 1963 2851 2014
rect 2903 1964 2915 2015
rect 2967 1965 2979 2016
rect 3031 1966 3043 2017
rect 3937 3027 3938 3079
rect 3990 3027 4020 3079
rect 4072 3027 4102 3079
rect 4154 3027 4184 3079
rect 4236 3027 4237 3079
rect 3937 3012 4237 3027
rect 3937 2960 3938 3012
rect 3990 2960 4020 3012
rect 4072 2960 4102 3012
rect 4154 2960 4184 3012
rect 4236 2960 4237 3012
rect 3937 2945 4237 2960
rect 3937 2893 3938 2945
rect 3990 2893 4020 2945
rect 4072 2893 4102 2945
rect 4154 2893 4184 2945
rect 4236 2893 4237 2945
rect 3937 2878 4237 2893
rect 3937 2826 3938 2878
rect 3990 2826 4020 2878
rect 4072 2826 4102 2878
rect 4154 2826 4184 2878
rect 4236 2826 4237 2878
rect 3937 2811 4237 2826
rect 3937 2759 3938 2811
rect 3990 2759 4020 2811
rect 4072 2759 4102 2811
rect 4154 2759 4184 2811
rect 4236 2759 4237 2811
rect 3937 2744 4237 2759
rect 3937 2692 3938 2744
rect 3990 2692 4020 2744
rect 4072 2692 4102 2744
rect 4154 2692 4184 2744
rect 4236 2692 4237 2744
rect 3937 2677 4237 2692
rect 3937 2625 3938 2677
rect 3990 2625 4020 2677
rect 4072 2625 4102 2677
rect 4154 2625 4184 2677
rect 4236 2625 4237 2677
rect 3937 2610 4237 2625
rect 3937 2558 3938 2610
rect 3990 2558 4020 2610
rect 4072 2558 4102 2610
rect 4154 2558 4184 2610
rect 4236 2558 4237 2610
rect 3937 2543 4237 2558
rect 3937 2491 3938 2543
rect 3990 2491 4020 2543
rect 4072 2491 4102 2543
rect 4154 2491 4184 2543
rect 4236 2491 4237 2543
rect 3937 2476 4237 2491
rect 3937 2424 3938 2476
rect 3990 2424 4020 2476
rect 4072 2424 4102 2476
rect 4154 2424 4184 2476
rect 4236 2424 4237 2476
rect 3937 2409 4237 2424
rect 3937 2357 3938 2409
rect 3990 2357 4020 2409
rect 4072 2357 4102 2409
rect 4154 2357 4184 2409
rect 4236 2357 4237 2409
rect 3937 2342 4237 2357
rect 3937 2290 3938 2342
rect 3990 2290 4020 2342
rect 4072 2290 4102 2342
rect 4154 2290 4184 2342
rect 4236 2290 4237 2342
rect 3937 2275 4237 2290
rect 3937 2223 3938 2275
rect 3990 2223 4020 2275
rect 4072 2223 4102 2275
rect 4154 2223 4184 2275
rect 4236 2223 4237 2275
rect 3937 2208 4237 2223
rect 3937 2156 3938 2208
rect 3990 2156 4020 2208
rect 4072 2156 4102 2208
rect 4154 2156 4184 2208
rect 4236 2156 4237 2208
rect 3937 2141 4237 2156
rect 3937 2089 3938 2141
rect 3990 2089 4020 2141
rect 4072 2089 4102 2141
rect 4154 2089 4184 2141
rect 4236 2089 4237 2141
rect 3937 2074 4237 2089
rect 3937 2022 3938 2074
rect 3990 2022 4020 2074
rect 4072 2022 4102 2074
rect 4154 2022 4184 2074
rect 4236 2022 4237 2074
rect 3937 2016 4237 2022
rect 4761 3410 5061 3416
rect 4761 3358 4762 3410
rect 4814 3358 4844 3410
rect 4896 3358 4926 3410
rect 4978 3358 5008 3410
rect 5060 3358 5061 3410
rect 4761 3344 5061 3358
rect 4761 3292 4762 3344
rect 4814 3292 4844 3344
rect 4896 3292 4926 3344
rect 4978 3292 5008 3344
rect 5060 3292 5061 3344
rect 4761 3278 5061 3292
rect 4761 3226 4762 3278
rect 4814 3226 4844 3278
rect 4896 3226 4926 3278
rect 4978 3226 5008 3278
rect 5060 3226 5061 3278
rect 4761 3212 5061 3226
rect 4761 3160 4762 3212
rect 4814 3160 4844 3212
rect 4896 3160 4926 3212
rect 4978 3160 5008 3212
rect 5060 3160 5061 3212
rect 4761 3146 5061 3160
rect 4761 3094 4762 3146
rect 4814 3094 4844 3146
rect 4896 3094 4926 3146
rect 4978 3094 5008 3146
rect 5060 3094 5061 3146
rect 4761 3079 5061 3094
rect 4761 3027 4762 3079
rect 4814 3027 4844 3079
rect 4896 3027 4926 3079
rect 4978 3027 5008 3079
rect 5060 3027 5061 3079
rect 4761 3012 5061 3027
rect 4761 2960 4762 3012
rect 4814 2960 4844 3012
rect 4896 2960 4926 3012
rect 4978 2960 5008 3012
rect 5060 2960 5061 3012
rect 4761 2945 5061 2960
rect 4761 2893 4762 2945
rect 4814 2893 4844 2945
rect 4896 2893 4926 2945
rect 4978 2893 5008 2945
rect 5060 2893 5061 2945
rect 4761 2878 5061 2893
rect 4761 2826 4762 2878
rect 4814 2826 4844 2878
rect 4896 2826 4926 2878
rect 4978 2826 5008 2878
rect 5060 2826 5061 2878
rect 4761 2811 5061 2826
rect 4761 2759 4762 2811
rect 4814 2759 4844 2811
rect 4896 2759 4926 2811
rect 4978 2759 5008 2811
rect 5060 2759 5061 2811
rect 4761 2744 5061 2759
rect 4761 2692 4762 2744
rect 4814 2692 4844 2744
rect 4896 2692 4926 2744
rect 4978 2692 5008 2744
rect 5060 2692 5061 2744
rect 4761 2677 5061 2692
rect 4761 2625 4762 2677
rect 4814 2625 4844 2677
rect 4896 2625 4926 2677
rect 4978 2625 5008 2677
rect 5060 2625 5061 2677
rect 4761 2610 5061 2625
rect 4761 2558 4762 2610
rect 4814 2558 4844 2610
rect 4896 2558 4926 2610
rect 4978 2558 5008 2610
rect 5060 2558 5061 2610
rect 4761 2543 5061 2558
rect 4761 2491 4762 2543
rect 4814 2491 4844 2543
rect 4896 2491 4926 2543
rect 4978 2491 5008 2543
rect 5060 2491 5061 2543
rect 4761 2476 5061 2491
rect 4761 2424 4762 2476
rect 4814 2424 4844 2476
rect 4896 2424 4926 2476
rect 4978 2424 5008 2476
rect 5060 2424 5061 2476
rect 4761 2409 5061 2424
rect 4761 2357 4762 2409
rect 4814 2357 4844 2409
rect 4896 2357 4926 2409
rect 4978 2357 5008 2409
rect 5060 2357 5061 2409
rect 4761 2342 5061 2357
rect 4761 2290 4762 2342
rect 4814 2290 4844 2342
rect 4896 2290 4926 2342
rect 4978 2290 5008 2342
rect 5060 2290 5061 2342
rect 4761 2275 5061 2290
rect 4761 2223 4762 2275
rect 4814 2223 4844 2275
rect 4896 2223 4926 2275
rect 4978 2223 5008 2275
rect 5060 2223 5061 2275
rect 4761 2208 5061 2223
rect 4761 2156 4762 2208
rect 4814 2156 4844 2208
rect 4896 2156 4926 2208
rect 4978 2156 5008 2208
rect 5060 2156 5061 2208
rect 4761 2141 5061 2156
rect 4761 2089 4762 2141
rect 4814 2089 4844 2141
rect 4896 2089 4926 2141
rect 4978 2089 5008 2141
rect 5060 2089 5061 2141
rect 4761 2074 5061 2089
rect 4761 2022 4762 2074
rect 4814 2022 4844 2074
rect 4896 2022 4926 2074
rect 4978 2022 5008 2074
rect 5060 2022 5061 2074
rect 4761 2016 5061 2022
rect 5585 3410 5885 3416
rect 5585 3358 5586 3410
rect 5638 3358 5668 3410
rect 5720 3358 5750 3410
rect 5802 3358 5832 3410
rect 5884 3358 5885 3410
rect 5585 3344 5885 3358
rect 5585 3292 5586 3344
rect 5638 3292 5668 3344
rect 5720 3292 5750 3344
rect 5802 3292 5832 3344
rect 5884 3292 5885 3344
rect 5585 3278 5885 3292
rect 5585 3226 5586 3278
rect 5638 3226 5668 3278
rect 5720 3226 5750 3278
rect 5802 3226 5832 3278
rect 5884 3226 5885 3278
rect 5585 3212 5885 3226
rect 5585 3160 5586 3212
rect 5638 3160 5668 3212
rect 5720 3160 5750 3212
rect 5802 3160 5832 3212
rect 5884 3160 5885 3212
rect 5585 3146 5885 3160
rect 5585 3094 5586 3146
rect 5638 3094 5668 3146
rect 5720 3094 5750 3146
rect 5802 3094 5832 3146
rect 5884 3094 5885 3146
rect 5585 3079 5885 3094
rect 5585 3027 5586 3079
rect 5638 3027 5668 3079
rect 5720 3027 5750 3079
rect 5802 3027 5832 3079
rect 5884 3027 5885 3079
rect 5585 3012 5885 3027
rect 5585 2960 5586 3012
rect 5638 2960 5668 3012
rect 5720 2960 5750 3012
rect 5802 2960 5832 3012
rect 5884 2960 5885 3012
rect 5585 2945 5885 2960
rect 5585 2893 5586 2945
rect 5638 2893 5668 2945
rect 5720 2893 5750 2945
rect 5802 2893 5832 2945
rect 5884 2893 5885 2945
rect 5585 2878 5885 2893
rect 5585 2826 5586 2878
rect 5638 2826 5668 2878
rect 5720 2826 5750 2878
rect 5802 2826 5832 2878
rect 5884 2826 5885 2878
rect 5585 2811 5885 2826
rect 5585 2759 5586 2811
rect 5638 2759 5668 2811
rect 5720 2759 5750 2811
rect 5802 2759 5832 2811
rect 5884 2759 5885 2811
rect 5585 2744 5885 2759
rect 5585 2692 5586 2744
rect 5638 2692 5668 2744
rect 5720 2692 5750 2744
rect 5802 2692 5832 2744
rect 5884 2692 5885 2744
rect 5585 2677 5885 2692
rect 5585 2625 5586 2677
rect 5638 2625 5668 2677
rect 5720 2625 5750 2677
rect 5802 2625 5832 2677
rect 5884 2625 5885 2677
rect 5585 2610 5885 2625
rect 5585 2558 5586 2610
rect 5638 2558 5668 2610
rect 5720 2558 5750 2610
rect 5802 2558 5832 2610
rect 5884 2558 5885 2610
rect 5585 2543 5885 2558
rect 5585 2491 5586 2543
rect 5638 2491 5668 2543
rect 5720 2491 5750 2543
rect 5802 2491 5832 2543
rect 5884 2491 5885 2543
rect 5585 2476 5885 2491
rect 5585 2424 5586 2476
rect 5638 2424 5668 2476
rect 5720 2424 5750 2476
rect 5802 2424 5832 2476
rect 5884 2424 5885 2476
rect 5585 2409 5885 2424
rect 5585 2357 5586 2409
rect 5638 2357 5668 2409
rect 5720 2357 5750 2409
rect 5802 2357 5832 2409
rect 5884 2357 5885 2409
rect 5585 2342 5885 2357
rect 5585 2290 5586 2342
rect 5638 2290 5668 2342
rect 5720 2290 5750 2342
rect 5802 2290 5832 2342
rect 5884 2290 5885 2342
rect 5585 2275 5885 2290
rect 5585 2223 5586 2275
rect 5638 2223 5668 2275
rect 5720 2223 5750 2275
rect 5802 2223 5832 2275
rect 5884 2223 5885 2275
rect 5585 2208 5885 2223
rect 5585 2156 5586 2208
rect 5638 2156 5668 2208
rect 5720 2156 5750 2208
rect 5802 2156 5832 2208
rect 5884 2156 5885 2208
rect 5585 2141 5885 2156
rect 5585 2089 5586 2141
rect 5638 2089 5668 2141
rect 5720 2089 5750 2141
rect 5802 2089 5832 2141
rect 5884 2089 5885 2141
rect 5585 2074 5885 2089
rect 5585 2022 5586 2074
rect 5638 2022 5668 2074
rect 5720 2022 5750 2074
rect 5802 2022 5832 2074
rect 5884 2022 5885 2074
rect 5585 2016 5885 2022
rect 6409 3410 6709 3416
rect 6409 3358 6410 3410
rect 6462 3358 6492 3410
rect 6544 3358 6574 3410
rect 6626 3358 6656 3410
rect 6708 3358 6709 3410
rect 6409 3344 6709 3358
rect 6409 3292 6410 3344
rect 6462 3292 6492 3344
rect 6544 3292 6574 3344
rect 6626 3292 6656 3344
rect 6708 3292 6709 3344
rect 6409 3278 6709 3292
rect 6409 3226 6410 3278
rect 6462 3226 6492 3278
rect 6544 3226 6574 3278
rect 6626 3226 6656 3278
rect 6708 3226 6709 3278
rect 6409 3212 6709 3226
rect 6409 3160 6410 3212
rect 6462 3160 6492 3212
rect 6544 3160 6574 3212
rect 6626 3160 6656 3212
rect 6708 3160 6709 3212
rect 6409 3146 6709 3160
rect 6409 3094 6410 3146
rect 6462 3094 6492 3146
rect 6544 3094 6574 3146
rect 6626 3094 6656 3146
rect 6708 3094 6709 3146
rect 6409 3079 6709 3094
rect 6409 3027 6410 3079
rect 6462 3027 6492 3079
rect 6544 3027 6574 3079
rect 6626 3027 6656 3079
rect 6708 3027 6709 3079
rect 6409 3012 6709 3027
rect 6409 2960 6410 3012
rect 6462 2960 6492 3012
rect 6544 2960 6574 3012
rect 6626 2960 6656 3012
rect 6708 2960 6709 3012
rect 6409 2945 6709 2960
rect 6409 2893 6410 2945
rect 6462 2893 6492 2945
rect 6544 2893 6574 2945
rect 6626 2893 6656 2945
rect 6708 2893 6709 2945
rect 6409 2878 6709 2893
rect 6409 2826 6410 2878
rect 6462 2826 6492 2878
rect 6544 2826 6574 2878
rect 6626 2826 6656 2878
rect 6708 2826 6709 2878
rect 6409 2811 6709 2826
rect 6409 2759 6410 2811
rect 6462 2759 6492 2811
rect 6544 2759 6574 2811
rect 6626 2759 6656 2811
rect 6708 2759 6709 2811
rect 6409 2744 6709 2759
rect 6409 2692 6410 2744
rect 6462 2692 6492 2744
rect 6544 2692 6574 2744
rect 6626 2692 6656 2744
rect 6708 2692 6709 2744
rect 6409 2677 6709 2692
rect 6409 2625 6410 2677
rect 6462 2625 6492 2677
rect 6544 2625 6574 2677
rect 6626 2625 6656 2677
rect 6708 2625 6709 2677
rect 6409 2610 6709 2625
rect 6409 2558 6410 2610
rect 6462 2558 6492 2610
rect 6544 2558 6574 2610
rect 6626 2558 6656 2610
rect 6708 2558 6709 2610
rect 6409 2543 6709 2558
rect 6409 2491 6410 2543
rect 6462 2491 6492 2543
rect 6544 2491 6574 2543
rect 6626 2491 6656 2543
rect 6708 2491 6709 2543
rect 6409 2476 6709 2491
rect 6409 2424 6410 2476
rect 6462 2424 6492 2476
rect 6544 2424 6574 2476
rect 6626 2424 6656 2476
rect 6708 2424 6709 2476
rect 6409 2409 6709 2424
rect 6409 2357 6410 2409
rect 6462 2357 6492 2409
rect 6544 2357 6574 2409
rect 6626 2357 6656 2409
rect 6708 2357 6709 2409
rect 6409 2342 6709 2357
rect 6409 2290 6410 2342
rect 6462 2290 6492 2342
rect 6544 2290 6574 2342
rect 6626 2290 6656 2342
rect 6708 2290 6709 2342
rect 6409 2275 6709 2290
rect 6409 2223 6410 2275
rect 6462 2223 6492 2275
rect 6544 2223 6574 2275
rect 6626 2223 6656 2275
rect 6708 2223 6709 2275
rect 6409 2208 6709 2223
rect 6409 2156 6410 2208
rect 6462 2156 6492 2208
rect 6544 2156 6574 2208
rect 6626 2156 6656 2208
rect 6708 2156 6709 2208
rect 6409 2141 6709 2156
rect 6409 2089 6410 2141
rect 6462 2089 6492 2141
rect 6544 2089 6574 2141
rect 6626 2089 6656 2141
rect 6708 2089 6709 2141
rect 6409 2074 6709 2089
rect 6409 2022 6410 2074
rect 6462 2022 6492 2074
rect 6544 2022 6574 2074
rect 6626 2022 6656 2074
rect 6708 2022 6709 2074
rect 6409 2016 6709 2022
rect 7523 3410 7823 3416
rect 7523 3358 7524 3410
rect 7576 3358 7606 3410
rect 7658 3358 7688 3410
rect 7740 3358 7770 3410
rect 7822 3358 7823 3410
rect 7523 3344 7823 3358
rect 7523 3292 7524 3344
rect 7576 3292 7606 3344
rect 7658 3292 7688 3344
rect 7740 3292 7770 3344
rect 7822 3292 7823 3344
rect 7523 3278 7823 3292
rect 7523 3226 7524 3278
rect 7576 3226 7606 3278
rect 7658 3226 7688 3278
rect 7740 3226 7770 3278
rect 7822 3226 7823 3278
rect 7523 3212 7823 3226
rect 7523 3160 7524 3212
rect 7576 3160 7606 3212
rect 7658 3160 7688 3212
rect 7740 3160 7770 3212
rect 7822 3160 7823 3212
rect 7523 3146 7823 3160
rect 7523 3094 7524 3146
rect 7576 3094 7606 3146
rect 7658 3094 7688 3146
rect 7740 3094 7770 3146
rect 7822 3094 7823 3146
rect 7523 3079 7823 3094
rect 7523 3027 7524 3079
rect 7576 3027 7606 3079
rect 7658 3027 7688 3079
rect 7740 3027 7770 3079
rect 7822 3027 7823 3079
rect 7523 3012 7823 3027
rect 7523 2960 7524 3012
rect 7576 2960 7606 3012
rect 7658 2960 7688 3012
rect 7740 2960 7770 3012
rect 7822 2960 7823 3012
rect 7523 2945 7823 2960
rect 7523 2893 7524 2945
rect 7576 2893 7606 2945
rect 7658 2893 7688 2945
rect 7740 2893 7770 2945
rect 7822 2893 7823 2945
rect 7523 2878 7823 2893
rect 7523 2826 7524 2878
rect 7576 2826 7606 2878
rect 7658 2826 7688 2878
rect 7740 2826 7770 2878
rect 7822 2826 7823 2878
rect 7523 2811 7823 2826
rect 7523 2759 7524 2811
rect 7576 2759 7606 2811
rect 7658 2759 7688 2811
rect 7740 2759 7770 2811
rect 7822 2759 7823 2811
rect 7523 2744 7823 2759
rect 7523 2692 7524 2744
rect 7576 2692 7606 2744
rect 7658 2692 7688 2744
rect 7740 2692 7770 2744
rect 7822 2692 7823 2744
rect 7523 2677 7823 2692
rect 7523 2625 7524 2677
rect 7576 2625 7606 2677
rect 7658 2625 7688 2677
rect 7740 2625 7770 2677
rect 7822 2625 7823 2677
rect 7523 2610 7823 2625
rect 7523 2558 7524 2610
rect 7576 2558 7606 2610
rect 7658 2558 7688 2610
rect 7740 2558 7770 2610
rect 7822 2558 7823 2610
rect 7523 2543 7823 2558
rect 7523 2491 7524 2543
rect 7576 2491 7606 2543
rect 7658 2491 7688 2543
rect 7740 2491 7770 2543
rect 7822 2491 7823 2543
rect 7523 2476 7823 2491
rect 7523 2424 7524 2476
rect 7576 2424 7606 2476
rect 7658 2424 7688 2476
rect 7740 2424 7770 2476
rect 7822 2424 7823 2476
rect 7523 2409 7823 2424
rect 7523 2357 7524 2409
rect 7576 2357 7606 2409
rect 7658 2357 7688 2409
rect 7740 2357 7770 2409
rect 7822 2357 7823 2409
rect 7523 2342 7823 2357
rect 7523 2290 7524 2342
rect 7576 2290 7606 2342
rect 7658 2290 7688 2342
rect 7740 2290 7770 2342
rect 7822 2290 7823 2342
rect 7523 2275 7823 2290
rect 7523 2223 7524 2275
rect 7576 2223 7606 2275
rect 7658 2223 7688 2275
rect 7740 2223 7770 2275
rect 7822 2223 7823 2275
rect 7523 2208 7823 2223
rect 7523 2156 7524 2208
rect 7576 2156 7606 2208
rect 7658 2156 7688 2208
rect 7740 2156 7770 2208
rect 7822 2156 7823 2208
rect 7523 2141 7823 2156
rect 7523 2089 7524 2141
rect 7576 2089 7606 2141
rect 7658 2089 7688 2141
rect 7740 2089 7770 2141
rect 7822 2089 7823 2141
rect 7523 2074 7823 2089
rect 7523 2022 7524 2074
rect 7576 2022 7606 2074
rect 7658 2022 7688 2074
rect 7740 2022 7770 2074
rect 7822 2022 7823 2074
rect 7523 2016 7823 2022
rect 8347 3410 8647 3416
rect 8347 3358 8348 3410
rect 8400 3358 8430 3410
rect 8482 3358 8512 3410
rect 8564 3358 8594 3410
rect 8646 3358 8647 3410
rect 8347 3344 8647 3358
rect 8347 3292 8348 3344
rect 8400 3292 8430 3344
rect 8482 3292 8512 3344
rect 8564 3292 8594 3344
rect 8646 3292 8647 3344
rect 8347 3278 8647 3292
rect 8347 3226 8348 3278
rect 8400 3226 8430 3278
rect 8482 3226 8512 3278
rect 8564 3226 8594 3278
rect 8646 3226 8647 3278
rect 8347 3212 8647 3226
rect 8347 3160 8348 3212
rect 8400 3160 8430 3212
rect 8482 3160 8512 3212
rect 8564 3160 8594 3212
rect 8646 3160 8647 3212
rect 8347 3146 8647 3160
rect 8347 3094 8348 3146
rect 8400 3094 8430 3146
rect 8482 3094 8512 3146
rect 8564 3094 8594 3146
rect 8646 3094 8647 3146
rect 8347 3079 8647 3094
rect 8347 3027 8348 3079
rect 8400 3027 8430 3079
rect 8482 3027 8512 3079
rect 8564 3027 8594 3079
rect 8646 3027 8647 3079
rect 8347 3012 8647 3027
rect 8347 2960 8348 3012
rect 8400 2960 8430 3012
rect 8482 2960 8512 3012
rect 8564 2960 8594 3012
rect 8646 2960 8647 3012
rect 8347 2945 8647 2960
rect 8347 2893 8348 2945
rect 8400 2893 8430 2945
rect 8482 2893 8512 2945
rect 8564 2893 8594 2945
rect 8646 2893 8647 2945
rect 8347 2878 8647 2893
rect 8347 2826 8348 2878
rect 8400 2826 8430 2878
rect 8482 2826 8512 2878
rect 8564 2826 8594 2878
rect 8646 2826 8647 2878
rect 8347 2811 8647 2826
rect 8347 2759 8348 2811
rect 8400 2759 8430 2811
rect 8482 2759 8512 2811
rect 8564 2759 8594 2811
rect 8646 2759 8647 2811
rect 8347 2744 8647 2759
rect 8347 2692 8348 2744
rect 8400 2692 8430 2744
rect 8482 2692 8512 2744
rect 8564 2692 8594 2744
rect 8646 2692 8647 2744
rect 8347 2677 8647 2692
rect 8347 2625 8348 2677
rect 8400 2625 8430 2677
rect 8482 2625 8512 2677
rect 8564 2625 8594 2677
rect 8646 2625 8647 2677
rect 8347 2610 8647 2625
rect 8347 2558 8348 2610
rect 8400 2558 8430 2610
rect 8482 2558 8512 2610
rect 8564 2558 8594 2610
rect 8646 2558 8647 2610
rect 8347 2543 8647 2558
rect 8347 2491 8348 2543
rect 8400 2491 8430 2543
rect 8482 2491 8512 2543
rect 8564 2491 8594 2543
rect 8646 2491 8647 2543
rect 8347 2476 8647 2491
rect 8347 2424 8348 2476
rect 8400 2424 8430 2476
rect 8482 2424 8512 2476
rect 8564 2424 8594 2476
rect 8646 2424 8647 2476
rect 8347 2409 8647 2424
rect 8347 2357 8348 2409
rect 8400 2357 8430 2409
rect 8482 2357 8512 2409
rect 8564 2357 8594 2409
rect 8646 2357 8647 2409
rect 8347 2342 8647 2357
rect 8347 2290 8348 2342
rect 8400 2290 8430 2342
rect 8482 2290 8512 2342
rect 8564 2290 8594 2342
rect 8646 2290 8647 2342
rect 8347 2275 8647 2290
rect 8347 2223 8348 2275
rect 8400 2223 8430 2275
rect 8482 2223 8512 2275
rect 8564 2223 8594 2275
rect 8646 2223 8647 2275
rect 8347 2208 8647 2223
rect 8347 2156 8348 2208
rect 8400 2156 8430 2208
rect 8482 2156 8512 2208
rect 8564 2156 8594 2208
rect 8646 2156 8647 2208
rect 8347 2141 8647 2156
rect 8347 2089 8348 2141
rect 8400 2089 8430 2141
rect 8482 2089 8512 2141
rect 8564 2089 8594 2141
rect 8646 2089 8647 2141
rect 8347 2074 8647 2089
rect 8347 2022 8348 2074
rect 8400 2022 8430 2074
rect 8482 2022 8512 2074
rect 8564 2022 8594 2074
rect 8646 2022 8647 2074
rect 8347 2016 8647 2022
rect 9171 3410 9471 3416
rect 9171 3358 9172 3410
rect 9224 3358 9254 3410
rect 9306 3358 9336 3410
rect 9388 3358 9418 3410
rect 9470 3358 9471 3410
rect 9171 3344 9471 3358
rect 9171 3292 9172 3344
rect 9224 3292 9254 3344
rect 9306 3292 9336 3344
rect 9388 3292 9418 3344
rect 9470 3292 9471 3344
rect 9171 3278 9471 3292
rect 9171 3226 9172 3278
rect 9224 3226 9254 3278
rect 9306 3226 9336 3278
rect 9388 3226 9418 3278
rect 9470 3226 9471 3278
rect 9171 3212 9471 3226
rect 9171 3160 9172 3212
rect 9224 3160 9254 3212
rect 9306 3160 9336 3212
rect 9388 3160 9418 3212
rect 9470 3160 9471 3212
rect 9171 3146 9471 3160
rect 9171 3094 9172 3146
rect 9224 3094 9254 3146
rect 9306 3094 9336 3146
rect 9388 3094 9418 3146
rect 9470 3094 9471 3146
rect 9171 3079 9471 3094
rect 9171 3027 9172 3079
rect 9224 3027 9254 3079
rect 9306 3027 9336 3079
rect 9388 3027 9418 3079
rect 9470 3027 9471 3079
rect 9171 3012 9471 3027
rect 9171 2960 9172 3012
rect 9224 2960 9254 3012
rect 9306 2960 9336 3012
rect 9388 2960 9418 3012
rect 9470 2960 9471 3012
rect 9171 2945 9471 2960
rect 9171 2893 9172 2945
rect 9224 2893 9254 2945
rect 9306 2893 9336 2945
rect 9388 2893 9418 2945
rect 9470 2893 9471 2945
rect 9171 2878 9471 2893
rect 9171 2826 9172 2878
rect 9224 2826 9254 2878
rect 9306 2826 9336 2878
rect 9388 2826 9418 2878
rect 9470 2826 9471 2878
rect 9171 2811 9471 2826
rect 9171 2759 9172 2811
rect 9224 2759 9254 2811
rect 9306 2759 9336 2811
rect 9388 2759 9418 2811
rect 9470 2759 9471 2811
rect 9171 2744 9471 2759
rect 9171 2692 9172 2744
rect 9224 2692 9254 2744
rect 9306 2692 9336 2744
rect 9388 2692 9418 2744
rect 9470 2692 9471 2744
rect 9171 2677 9471 2692
rect 9171 2625 9172 2677
rect 9224 2625 9254 2677
rect 9306 2625 9336 2677
rect 9388 2625 9418 2677
rect 9470 2625 9471 2677
rect 9171 2610 9471 2625
rect 9171 2558 9172 2610
rect 9224 2558 9254 2610
rect 9306 2558 9336 2610
rect 9388 2558 9418 2610
rect 9470 2558 9471 2610
rect 9171 2543 9471 2558
rect 9171 2491 9172 2543
rect 9224 2491 9254 2543
rect 9306 2491 9336 2543
rect 9388 2491 9418 2543
rect 9470 2491 9471 2543
rect 9171 2476 9471 2491
rect 9171 2424 9172 2476
rect 9224 2424 9254 2476
rect 9306 2424 9336 2476
rect 9388 2424 9418 2476
rect 9470 2424 9471 2476
rect 9171 2409 9471 2424
rect 9171 2357 9172 2409
rect 9224 2357 9254 2409
rect 9306 2357 9336 2409
rect 9388 2357 9418 2409
rect 9470 2357 9471 2409
rect 9171 2342 9471 2357
rect 9171 2290 9172 2342
rect 9224 2290 9254 2342
rect 9306 2290 9336 2342
rect 9388 2290 9418 2342
rect 9470 2290 9471 2342
rect 9171 2275 9471 2290
rect 9171 2223 9172 2275
rect 9224 2223 9254 2275
rect 9306 2223 9336 2275
rect 9388 2223 9418 2275
rect 9470 2223 9471 2275
rect 9171 2208 9471 2223
rect 9171 2156 9172 2208
rect 9224 2156 9254 2208
rect 9306 2156 9336 2208
rect 9388 2156 9418 2208
rect 9470 2156 9471 2208
rect 9171 2141 9471 2156
rect 9171 2089 9172 2141
rect 9224 2089 9254 2141
rect 9306 2089 9336 2141
rect 9388 2089 9418 2141
rect 9470 2089 9471 2141
rect 9171 2074 9471 2089
rect 9171 2022 9172 2074
rect 9224 2022 9254 2074
rect 9306 2022 9336 2074
rect 9388 2022 9418 2074
rect 9470 2022 9471 2074
rect 9171 2016 9471 2022
rect 9995 3410 10295 3416
rect 9995 3358 9996 3410
rect 10048 3358 10078 3410
rect 10130 3358 10160 3410
rect 10212 3358 10242 3410
rect 10294 3358 10295 3410
rect 9995 3344 10295 3358
rect 9995 3292 9996 3344
rect 10048 3292 10078 3344
rect 10130 3292 10160 3344
rect 10212 3292 10242 3344
rect 10294 3292 10295 3344
rect 9995 3278 10295 3292
rect 9995 3226 9996 3278
rect 10048 3226 10078 3278
rect 10130 3226 10160 3278
rect 10212 3226 10242 3278
rect 10294 3226 10295 3278
rect 9995 3212 10295 3226
rect 9995 3160 9996 3212
rect 10048 3160 10078 3212
rect 10130 3160 10160 3212
rect 10212 3160 10242 3212
rect 10294 3160 10295 3212
rect 9995 3146 10295 3160
rect 9995 3094 9996 3146
rect 10048 3094 10078 3146
rect 10130 3094 10160 3146
rect 10212 3094 10242 3146
rect 10294 3094 10295 3146
rect 9995 3079 10295 3094
rect 9995 3027 9996 3079
rect 10048 3027 10078 3079
rect 10130 3027 10160 3079
rect 10212 3027 10242 3079
rect 10294 3027 10295 3079
rect 9995 3012 10295 3027
rect 9995 2960 9996 3012
rect 10048 2960 10078 3012
rect 10130 2960 10160 3012
rect 10212 2960 10242 3012
rect 10294 2960 10295 3012
rect 9995 2945 10295 2960
rect 9995 2893 9996 2945
rect 10048 2893 10078 2945
rect 10130 2893 10160 2945
rect 10212 2893 10242 2945
rect 10294 2893 10295 2945
rect 9995 2878 10295 2893
rect 9995 2826 9996 2878
rect 10048 2826 10078 2878
rect 10130 2826 10160 2878
rect 10212 2826 10242 2878
rect 10294 2826 10295 2878
rect 9995 2811 10295 2826
rect 9995 2759 9996 2811
rect 10048 2759 10078 2811
rect 10130 2759 10160 2811
rect 10212 2759 10242 2811
rect 10294 2759 10295 2811
rect 9995 2744 10295 2759
rect 9995 2692 9996 2744
rect 10048 2692 10078 2744
rect 10130 2692 10160 2744
rect 10212 2692 10242 2744
rect 10294 2692 10295 2744
rect 9995 2677 10295 2692
rect 9995 2625 9996 2677
rect 10048 2625 10078 2677
rect 10130 2625 10160 2677
rect 10212 2625 10242 2677
rect 10294 2625 10295 2677
rect 9995 2610 10295 2625
rect 9995 2558 9996 2610
rect 10048 2558 10078 2610
rect 10130 2558 10160 2610
rect 10212 2558 10242 2610
rect 10294 2558 10295 2610
rect 9995 2543 10295 2558
rect 9995 2491 9996 2543
rect 10048 2491 10078 2543
rect 10130 2491 10160 2543
rect 10212 2491 10242 2543
rect 10294 2491 10295 2543
rect 9995 2476 10295 2491
rect 9995 2424 9996 2476
rect 10048 2424 10078 2476
rect 10130 2424 10160 2476
rect 10212 2424 10242 2476
rect 10294 2424 10295 2476
rect 9995 2409 10295 2424
rect 9995 2357 9996 2409
rect 10048 2357 10078 2409
rect 10130 2357 10160 2409
rect 10212 2357 10242 2409
rect 10294 2357 10295 2409
rect 9995 2342 10295 2357
rect 9995 2290 9996 2342
rect 10048 2290 10078 2342
rect 10130 2290 10160 2342
rect 10212 2290 10242 2342
rect 10294 2290 10295 2342
rect 9995 2275 10295 2290
rect 9995 2223 9996 2275
rect 10048 2223 10078 2275
rect 10130 2223 10160 2275
rect 10212 2223 10242 2275
rect 10294 2223 10295 2275
rect 9995 2208 10295 2223
rect 9995 2156 9996 2208
rect 10048 2156 10078 2208
rect 10130 2156 10160 2208
rect 10212 2156 10242 2208
rect 10294 2156 10295 2208
rect 9995 2141 10295 2156
rect 9995 2089 9996 2141
rect 10048 2089 10078 2141
rect 10130 2089 10160 2141
rect 10212 2089 10242 2141
rect 10294 2089 10295 2141
rect 9995 2074 10295 2089
rect 9995 2022 9996 2074
rect 10048 2022 10078 2074
rect 10130 2022 10160 2074
rect 10212 2022 10242 2074
rect 10294 2022 10295 2074
rect 9995 2016 10295 2022
rect 10819 3410 11119 3416
rect 10819 3358 10820 3410
rect 10872 3358 10902 3410
rect 10954 3358 10984 3410
rect 11036 3358 11066 3410
rect 11118 3358 11119 3410
rect 10819 3344 11119 3358
rect 10819 3292 10820 3344
rect 10872 3292 10902 3344
rect 10954 3292 10984 3344
rect 11036 3292 11066 3344
rect 11118 3292 11119 3344
rect 10819 3278 11119 3292
rect 10819 3226 10820 3278
rect 10872 3226 10902 3278
rect 10954 3226 10984 3278
rect 11036 3226 11066 3278
rect 11118 3226 11119 3278
rect 11384 3379 11514 3739
rect 11384 3273 11396 3379
rect 11502 3273 11514 3379
rect 11384 3267 11514 3273
rect 10819 3212 11119 3226
rect 10819 3160 10820 3212
rect 10872 3160 10902 3212
rect 10954 3160 10984 3212
rect 11036 3160 11066 3212
rect 11118 3160 11119 3212
rect 10819 3146 11119 3160
rect 10819 3094 10820 3146
rect 10872 3094 10902 3146
rect 10954 3094 10984 3146
rect 11036 3094 11066 3146
rect 11118 3094 11119 3146
rect 10819 3079 11119 3094
rect 10819 3027 10820 3079
rect 10872 3027 10902 3079
rect 10954 3027 10984 3079
rect 11036 3027 11066 3079
rect 11118 3027 11119 3079
rect 10819 3012 11119 3027
rect 10819 2960 10820 3012
rect 10872 2960 10902 3012
rect 10954 2960 10984 3012
rect 11036 2960 11066 3012
rect 11118 2960 11119 3012
rect 10819 2945 11119 2960
rect 10819 2893 10820 2945
rect 10872 2893 10902 2945
rect 10954 2893 10984 2945
rect 11036 2893 11066 2945
rect 11118 2893 11119 2945
rect 10819 2878 11119 2893
rect 10819 2826 10820 2878
rect 10872 2826 10902 2878
rect 10954 2826 10984 2878
rect 11036 2826 11066 2878
rect 11118 2826 11119 2878
rect 10819 2811 11119 2826
rect 10819 2759 10820 2811
rect 10872 2759 10902 2811
rect 10954 2759 10984 2811
rect 11036 2759 11066 2811
rect 11118 2759 11119 2811
rect 10819 2744 11119 2759
rect 10819 2692 10820 2744
rect 10872 2692 10902 2744
rect 10954 2692 10984 2744
rect 11036 2692 11066 2744
rect 11118 2692 11119 2744
rect 10819 2677 11119 2692
rect 10819 2625 10820 2677
rect 10872 2625 10902 2677
rect 10954 2625 10984 2677
rect 11036 2625 11066 2677
rect 11118 2625 11119 2677
rect 10819 2610 11119 2625
rect 10819 2558 10820 2610
rect 10872 2558 10902 2610
rect 10954 2558 10984 2610
rect 11036 2558 11066 2610
rect 11118 2558 11119 2610
rect 10819 2543 11119 2558
rect 10819 2491 10820 2543
rect 10872 2491 10902 2543
rect 10954 2491 10984 2543
rect 11036 2491 11066 2543
rect 11118 2491 11119 2543
rect 10819 2476 11119 2491
rect 10819 2424 10820 2476
rect 10872 2424 10902 2476
rect 10954 2424 10984 2476
rect 11036 2424 11066 2476
rect 11118 2424 11119 2476
rect 10819 2409 11119 2424
rect 10819 2357 10820 2409
rect 10872 2357 10902 2409
rect 10954 2357 10984 2409
rect 11036 2357 11066 2409
rect 11118 2357 11119 2409
rect 10819 2342 11119 2357
rect 10819 2290 10820 2342
rect 10872 2290 10902 2342
rect 10954 2290 10984 2342
rect 11036 2290 11066 2342
rect 11118 2290 11119 2342
rect 10819 2275 11119 2290
rect 10819 2223 10820 2275
rect 10872 2223 10902 2275
rect 10954 2223 10984 2275
rect 11036 2223 11066 2275
rect 11118 2223 11119 2275
rect 10819 2208 11119 2223
rect 10819 2156 10820 2208
rect 10872 2156 10902 2208
rect 10954 2156 10984 2208
rect 11036 2156 11066 2208
rect 11118 2156 11119 2208
rect 10819 2141 11119 2156
rect 10819 2089 10820 2141
rect 10872 2089 10902 2141
rect 10954 2089 10984 2141
rect 11036 2089 11066 2141
rect 11118 2089 11119 2141
rect 10819 2074 11119 2089
rect 10819 2022 10820 2074
rect 10872 2022 10902 2074
rect 10954 2022 10984 2074
rect 11036 2022 11066 2074
rect 11118 2022 11119 2074
rect 10819 2016 11119 2022
rect 3031 1965 3107 1966
rect 2967 1964 3107 1965
rect 2903 1963 3107 1964
rect 2839 1962 3107 1963
rect 2775 1961 3107 1962
rect 2711 1960 3107 1961
rect 2647 1959 3107 1960
rect 1933 1953 3107 1959
rect 1933 1952 3043 1953
rect 1933 1951 2979 1952
rect 1933 1950 2915 1951
rect 1933 1949 2851 1950
rect 1933 1897 2403 1949
rect 2455 1948 2787 1949
rect 2455 1897 2467 1948
rect 1933 1896 2467 1897
rect 2519 1947 2723 1948
rect 2519 1896 2531 1947
rect 1933 1895 2531 1896
rect 2583 1946 2659 1947
rect 2583 1895 2595 1946
rect 1933 1894 2595 1895
rect 2647 1895 2659 1946
rect 2711 1896 2723 1947
rect 2775 1897 2787 1948
rect 2839 1898 2851 1949
rect 2903 1899 2915 1950
rect 2967 1900 2979 1951
rect 3031 1901 3043 1952
rect 3095 1902 3107 1953
rect 3095 1901 3223 1902
rect 3031 1900 3223 1901
rect 2967 1899 3223 1900
rect 2903 1898 3223 1899
rect 2839 1897 3223 1898
rect 2775 1896 3223 1897
rect 2711 1895 3223 1896
rect 2647 1894 3223 1895
rect 1933 1889 3223 1894
rect 1933 1888 3107 1889
rect 1933 1887 3043 1888
rect 1933 1886 2979 1887
rect 1933 1885 2915 1886
rect 1933 1884 2851 1885
rect 1933 1832 2403 1884
rect 2455 1883 2787 1884
rect 2455 1832 2467 1883
rect 1933 1831 2467 1832
rect 2519 1882 2723 1883
rect 2519 1831 2531 1882
rect 1933 1830 2531 1831
rect 2583 1881 2659 1882
rect 2583 1830 2595 1881
rect 1933 1829 2595 1830
rect 2647 1830 2659 1881
rect 2711 1831 2723 1882
rect 2775 1832 2787 1883
rect 2839 1833 2851 1884
rect 2903 1834 2915 1885
rect 2967 1835 2979 1886
rect 3031 1836 3043 1887
rect 3095 1837 3107 1888
rect 3159 1837 3171 1889
rect 3095 1836 3223 1837
rect 3031 1835 3223 1836
rect 2967 1834 3223 1835
rect 2903 1833 3223 1834
rect 2839 1832 3223 1833
rect 2775 1831 3223 1832
rect 2711 1830 3223 1831
rect 2647 1829 3223 1830
rect 1933 1824 3223 1829
rect 1933 1823 3107 1824
rect 1933 1822 3043 1823
rect 1933 1821 2979 1822
rect 1933 1820 2915 1821
rect 1933 1819 2851 1820
rect 1933 1818 2787 1819
rect 1933 1766 2403 1818
rect 2455 1766 2467 1818
rect 2519 1817 2723 1818
rect 2519 1766 2531 1817
rect 1933 1765 2531 1766
rect 2583 1816 2659 1817
rect 2583 1765 2595 1816
rect 1933 1764 2595 1765
rect 2647 1765 2659 1816
rect 2711 1766 2723 1817
rect 2775 1767 2787 1818
rect 2839 1768 2851 1819
rect 2903 1769 2915 1820
rect 2967 1770 2979 1821
rect 3031 1771 3043 1822
rect 3095 1772 3107 1823
rect 3159 1772 3171 1824
rect 3095 1771 3223 1772
rect 3031 1770 3223 1771
rect 2967 1769 3223 1770
rect 2903 1768 3223 1769
rect 2839 1767 3223 1768
rect 2775 1766 3223 1767
rect 2711 1765 3223 1766
rect 2647 1764 3223 1765
rect 1933 1759 3223 1764
rect 1933 1758 3107 1759
rect 1933 1757 3043 1758
rect 1933 1756 2979 1757
rect 1933 1755 2915 1756
rect 1933 1754 2851 1755
rect 1933 1753 2787 1754
rect 1933 1752 2467 1753
rect 1933 1700 2403 1752
rect 2455 1701 2467 1752
rect 2519 1752 2723 1753
rect 2519 1701 2531 1752
rect 2455 1700 2531 1701
rect 2583 1751 2659 1752
rect 2583 1700 2595 1751
rect 1933 1699 2595 1700
rect 2647 1700 2659 1751
rect 2711 1701 2723 1752
rect 2775 1702 2787 1753
rect 2839 1703 2851 1754
rect 2903 1704 2915 1755
rect 2967 1705 2979 1756
rect 3031 1706 3043 1757
rect 3095 1707 3107 1758
rect 3159 1707 3171 1759
rect 3095 1706 3223 1707
rect 3031 1705 3223 1706
rect 2967 1704 3223 1705
rect 2903 1703 3223 1704
rect 2839 1702 3223 1703
rect 2775 1701 3223 1702
rect 2711 1700 3223 1701
rect 2647 1699 3223 1700
rect 1933 1694 3223 1699
rect 1933 1693 3107 1694
rect 1933 1692 3043 1693
rect 1933 1691 2979 1692
rect 1933 1690 2915 1691
rect 1933 1689 2851 1690
rect 1933 1688 2787 1689
rect 1933 1686 2467 1688
rect 1933 1634 2403 1686
rect 2455 1636 2467 1686
rect 2519 1687 2723 1688
rect 2519 1636 2531 1687
rect 2455 1635 2531 1636
rect 2583 1686 2659 1687
rect 2583 1635 2595 1686
rect 2455 1634 2595 1635
rect 2647 1635 2659 1686
rect 2711 1636 2723 1687
rect 2775 1637 2787 1688
rect 2839 1638 2851 1689
rect 2903 1639 2915 1690
rect 2967 1640 2979 1691
rect 3031 1641 3043 1692
rect 3095 1642 3107 1693
rect 3159 1642 3171 1694
rect 3095 1641 3223 1642
rect 3031 1640 3223 1641
rect 2967 1639 3223 1640
rect 2903 1638 3223 1639
rect 2839 1637 3223 1638
rect 2775 1636 3223 1637
rect 2711 1635 3223 1636
rect 2647 1634 3223 1635
rect 1933 1629 3223 1634
rect 1933 1628 3107 1629
rect 1933 1627 3043 1628
rect 1933 1626 2979 1627
rect 1933 1625 2915 1626
rect 1933 1624 2851 1625
rect 1933 1623 2787 1624
rect 1933 1622 2723 1623
rect 1933 1620 2467 1622
rect 1933 1568 2403 1620
rect 2455 1570 2467 1620
rect 2519 1570 2531 1622
rect 2583 1621 2659 1622
rect 2583 1570 2595 1621
rect 2455 1569 2595 1570
rect 2647 1570 2659 1621
rect 2711 1571 2723 1622
rect 2775 1572 2787 1623
rect 2839 1573 2851 1624
rect 2903 1574 2915 1625
rect 2967 1575 2979 1626
rect 3031 1576 3043 1627
rect 3095 1577 3107 1628
rect 3159 1577 3171 1629
rect 3095 1576 3223 1577
rect 3031 1575 3223 1576
rect 2967 1574 3223 1575
rect 2903 1573 3223 1574
rect 2839 1572 3223 1573
rect 2775 1571 3223 1572
rect 2711 1570 3223 1571
rect 2647 1569 3223 1570
rect 2455 1568 3223 1569
rect 1933 1564 3223 1568
rect 1933 1563 3107 1564
rect 1933 1562 3043 1563
rect 1933 1561 2979 1562
rect 1933 1560 2915 1561
rect 1933 1559 2851 1560
rect 1933 1558 2787 1559
rect 1933 1557 2723 1558
rect 1933 1556 2531 1557
rect 1933 1554 2467 1556
rect 1933 1502 2403 1554
rect 2455 1504 2467 1554
rect 2519 1505 2531 1556
rect 2583 1556 2659 1557
rect 2583 1505 2595 1556
rect 2519 1504 2595 1505
rect 2647 1505 2659 1556
rect 2711 1506 2723 1557
rect 2775 1507 2787 1558
rect 2839 1508 2851 1559
rect 2903 1509 2915 1560
rect 2967 1510 2979 1561
rect 3031 1511 3043 1562
rect 3095 1512 3107 1563
rect 3159 1512 3171 1564
rect 3095 1511 3223 1512
rect 3031 1510 3223 1511
rect 2967 1509 3223 1510
rect 2903 1508 3223 1509
rect 2839 1507 3223 1508
rect 2775 1506 3223 1507
rect 2711 1505 3223 1506
rect 2647 1504 3223 1505
rect 2455 1502 3223 1504
rect 1933 1499 3223 1502
rect 1933 1498 3107 1499
rect 1933 1497 3043 1498
rect 1933 1496 2979 1497
rect 1933 1495 2915 1496
rect 1933 1494 2851 1495
rect 1933 1493 2787 1494
rect 1933 1492 2723 1493
rect 1933 1490 2531 1492
rect 1933 1488 2467 1490
rect 1933 1436 1939 1488
rect 1991 1436 2006 1488
rect 2058 1436 2073 1488
rect 2125 1436 2139 1488
rect 2191 1436 2205 1488
rect 2257 1436 2271 1488
rect 2323 1436 2337 1488
rect 2389 1436 2403 1488
rect 2455 1438 2467 1488
rect 2519 1440 2531 1490
rect 2583 1491 2659 1492
rect 2583 1440 2595 1491
rect 2519 1439 2595 1440
rect 2647 1440 2659 1491
rect 2711 1441 2723 1492
rect 2775 1442 2787 1493
rect 2839 1443 2851 1494
rect 2903 1444 2915 1495
rect 2967 1445 2979 1496
rect 3031 1446 3043 1497
rect 3095 1447 3107 1498
rect 3159 1447 3171 1499
rect 3095 1446 3223 1447
rect 3031 1445 3223 1446
rect 2967 1444 3223 1445
rect 2903 1443 3223 1444
rect 2839 1442 3223 1443
rect 2775 1441 3223 1442
rect 2711 1440 3223 1441
rect 2647 1439 3223 1440
rect 2519 1438 3223 1439
rect 2455 1436 3223 1438
rect 1933 1434 3223 1436
rect 1933 1433 3107 1434
rect 1933 1432 3043 1433
rect 1933 1431 2979 1432
rect 1933 1430 2915 1431
rect 1933 1429 2851 1430
rect 1933 1428 2787 1429
rect 1933 1427 2723 1428
rect 1933 1426 2659 1427
rect 1933 1424 2531 1426
rect 1933 1372 1939 1424
rect 1991 1372 2005 1424
rect 2057 1372 2071 1424
rect 2123 1372 2137 1424
rect 2189 1372 2203 1424
rect 2255 1372 2269 1424
rect 2321 1372 2335 1424
rect 2387 1372 2401 1424
rect 2453 1372 2467 1424
rect 2519 1374 2531 1424
rect 2583 1374 2595 1426
rect 2647 1375 2659 1426
rect 2711 1376 2723 1427
rect 2775 1377 2787 1428
rect 2839 1378 2851 1429
rect 2903 1379 2915 1430
rect 2967 1380 2979 1431
rect 3031 1381 3043 1432
rect 3095 1382 3107 1433
rect 3159 1382 3171 1434
rect 3095 1381 3223 1382
rect 3031 1380 3223 1381
rect 2967 1379 3223 1380
rect 2903 1378 3223 1379
rect 2839 1377 3223 1378
rect 2775 1376 3223 1377
rect 2711 1375 3223 1376
rect 2647 1374 3223 1375
rect 2519 1372 3223 1374
rect 1933 1369 3223 1372
rect 1933 1368 3107 1369
rect 1933 1367 3043 1368
rect 1933 1366 2979 1367
rect 1933 1365 2915 1366
rect 1933 1364 2851 1365
rect 1933 1363 2787 1364
rect 1933 1362 2723 1363
rect 1933 1361 2659 1362
rect 1933 1360 2595 1361
rect 1933 1308 1939 1360
rect 1991 1308 2005 1360
rect 2057 1308 2071 1360
rect 2123 1308 2137 1360
rect 2189 1308 2203 1360
rect 2255 1308 2269 1360
rect 2321 1308 2335 1360
rect 2387 1308 2401 1360
rect 2453 1308 2466 1360
rect 2518 1308 2531 1360
rect 2583 1309 2595 1360
rect 2647 1310 2659 1361
rect 2711 1311 2723 1362
rect 2775 1312 2787 1363
rect 2839 1313 2851 1364
rect 2903 1314 2915 1365
rect 2967 1315 2979 1366
rect 3031 1316 3043 1367
rect 3095 1317 3107 1368
rect 3159 1317 3171 1369
rect 3095 1316 3223 1317
rect 3031 1315 3223 1316
rect 2967 1314 3223 1315
rect 2903 1313 3223 1314
rect 2839 1312 3223 1313
rect 2775 1311 3223 1312
rect 2711 1310 3223 1311
rect 2647 1309 3223 1310
rect 2583 1308 3223 1309
rect 1933 1304 3223 1308
rect 1933 1303 3107 1304
rect 1933 1302 3043 1303
rect 1933 1301 2979 1302
rect 1933 1300 2915 1301
rect 1933 1299 2851 1300
rect 1933 1298 2787 1299
rect 1933 1297 2723 1298
rect 1933 1296 2659 1297
rect 1933 1244 1939 1296
rect 1991 1244 2005 1296
rect 2057 1244 2071 1296
rect 2123 1244 2137 1296
rect 2189 1244 2203 1296
rect 2255 1244 2269 1296
rect 2321 1244 2335 1296
rect 2387 1244 2400 1296
rect 2452 1244 2465 1296
rect 2517 1244 2530 1296
rect 2582 1244 2595 1296
rect 2647 1245 2659 1296
rect 2711 1246 2723 1297
rect 2775 1247 2787 1298
rect 2839 1248 2851 1299
rect 2903 1249 2915 1300
rect 2967 1250 2979 1301
rect 3031 1251 3043 1302
rect 3095 1252 3107 1303
rect 3159 1252 3171 1304
rect 3095 1251 3223 1252
rect 3031 1250 3223 1251
rect 2967 1249 3223 1250
rect 2903 1248 3223 1249
rect 2839 1247 3223 1248
rect 2775 1246 3223 1247
rect 2711 1245 3223 1246
rect 2647 1244 3223 1245
rect 1933 1239 3223 1244
rect 1933 1238 3107 1239
rect 1933 1237 3043 1238
rect 1933 1236 2979 1237
rect 1933 1235 2915 1236
rect 1933 1234 2851 1235
rect 1933 1233 2787 1234
rect 1933 1232 2723 1233
rect 1933 1180 1939 1232
rect 1991 1180 2005 1232
rect 2057 1180 2071 1232
rect 2123 1180 2137 1232
rect 2189 1180 2203 1232
rect 2255 1180 2269 1232
rect 2321 1180 2334 1232
rect 2386 1180 2399 1232
rect 2451 1180 2464 1232
rect 2516 1180 2529 1232
rect 2581 1180 2594 1232
rect 2646 1180 2659 1232
rect 2711 1181 2723 1232
rect 2775 1182 2787 1233
rect 2839 1183 2851 1234
rect 2903 1184 2915 1235
rect 2967 1185 2979 1236
rect 3031 1186 3043 1237
rect 3095 1187 3107 1238
rect 3159 1187 3171 1239
rect 3095 1186 3223 1187
rect 3031 1185 3223 1186
rect 2967 1184 3223 1185
rect 2903 1183 3223 1184
rect 2839 1182 3223 1183
rect 2775 1181 3223 1182
rect 2711 1180 3223 1181
rect 1933 1174 3223 1180
rect 1933 1173 3107 1174
rect 1933 1172 3043 1173
rect 1933 1171 2979 1172
rect 1933 1170 2915 1171
rect 1933 1169 2851 1170
rect 1933 1168 2787 1169
rect 1933 1116 1939 1168
rect 1991 1116 2005 1168
rect 2057 1116 2071 1168
rect 2123 1116 2137 1168
rect 2189 1116 2203 1168
rect 2255 1116 2268 1168
rect 2320 1116 2333 1168
rect 2385 1116 2398 1168
rect 2450 1116 2463 1168
rect 2515 1116 2528 1168
rect 2580 1116 2593 1168
rect 2645 1116 2658 1168
rect 2710 1116 2723 1168
rect 2775 1117 2787 1168
rect 2839 1118 2851 1169
rect 2903 1119 2915 1170
rect 2967 1120 2979 1171
rect 3031 1121 3043 1172
rect 3095 1122 3107 1173
rect 3159 1122 3171 1174
rect 3095 1121 3223 1122
rect 3031 1120 3223 1121
rect 2967 1119 3223 1120
rect 2903 1118 3223 1119
rect 2839 1117 3223 1118
rect 2775 1116 3223 1117
rect 1933 1109 3223 1116
rect 1933 1108 3107 1109
rect 1933 1107 3043 1108
rect 1933 1106 2979 1107
rect 1933 1105 2915 1106
rect 1933 1104 2851 1105
rect 1933 1052 1939 1104
rect 1991 1052 2005 1104
rect 2057 1052 2071 1104
rect 2123 1052 2137 1104
rect 2189 1052 2202 1104
rect 2254 1052 2267 1104
rect 2319 1052 2332 1104
rect 2384 1052 2397 1104
rect 2449 1052 2462 1104
rect 2514 1052 2527 1104
rect 2579 1052 2592 1104
rect 2644 1052 2657 1104
rect 2709 1052 2722 1104
rect 2774 1052 2787 1104
rect 2839 1053 2851 1104
rect 2903 1054 2915 1105
rect 2967 1055 2979 1106
rect 3031 1056 3043 1107
rect 3095 1057 3107 1108
rect 3159 1057 3171 1109
rect 3095 1056 3223 1057
rect 3031 1055 3223 1056
rect 2967 1054 3223 1055
rect 2903 1053 3223 1054
rect 2839 1052 3223 1053
rect 1933 1044 3223 1052
rect 1933 1043 3107 1044
rect 1933 1042 3043 1043
rect 1933 1041 2979 1042
rect 1933 1040 2915 1041
rect 1933 988 1939 1040
rect 1991 988 2005 1040
rect 2057 988 2071 1040
rect 2123 988 2136 1040
rect 2188 988 2201 1040
rect 2253 988 2266 1040
rect 2318 988 2331 1040
rect 2383 988 2396 1040
rect 2448 988 2461 1040
rect 2513 988 2526 1040
rect 2578 988 2591 1040
rect 2643 988 2656 1040
rect 2708 988 2721 1040
rect 2773 988 2786 1040
rect 2838 988 2851 1040
rect 2903 989 2915 1040
rect 2967 990 2979 1041
rect 3031 991 3043 1042
rect 3095 992 3107 1043
rect 3159 992 3171 1044
rect 3526 1902 3824 1908
rect 3578 1850 3608 1902
rect 3660 1850 3690 1902
rect 3742 1850 3772 1902
rect 3526 1834 3824 1850
rect 3578 1782 3608 1834
rect 3660 1782 3690 1834
rect 3742 1782 3772 1834
rect 3526 1766 3824 1782
rect 3578 1714 3608 1766
rect 3660 1714 3690 1766
rect 3742 1714 3772 1766
rect 3526 1698 3824 1714
rect 3578 1646 3608 1698
rect 3660 1646 3690 1698
rect 3742 1646 3772 1698
rect 3526 1630 3824 1646
rect 3578 1578 3608 1630
rect 3660 1578 3690 1630
rect 3742 1578 3772 1630
rect 3526 1562 3824 1578
rect 3578 1510 3608 1562
rect 3660 1510 3690 1562
rect 3742 1510 3772 1562
rect 3526 1494 3824 1510
rect 3578 1442 3608 1494
rect 3660 1442 3690 1494
rect 3742 1442 3772 1494
rect 3526 1426 3824 1442
rect 3578 1374 3608 1426
rect 3660 1374 3690 1426
rect 3742 1374 3772 1426
rect 3526 1358 3824 1374
rect 3578 1306 3608 1358
rect 3660 1306 3690 1358
rect 3742 1306 3772 1358
rect 3526 1289 3824 1306
rect 3578 1237 3608 1289
rect 3660 1237 3690 1289
rect 3742 1237 3772 1289
rect 3526 1220 3824 1237
rect 3578 1168 3608 1220
rect 3660 1168 3690 1220
rect 3742 1168 3772 1220
rect 3526 1151 3824 1168
rect 3578 1099 3608 1151
rect 3660 1099 3690 1151
rect 3742 1099 3772 1151
rect 3526 1082 3824 1099
rect 3578 1030 3608 1082
rect 3660 1030 3690 1082
rect 3742 1030 3772 1082
rect 3526 1024 3824 1030
rect 4349 1902 4649 1908
rect 4349 1850 4350 1902
rect 4402 1850 4432 1902
rect 4484 1850 4514 1902
rect 4566 1850 4596 1902
rect 4648 1850 4649 1902
rect 4349 1838 4649 1850
rect 4349 1786 4350 1838
rect 4402 1786 4432 1838
rect 4484 1786 4514 1838
rect 4566 1786 4596 1838
rect 4648 1786 4649 1838
rect 4349 1774 4649 1786
rect 4349 1722 4350 1774
rect 4402 1722 4432 1774
rect 4484 1722 4514 1774
rect 4566 1722 4596 1774
rect 4648 1722 4649 1774
rect 4349 1710 4649 1722
rect 4349 1658 4350 1710
rect 4402 1658 4432 1710
rect 4484 1658 4514 1710
rect 4566 1658 4596 1710
rect 4648 1658 4649 1710
rect 4349 1646 4649 1658
rect 4349 1594 4350 1646
rect 4402 1594 4432 1646
rect 4484 1594 4514 1646
rect 4566 1594 4596 1646
rect 4648 1594 4649 1646
rect 4349 1582 4649 1594
rect 4349 1530 4350 1582
rect 4402 1530 4432 1582
rect 4484 1530 4514 1582
rect 4566 1530 4596 1582
rect 4648 1530 4649 1582
rect 4349 1518 4649 1530
rect 4349 1466 4350 1518
rect 4402 1466 4432 1518
rect 4484 1466 4514 1518
rect 4566 1466 4596 1518
rect 4648 1466 4649 1518
rect 4349 1454 4649 1466
rect 4349 1402 4350 1454
rect 4402 1402 4432 1454
rect 4484 1402 4514 1454
rect 4566 1402 4596 1454
rect 4648 1402 4649 1454
rect 4349 1390 4649 1402
rect 4349 1338 4350 1390
rect 4402 1338 4432 1390
rect 4484 1338 4514 1390
rect 4566 1338 4596 1390
rect 4648 1338 4649 1390
rect 4349 1326 4649 1338
rect 4349 1274 4350 1326
rect 4402 1274 4432 1326
rect 4484 1274 4514 1326
rect 4566 1274 4596 1326
rect 4648 1274 4649 1326
rect 4349 1262 4649 1274
rect 4349 1210 4350 1262
rect 4402 1210 4432 1262
rect 4484 1210 4514 1262
rect 4566 1210 4596 1262
rect 4648 1210 4649 1262
rect 4349 1198 4649 1210
rect 4349 1146 4350 1198
rect 4402 1146 4432 1198
rect 4484 1146 4514 1198
rect 4566 1146 4596 1198
rect 4648 1146 4649 1198
rect 4349 1134 4649 1146
rect 4349 1082 4350 1134
rect 4402 1082 4432 1134
rect 4484 1082 4514 1134
rect 4566 1082 4596 1134
rect 4648 1082 4649 1134
rect 4349 1070 4649 1082
rect 4349 1018 4350 1070
rect 4402 1018 4432 1070
rect 4484 1018 4514 1070
rect 4566 1018 4596 1070
rect 4648 1018 4649 1070
rect 3095 991 3223 992
rect 3031 990 3223 991
rect 2967 989 3223 990
rect 2903 988 3223 989
rect 1933 979 3223 988
rect 1933 978 3107 979
rect 1933 977 3043 978
rect 1933 976 2979 977
rect 1933 924 1939 976
rect 1991 924 2005 976
rect 2057 924 2070 976
rect 2122 924 2135 976
rect 2187 924 2200 976
rect 2252 924 2265 976
rect 2317 924 2330 976
rect 2382 924 2395 976
rect 2447 924 2460 976
rect 2512 924 2525 976
rect 2577 924 2590 976
rect 2642 924 2655 976
rect 2707 924 2720 976
rect 2772 924 2785 976
rect 2837 924 2850 976
rect 2902 924 2915 976
rect 2967 925 2979 976
rect 3031 926 3043 977
rect 3095 927 3107 978
rect 3159 927 3171 979
rect 3584 966 3590 1018
rect 3642 966 3678 1018
rect 3730 966 3766 1018
rect 3818 966 3824 1018
rect 4349 1006 4649 1018
rect 4349 954 4350 1006
rect 4402 954 4432 1006
rect 4484 954 4514 1006
rect 4566 954 4596 1006
rect 4648 954 4649 1006
rect 3095 926 3223 927
rect 3031 925 3223 926
rect 2967 924 3223 925
rect 1933 914 3223 924
rect 1933 913 3107 914
rect 1933 912 3043 913
rect 1933 860 1939 912
rect 1991 860 2004 912
rect 2056 860 2069 912
rect 2121 860 2134 912
rect 2186 860 2199 912
rect 2251 860 2264 912
rect 2316 860 2329 912
rect 2381 860 2394 912
rect 2446 860 2459 912
rect 2511 860 2524 912
rect 2576 860 2589 912
rect 2641 860 2654 912
rect 2706 860 2719 912
rect 2771 860 2784 912
rect 2836 860 2849 912
rect 2901 860 2914 912
rect 2966 860 2979 912
rect 3031 861 3043 912
rect 3095 862 3107 913
rect 3159 862 3171 914
rect 3654 901 3660 953
rect 3712 901 3766 953
rect 3818 901 3824 953
rect 4349 942 4649 954
rect 4349 890 4350 942
rect 4402 890 4432 942
rect 4484 890 4514 942
rect 4566 890 4596 942
rect 4648 890 4649 942
rect 4349 878 4649 890
rect 3095 861 3223 862
rect 3031 860 3223 861
rect 1933 849 3223 860
rect 1933 848 3107 849
rect 1933 796 1939 848
rect 1991 796 2004 848
rect 2056 796 2069 848
rect 2121 796 2134 848
rect 2186 796 2199 848
rect 2251 796 2264 848
rect 2316 796 2329 848
rect 2381 796 2394 848
rect 2446 796 2459 848
rect 2511 796 2524 848
rect 2576 796 2589 848
rect 2641 796 2654 848
rect 2706 796 2719 848
rect 2771 796 2784 848
rect 2836 796 2849 848
rect 2901 796 2914 848
rect 2966 796 2979 848
rect 1933 784 2979 796
rect 3095 797 3107 848
rect 3159 797 3171 849
rect 3747 815 3753 867
rect 3805 815 3816 867
rect 4349 826 4350 878
rect 4402 826 4432 878
rect 4484 826 4514 878
rect 4566 826 4596 878
rect 4648 826 4649 878
rect 3095 784 3223 797
rect 1933 732 1939 784
rect 1991 732 2004 784
rect 2056 732 2069 784
rect 2121 732 2134 784
rect 2186 732 2199 784
rect 2251 732 2264 784
rect 2316 732 2329 784
rect 2381 732 2394 784
rect 2446 732 2459 784
rect 2511 732 2524 784
rect 2576 732 2589 784
rect 2641 732 2654 784
rect 2706 732 2719 784
rect 2771 732 2784 784
rect 2836 732 2849 784
rect 2901 732 2914 784
rect 2966 732 2979 784
rect 1933 720 2979 732
rect 1933 668 1939 720
rect 1991 668 2004 720
rect 2056 668 2069 720
rect 2121 668 2134 720
rect 2186 668 2199 720
rect 2251 668 2264 720
rect 2316 668 2329 720
rect 2381 668 2394 720
rect 2446 668 2459 720
rect 2511 668 2524 720
rect 2576 668 2589 720
rect 2641 668 2654 720
rect 2706 668 2719 720
rect 2771 668 2784 720
rect 2836 668 2849 720
rect 2901 668 2914 720
rect 2966 668 2979 720
rect 3159 732 3171 784
rect 3159 668 3223 732
rect 4349 814 4649 826
rect 4349 762 4350 814
rect 4402 762 4432 814
rect 4484 762 4514 814
rect 4566 762 4596 814
rect 4648 762 4649 814
rect 4349 750 4649 762
rect 4349 698 4350 750
rect 4402 698 4432 750
rect 4484 698 4514 750
rect 4566 698 4596 750
rect 4648 698 4649 750
rect 4349 685 4649 698
tri 1825 656 1827 658 sw
rect 1711 652 1827 656
rect 1671 649 1827 652
tri 1827 649 1834 656 sw
rect 1671 615 1785 649
rect 1819 644 1834 649
tri 1834 644 1839 649 sw
rect 1819 619 1839 644
tri 1839 619 1864 644 sw
tri 3306 619 3331 644 se
rect 1819 615 1864 619
rect 1671 613 1864 615
rect 1671 579 1677 613
rect 1711 594 1864 613
tri 1864 594 1889 619 sw
tri 3281 594 3306 619 se
rect 3306 609 3331 619
rect 4349 633 4350 685
rect 4402 633 4432 685
rect 4484 633 4514 685
rect 4566 633 4596 685
rect 4648 633 4649 685
rect 4349 620 4649 633
rect 3306 594 3413 609
rect 1711 588 1889 594
tri 1889 588 1895 594 sw
tri 3275 588 3281 594 se
rect 3281 588 3413 594
rect 1711 584 3413 588
tri 3516 585 3525 594 se
tri 3515 584 3516 585 se
rect 3516 584 3525 585
rect 1711 582 3403 584
rect 1711 579 1892 582
rect 1671 576 1892 579
rect 1671 542 1785 576
rect 1819 548 1892 576
rect 1926 548 1967 582
rect 2001 548 2042 582
rect 2076 548 2117 582
rect 2151 548 2192 582
rect 2226 548 2266 582
rect 2300 548 2340 582
rect 2374 548 2414 582
rect 2448 548 2488 582
rect 2522 548 2562 582
rect 2596 548 2636 582
rect 2670 548 2710 582
rect 2744 548 2784 582
rect 2818 548 2858 582
rect 2892 548 2932 582
rect 2966 548 3006 582
rect 3040 548 3080 582
rect 3114 548 3154 582
rect 3188 548 3228 582
rect 3262 574 3403 582
tri 3403 574 3413 584 nw
tri 3505 574 3515 584 se
rect 3515 574 3525 584
rect 3262 548 3373 574
rect 1819 544 3373 548
tri 3373 544 3403 574 nw
tri 3475 544 3505 574 se
rect 3505 544 3525 574
rect 1819 542 3339 544
rect 1671 540 3339 542
rect 1671 506 1677 540
rect 1711 510 3339 540
tri 3339 510 3373 544 nw
tri 3441 510 3475 544 se
rect 3475 510 3525 544
rect 1711 506 1892 510
rect 1671 503 1892 506
rect 1671 469 1785 503
rect 1819 476 1892 503
rect 1926 476 1967 510
rect 2001 476 2042 510
rect 2076 476 2117 510
rect 2151 476 2192 510
rect 2226 476 2266 510
rect 2300 476 2340 510
rect 2374 476 2414 510
rect 2448 476 2488 510
rect 2522 476 2562 510
rect 2596 476 2636 510
rect 2670 476 2710 510
rect 2744 476 2784 510
rect 2818 476 2858 510
rect 2892 476 2932 510
rect 2966 476 3006 510
rect 3040 476 3080 510
rect 3114 476 3154 510
rect 3188 476 3228 510
rect 3262 499 3328 510
tri 3328 499 3339 510 nw
tri 3430 499 3441 510 se
rect 3441 499 3525 510
rect 3262 482 3311 499
tri 3311 482 3328 499 nw
tri 3413 482 3430 499 se
rect 3430 482 3525 499
rect 3262 476 3299 482
rect 1819 470 3299 476
tri 3299 470 3311 482 nw
tri 3401 470 3413 482 se
rect 3413 470 3525 482
rect 1819 469 3297 470
rect 1671 468 3297 469
tri 3297 468 3299 470 nw
tri 3399 468 3401 470 se
rect 3401 468 3525 470
rect 1671 467 3287 468
rect 1671 433 1677 467
rect 1711 458 3287 467
tri 3287 458 3297 468 nw
tri 3389 458 3399 468 se
rect 3399 458 3525 468
rect 1711 433 3276 458
tri 3276 447 3287 458 nw
tri 3378 447 3389 458 se
rect 3389 447 3525 458
rect 1671 430 3276 433
rect 1671 396 1785 430
rect 1819 396 1860 430
rect 1894 396 1935 430
rect 1969 396 2010 430
rect 2044 396 2085 430
rect 2119 396 2160 430
rect 2194 396 2235 430
rect 2269 396 2310 430
rect 2344 396 2385 430
rect 2419 396 2460 430
rect 2494 396 2535 430
rect 2569 396 2610 430
rect 2644 396 2685 430
rect 2719 396 2760 430
rect 2794 396 2835 430
rect 2869 396 2910 430
rect 2944 396 2985 430
rect 3019 396 3060 430
rect 3094 396 3135 430
rect 3169 396 3210 430
rect 3244 396 3276 430
tri 3355 424 3378 447 se
rect 3378 424 3525 447
tri 3331 400 3355 424 se
rect 3355 400 3525 424
rect 4349 568 4350 620
rect 4402 568 4432 620
rect 4484 568 4514 620
rect 4566 568 4596 620
rect 4648 568 4649 620
rect 4349 555 4649 568
rect 4349 503 4350 555
rect 4402 503 4432 555
rect 4484 503 4514 555
rect 4566 503 4596 555
rect 4648 503 4649 555
rect 4349 490 4649 503
rect 4349 438 4350 490
rect 4402 438 4432 490
rect 4484 438 4514 490
rect 4566 438 4596 490
rect 4648 438 4649 490
rect 4349 425 4649 438
rect 1671 394 3276 396
rect 1671 360 1677 394
rect 1711 360 3276 394
rect 4349 373 4350 425
rect 4402 373 4432 425
rect 4484 373 4514 425
rect 4566 373 4596 425
rect 4648 373 4649 425
rect 4349 367 4649 373
rect 5173 1902 5473 1908
rect 5173 1850 5174 1902
rect 5226 1850 5256 1902
rect 5308 1850 5338 1902
rect 5390 1850 5420 1902
rect 5472 1850 5473 1902
rect 5173 1838 5473 1850
rect 5173 1786 5174 1838
rect 5226 1786 5256 1838
rect 5308 1786 5338 1838
rect 5390 1786 5420 1838
rect 5472 1786 5473 1838
rect 5173 1774 5473 1786
rect 5173 1722 5174 1774
rect 5226 1722 5256 1774
rect 5308 1722 5338 1774
rect 5390 1722 5420 1774
rect 5472 1722 5473 1774
rect 5173 1710 5473 1722
rect 5173 1658 5174 1710
rect 5226 1658 5256 1710
rect 5308 1658 5338 1710
rect 5390 1658 5420 1710
rect 5472 1658 5473 1710
rect 5173 1646 5473 1658
rect 5173 1594 5174 1646
rect 5226 1594 5256 1646
rect 5308 1594 5338 1646
rect 5390 1594 5420 1646
rect 5472 1594 5473 1646
rect 5173 1582 5473 1594
rect 5173 1530 5174 1582
rect 5226 1530 5256 1582
rect 5308 1530 5338 1582
rect 5390 1530 5420 1582
rect 5472 1530 5473 1582
rect 5173 1518 5473 1530
rect 5173 1466 5174 1518
rect 5226 1466 5256 1518
rect 5308 1466 5338 1518
rect 5390 1466 5420 1518
rect 5472 1466 5473 1518
rect 5173 1454 5473 1466
rect 5173 1402 5174 1454
rect 5226 1402 5256 1454
rect 5308 1402 5338 1454
rect 5390 1402 5420 1454
rect 5472 1402 5473 1454
rect 5173 1390 5473 1402
rect 5173 1338 5174 1390
rect 5226 1338 5256 1390
rect 5308 1338 5338 1390
rect 5390 1338 5420 1390
rect 5472 1338 5473 1390
rect 5173 1326 5473 1338
rect 5173 1274 5174 1326
rect 5226 1274 5256 1326
rect 5308 1274 5338 1326
rect 5390 1274 5420 1326
rect 5472 1274 5473 1326
rect 5173 1262 5473 1274
rect 5173 1210 5174 1262
rect 5226 1210 5256 1262
rect 5308 1210 5338 1262
rect 5390 1210 5420 1262
rect 5472 1210 5473 1262
rect 5173 1198 5473 1210
rect 5173 1146 5174 1198
rect 5226 1146 5256 1198
rect 5308 1146 5338 1198
rect 5390 1146 5420 1198
rect 5472 1146 5473 1198
rect 5173 1134 5473 1146
rect 5173 1082 5174 1134
rect 5226 1082 5256 1134
rect 5308 1082 5338 1134
rect 5390 1082 5420 1134
rect 5472 1082 5473 1134
rect 5173 1070 5473 1082
rect 5173 1018 5174 1070
rect 5226 1018 5256 1070
rect 5308 1018 5338 1070
rect 5390 1018 5420 1070
rect 5472 1018 5473 1070
rect 5173 1006 5473 1018
rect 5173 954 5174 1006
rect 5226 954 5256 1006
rect 5308 954 5338 1006
rect 5390 954 5420 1006
rect 5472 954 5473 1006
rect 5173 942 5473 954
rect 5173 890 5174 942
rect 5226 890 5256 942
rect 5308 890 5338 942
rect 5390 890 5420 942
rect 5472 890 5473 942
rect 5173 878 5473 890
rect 5173 826 5174 878
rect 5226 826 5256 878
rect 5308 826 5338 878
rect 5390 826 5420 878
rect 5472 826 5473 878
rect 5173 814 5473 826
rect 5173 762 5174 814
rect 5226 762 5256 814
rect 5308 762 5338 814
rect 5390 762 5420 814
rect 5472 762 5473 814
rect 5173 750 5473 762
rect 5173 698 5174 750
rect 5226 698 5256 750
rect 5308 698 5338 750
rect 5390 698 5420 750
rect 5472 698 5473 750
rect 5173 685 5473 698
rect 5173 633 5174 685
rect 5226 633 5256 685
rect 5308 633 5338 685
rect 5390 633 5420 685
rect 5472 633 5473 685
rect 5173 620 5473 633
rect 5173 568 5174 620
rect 5226 568 5256 620
rect 5308 568 5338 620
rect 5390 568 5420 620
rect 5472 568 5473 620
rect 5173 555 5473 568
rect 5173 503 5174 555
rect 5226 503 5256 555
rect 5308 503 5338 555
rect 5390 503 5420 555
rect 5472 503 5473 555
rect 5173 490 5473 503
rect 5173 438 5174 490
rect 5226 438 5256 490
rect 5308 438 5338 490
rect 5390 438 5420 490
rect 5472 438 5473 490
rect 5173 425 5473 438
rect 5173 373 5174 425
rect 5226 373 5256 425
rect 5308 373 5338 425
rect 5390 373 5420 425
rect 5472 373 5473 425
rect 5173 367 5473 373
rect 5997 1902 6297 1908
rect 5997 1850 5998 1902
rect 6050 1850 6080 1902
rect 6132 1850 6162 1902
rect 6214 1850 6244 1902
rect 6296 1850 6297 1902
rect 5997 1838 6297 1850
rect 5997 1786 5998 1838
rect 6050 1786 6080 1838
rect 6132 1786 6162 1838
rect 6214 1786 6244 1838
rect 6296 1786 6297 1838
rect 5997 1774 6297 1786
rect 5997 1722 5998 1774
rect 6050 1722 6080 1774
rect 6132 1722 6162 1774
rect 6214 1722 6244 1774
rect 6296 1722 6297 1774
rect 5997 1710 6297 1722
rect 5997 1658 5998 1710
rect 6050 1658 6080 1710
rect 6132 1658 6162 1710
rect 6214 1658 6244 1710
rect 6296 1658 6297 1710
rect 5997 1646 6297 1658
rect 5997 1594 5998 1646
rect 6050 1594 6080 1646
rect 6132 1594 6162 1646
rect 6214 1594 6244 1646
rect 6296 1594 6297 1646
rect 5997 1582 6297 1594
rect 5997 1530 5998 1582
rect 6050 1530 6080 1582
rect 6132 1530 6162 1582
rect 6214 1530 6244 1582
rect 6296 1530 6297 1582
rect 5997 1518 6297 1530
rect 5997 1466 5998 1518
rect 6050 1466 6080 1518
rect 6132 1466 6162 1518
rect 6214 1466 6244 1518
rect 6296 1466 6297 1518
rect 5997 1454 6297 1466
rect 5997 1402 5998 1454
rect 6050 1402 6080 1454
rect 6132 1402 6162 1454
rect 6214 1402 6244 1454
rect 6296 1402 6297 1454
rect 5997 1390 6297 1402
rect 5997 1338 5998 1390
rect 6050 1338 6080 1390
rect 6132 1338 6162 1390
rect 6214 1338 6244 1390
rect 6296 1338 6297 1390
rect 5997 1326 6297 1338
rect 5997 1274 5998 1326
rect 6050 1274 6080 1326
rect 6132 1274 6162 1326
rect 6214 1274 6244 1326
rect 6296 1274 6297 1326
rect 5997 1262 6297 1274
rect 5997 1210 5998 1262
rect 6050 1210 6080 1262
rect 6132 1210 6162 1262
rect 6214 1210 6244 1262
rect 6296 1210 6297 1262
rect 5997 1198 6297 1210
rect 5997 1146 5998 1198
rect 6050 1146 6080 1198
rect 6132 1146 6162 1198
rect 6214 1146 6244 1198
rect 6296 1146 6297 1198
rect 5997 1134 6297 1146
rect 5997 1082 5998 1134
rect 6050 1082 6080 1134
rect 6132 1082 6162 1134
rect 6214 1082 6244 1134
rect 6296 1082 6297 1134
rect 5997 1070 6297 1082
rect 5997 1018 5998 1070
rect 6050 1018 6080 1070
rect 6132 1018 6162 1070
rect 6214 1018 6244 1070
rect 6296 1018 6297 1070
rect 5997 1006 6297 1018
rect 5997 954 5998 1006
rect 6050 954 6080 1006
rect 6132 954 6162 1006
rect 6214 954 6244 1006
rect 6296 954 6297 1006
rect 5997 942 6297 954
rect 5997 890 5998 942
rect 6050 890 6080 942
rect 6132 890 6162 942
rect 6214 890 6244 942
rect 6296 890 6297 942
rect 5997 878 6297 890
rect 5997 826 5998 878
rect 6050 826 6080 878
rect 6132 826 6162 878
rect 6214 826 6244 878
rect 6296 826 6297 878
rect 5997 814 6297 826
rect 5997 762 5998 814
rect 6050 762 6080 814
rect 6132 762 6162 814
rect 6214 762 6244 814
rect 6296 762 6297 814
rect 5997 750 6297 762
rect 5997 698 5998 750
rect 6050 698 6080 750
rect 6132 698 6162 750
rect 6214 698 6244 750
rect 6296 698 6297 750
rect 5997 685 6297 698
rect 5997 633 5998 685
rect 6050 633 6080 685
rect 6132 633 6162 685
rect 6214 633 6244 685
rect 6296 633 6297 685
rect 5997 620 6297 633
rect 5997 568 5998 620
rect 6050 568 6080 620
rect 6132 568 6162 620
rect 6214 568 6244 620
rect 6296 568 6297 620
rect 5997 555 6297 568
rect 5997 503 5998 555
rect 6050 503 6080 555
rect 6132 503 6162 555
rect 6214 503 6244 555
rect 6296 503 6297 555
rect 5997 490 6297 503
rect 5997 438 5998 490
rect 6050 438 6080 490
rect 6132 438 6162 490
rect 6214 438 6244 490
rect 6296 438 6297 490
rect 5997 425 6297 438
rect 5997 373 5998 425
rect 6050 373 6080 425
rect 6132 373 6162 425
rect 6214 373 6244 425
rect 6296 373 6297 425
rect 5997 367 6297 373
rect 6821 1902 7121 1908
rect 6821 1850 6822 1902
rect 6874 1850 6904 1902
rect 6956 1850 6986 1902
rect 7038 1850 7068 1902
rect 7120 1850 7121 1902
rect 6821 1838 7121 1850
rect 6821 1786 6822 1838
rect 6874 1786 6904 1838
rect 6956 1786 6986 1838
rect 7038 1786 7068 1838
rect 7120 1786 7121 1838
rect 6821 1774 7121 1786
rect 6821 1722 6822 1774
rect 6874 1722 6904 1774
rect 6956 1722 6986 1774
rect 7038 1722 7068 1774
rect 7120 1722 7121 1774
rect 6821 1710 7121 1722
rect 6821 1658 6822 1710
rect 6874 1658 6904 1710
rect 6956 1658 6986 1710
rect 7038 1658 7068 1710
rect 7120 1658 7121 1710
rect 6821 1646 7121 1658
rect 6821 1594 6822 1646
rect 6874 1594 6904 1646
rect 6956 1594 6986 1646
rect 7038 1594 7068 1646
rect 7120 1594 7121 1646
rect 6821 1582 7121 1594
rect 6821 1530 6822 1582
rect 6874 1530 6904 1582
rect 6956 1530 6986 1582
rect 7038 1530 7068 1582
rect 7120 1530 7121 1582
rect 6821 1518 7121 1530
rect 6821 1466 6822 1518
rect 6874 1466 6904 1518
rect 6956 1466 6986 1518
rect 7038 1466 7068 1518
rect 7120 1466 7121 1518
rect 6821 1454 7121 1466
rect 6821 1402 6822 1454
rect 6874 1402 6904 1454
rect 6956 1402 6986 1454
rect 7038 1402 7068 1454
rect 7120 1402 7121 1454
rect 6821 1390 7121 1402
rect 6821 1338 6822 1390
rect 6874 1338 6904 1390
rect 6956 1338 6986 1390
rect 7038 1338 7068 1390
rect 7120 1338 7121 1390
rect 6821 1326 7121 1338
rect 6821 1274 6822 1326
rect 6874 1274 6904 1326
rect 6956 1274 6986 1326
rect 7038 1274 7068 1326
rect 7120 1274 7121 1326
rect 6821 1262 7121 1274
rect 6821 1210 6822 1262
rect 6874 1210 6904 1262
rect 6956 1210 6986 1262
rect 7038 1210 7068 1262
rect 7120 1210 7121 1262
rect 6821 1198 7121 1210
rect 6821 1146 6822 1198
rect 6874 1146 6904 1198
rect 6956 1146 6986 1198
rect 7038 1146 7068 1198
rect 7120 1146 7121 1198
rect 6821 1134 7121 1146
rect 6821 1082 6822 1134
rect 6874 1082 6904 1134
rect 6956 1082 6986 1134
rect 7038 1082 7068 1134
rect 7120 1082 7121 1134
rect 6821 1070 7121 1082
rect 6821 1018 6822 1070
rect 6874 1018 6904 1070
rect 6956 1018 6986 1070
rect 7038 1018 7068 1070
rect 7120 1018 7121 1070
rect 6821 1006 7121 1018
rect 6821 954 6822 1006
rect 6874 954 6904 1006
rect 6956 954 6986 1006
rect 7038 954 7068 1006
rect 7120 954 7121 1006
rect 6821 942 7121 954
rect 6821 890 6822 942
rect 6874 890 6904 942
rect 6956 890 6986 942
rect 7038 890 7068 942
rect 7120 890 7121 942
rect 6821 878 7121 890
rect 6821 826 6822 878
rect 6874 826 6904 878
rect 6956 826 6986 878
rect 7038 826 7068 878
rect 7120 826 7121 878
rect 6821 814 7121 826
rect 6821 762 6822 814
rect 6874 762 6904 814
rect 6956 762 6986 814
rect 7038 762 7068 814
rect 7120 762 7121 814
rect 6821 750 7121 762
rect 6821 698 6822 750
rect 6874 698 6904 750
rect 6956 698 6986 750
rect 7038 698 7068 750
rect 7120 698 7121 750
rect 6821 685 7121 698
rect 6821 633 6822 685
rect 6874 633 6904 685
rect 6956 633 6986 685
rect 7038 633 7068 685
rect 7120 633 7121 685
rect 6821 620 7121 633
rect 6821 568 6822 620
rect 6874 568 6904 620
rect 6956 568 6986 620
rect 7038 568 7068 620
rect 7120 568 7121 620
rect 6821 555 7121 568
rect 6821 503 6822 555
rect 6874 503 6904 555
rect 6956 503 6986 555
rect 7038 503 7068 555
rect 7120 503 7121 555
rect 6821 490 7121 503
rect 6821 438 6822 490
rect 6874 438 6904 490
rect 6956 438 6986 490
rect 7038 438 7068 490
rect 7120 438 7121 490
rect 6821 425 7121 438
rect 6821 373 6822 425
rect 6874 373 6904 425
rect 6956 373 6986 425
rect 7038 373 7068 425
rect 7120 373 7121 425
rect 6821 367 7121 373
rect 7935 1902 8235 1908
rect 7935 1850 7936 1902
rect 7988 1850 8018 1902
rect 8070 1850 8100 1902
rect 8152 1850 8182 1902
rect 8234 1850 8235 1902
rect 7935 1838 8235 1850
rect 7935 1786 7936 1838
rect 7988 1786 8018 1838
rect 8070 1786 8100 1838
rect 8152 1786 8182 1838
rect 8234 1786 8235 1838
rect 7935 1774 8235 1786
rect 7935 1722 7936 1774
rect 7988 1722 8018 1774
rect 8070 1722 8100 1774
rect 8152 1722 8182 1774
rect 8234 1722 8235 1774
rect 7935 1710 8235 1722
rect 7935 1658 7936 1710
rect 7988 1658 8018 1710
rect 8070 1658 8100 1710
rect 8152 1658 8182 1710
rect 8234 1658 8235 1710
rect 7935 1646 8235 1658
rect 7935 1594 7936 1646
rect 7988 1594 8018 1646
rect 8070 1594 8100 1646
rect 8152 1594 8182 1646
rect 8234 1594 8235 1646
rect 7935 1582 8235 1594
rect 7935 1530 7936 1582
rect 7988 1530 8018 1582
rect 8070 1530 8100 1582
rect 8152 1530 8182 1582
rect 8234 1530 8235 1582
rect 7935 1518 8235 1530
rect 7935 1466 7936 1518
rect 7988 1466 8018 1518
rect 8070 1466 8100 1518
rect 8152 1466 8182 1518
rect 8234 1466 8235 1518
rect 7935 1454 8235 1466
rect 7935 1402 7936 1454
rect 7988 1402 8018 1454
rect 8070 1402 8100 1454
rect 8152 1402 8182 1454
rect 8234 1402 8235 1454
rect 7935 1390 8235 1402
rect 7935 1338 7936 1390
rect 7988 1338 8018 1390
rect 8070 1338 8100 1390
rect 8152 1338 8182 1390
rect 8234 1338 8235 1390
rect 7935 1326 8235 1338
rect 7935 1274 7936 1326
rect 7988 1274 8018 1326
rect 8070 1274 8100 1326
rect 8152 1274 8182 1326
rect 8234 1274 8235 1326
rect 7935 1262 8235 1274
rect 7935 1210 7936 1262
rect 7988 1210 8018 1262
rect 8070 1210 8100 1262
rect 8152 1210 8182 1262
rect 8234 1210 8235 1262
rect 7935 1198 8235 1210
rect 7935 1146 7936 1198
rect 7988 1146 8018 1198
rect 8070 1146 8100 1198
rect 8152 1146 8182 1198
rect 8234 1146 8235 1198
rect 7935 1134 8235 1146
rect 7935 1082 7936 1134
rect 7988 1082 8018 1134
rect 8070 1082 8100 1134
rect 8152 1082 8182 1134
rect 8234 1082 8235 1134
rect 7935 1070 8235 1082
rect 7935 1018 7936 1070
rect 7988 1018 8018 1070
rect 8070 1018 8100 1070
rect 8152 1018 8182 1070
rect 8234 1018 8235 1070
rect 7935 1006 8235 1018
rect 7935 954 7936 1006
rect 7988 954 8018 1006
rect 8070 954 8100 1006
rect 8152 954 8182 1006
rect 8234 954 8235 1006
rect 7935 942 8235 954
rect 7935 890 7936 942
rect 7988 890 8018 942
rect 8070 890 8100 942
rect 8152 890 8182 942
rect 8234 890 8235 942
rect 7935 878 8235 890
rect 7935 826 7936 878
rect 7988 826 8018 878
rect 8070 826 8100 878
rect 8152 826 8182 878
rect 8234 826 8235 878
rect 7935 814 8235 826
rect 7935 762 7936 814
rect 7988 762 8018 814
rect 8070 762 8100 814
rect 8152 762 8182 814
rect 8234 762 8235 814
rect 7935 750 8235 762
rect 7935 698 7936 750
rect 7988 698 8018 750
rect 8070 698 8100 750
rect 8152 698 8182 750
rect 8234 698 8235 750
rect 7935 685 8235 698
rect 7935 633 7936 685
rect 7988 633 8018 685
rect 8070 633 8100 685
rect 8152 633 8182 685
rect 8234 633 8235 685
rect 7935 620 8235 633
rect 7935 568 7936 620
rect 7988 568 8018 620
rect 8070 568 8100 620
rect 8152 568 8182 620
rect 8234 568 8235 620
rect 7935 555 8235 568
rect 7935 503 7936 555
rect 7988 503 8018 555
rect 8070 503 8100 555
rect 8152 503 8182 555
rect 8234 503 8235 555
rect 7935 490 8235 503
rect 7935 438 7936 490
rect 7988 438 8018 490
rect 8070 438 8100 490
rect 8152 438 8182 490
rect 8234 438 8235 490
rect 7935 425 8235 438
rect 7935 373 7936 425
rect 7988 373 8018 425
rect 8070 373 8100 425
rect 8152 373 8182 425
rect 8234 373 8235 425
rect 7935 367 8235 373
rect 8759 1902 9059 1908
rect 8759 1850 8760 1902
rect 8812 1850 8842 1902
rect 8894 1850 8924 1902
rect 8976 1850 9006 1902
rect 9058 1850 9059 1902
rect 8759 1838 9059 1850
rect 8759 1786 8760 1838
rect 8812 1786 8842 1838
rect 8894 1786 8924 1838
rect 8976 1786 9006 1838
rect 9058 1786 9059 1838
rect 8759 1774 9059 1786
rect 8759 1722 8760 1774
rect 8812 1722 8842 1774
rect 8894 1722 8924 1774
rect 8976 1722 9006 1774
rect 9058 1722 9059 1774
rect 8759 1710 9059 1722
rect 8759 1658 8760 1710
rect 8812 1658 8842 1710
rect 8894 1658 8924 1710
rect 8976 1658 9006 1710
rect 9058 1658 9059 1710
rect 8759 1646 9059 1658
rect 8759 1594 8760 1646
rect 8812 1594 8842 1646
rect 8894 1594 8924 1646
rect 8976 1594 9006 1646
rect 9058 1594 9059 1646
rect 8759 1582 9059 1594
rect 8759 1530 8760 1582
rect 8812 1530 8842 1582
rect 8894 1530 8924 1582
rect 8976 1530 9006 1582
rect 9058 1530 9059 1582
rect 8759 1518 9059 1530
rect 8759 1466 8760 1518
rect 8812 1466 8842 1518
rect 8894 1466 8924 1518
rect 8976 1466 9006 1518
rect 9058 1466 9059 1518
rect 8759 1454 9059 1466
rect 8759 1402 8760 1454
rect 8812 1402 8842 1454
rect 8894 1402 8924 1454
rect 8976 1402 9006 1454
rect 9058 1402 9059 1454
rect 8759 1390 9059 1402
rect 8759 1338 8760 1390
rect 8812 1338 8842 1390
rect 8894 1338 8924 1390
rect 8976 1338 9006 1390
rect 9058 1338 9059 1390
rect 8759 1326 9059 1338
rect 8759 1274 8760 1326
rect 8812 1274 8842 1326
rect 8894 1274 8924 1326
rect 8976 1274 9006 1326
rect 9058 1274 9059 1326
rect 8759 1262 9059 1274
rect 8759 1210 8760 1262
rect 8812 1210 8842 1262
rect 8894 1210 8924 1262
rect 8976 1210 9006 1262
rect 9058 1210 9059 1262
rect 8759 1198 9059 1210
rect 8759 1146 8760 1198
rect 8812 1146 8842 1198
rect 8894 1146 8924 1198
rect 8976 1146 9006 1198
rect 9058 1146 9059 1198
rect 8759 1134 9059 1146
rect 8759 1082 8760 1134
rect 8812 1082 8842 1134
rect 8894 1082 8924 1134
rect 8976 1082 9006 1134
rect 9058 1082 9059 1134
rect 8759 1070 9059 1082
rect 8759 1018 8760 1070
rect 8812 1018 8842 1070
rect 8894 1018 8924 1070
rect 8976 1018 9006 1070
rect 9058 1018 9059 1070
rect 8759 1006 9059 1018
rect 8759 954 8760 1006
rect 8812 954 8842 1006
rect 8894 954 8924 1006
rect 8976 954 9006 1006
rect 9058 954 9059 1006
rect 8759 942 9059 954
rect 8759 890 8760 942
rect 8812 890 8842 942
rect 8894 890 8924 942
rect 8976 890 9006 942
rect 9058 890 9059 942
rect 8759 878 9059 890
rect 8759 826 8760 878
rect 8812 826 8842 878
rect 8894 826 8924 878
rect 8976 826 9006 878
rect 9058 826 9059 878
rect 8759 814 9059 826
rect 8759 762 8760 814
rect 8812 762 8842 814
rect 8894 762 8924 814
rect 8976 762 9006 814
rect 9058 762 9059 814
rect 8759 750 9059 762
rect 8759 698 8760 750
rect 8812 698 8842 750
rect 8894 698 8924 750
rect 8976 698 9006 750
rect 9058 698 9059 750
rect 8759 685 9059 698
rect 8759 633 8760 685
rect 8812 633 8842 685
rect 8894 633 8924 685
rect 8976 633 9006 685
rect 9058 633 9059 685
rect 8759 620 9059 633
rect 8759 568 8760 620
rect 8812 568 8842 620
rect 8894 568 8924 620
rect 8976 568 9006 620
rect 9058 568 9059 620
rect 8759 555 9059 568
rect 8759 503 8760 555
rect 8812 503 8842 555
rect 8894 503 8924 555
rect 8976 503 9006 555
rect 9058 503 9059 555
rect 8759 490 9059 503
rect 8759 438 8760 490
rect 8812 438 8842 490
rect 8894 438 8924 490
rect 8976 438 9006 490
rect 9058 438 9059 490
rect 8759 425 9059 438
rect 8759 373 8760 425
rect 8812 373 8842 425
rect 8894 373 8924 425
rect 8976 373 9006 425
rect 9058 373 9059 425
rect 8759 367 9059 373
rect 9583 1902 9883 1908
rect 9583 1850 9584 1902
rect 9636 1850 9666 1902
rect 9718 1850 9748 1902
rect 9800 1850 9830 1902
rect 9882 1850 9883 1902
rect 9583 1838 9883 1850
rect 9583 1786 9584 1838
rect 9636 1786 9666 1838
rect 9718 1786 9748 1838
rect 9800 1786 9830 1838
rect 9882 1786 9883 1838
rect 9583 1774 9883 1786
rect 9583 1722 9584 1774
rect 9636 1722 9666 1774
rect 9718 1722 9748 1774
rect 9800 1722 9830 1774
rect 9882 1722 9883 1774
rect 9583 1710 9883 1722
rect 9583 1658 9584 1710
rect 9636 1658 9666 1710
rect 9718 1658 9748 1710
rect 9800 1658 9830 1710
rect 9882 1658 9883 1710
rect 9583 1646 9883 1658
rect 9583 1594 9584 1646
rect 9636 1594 9666 1646
rect 9718 1594 9748 1646
rect 9800 1594 9830 1646
rect 9882 1594 9883 1646
rect 9583 1582 9883 1594
rect 9583 1530 9584 1582
rect 9636 1530 9666 1582
rect 9718 1530 9748 1582
rect 9800 1530 9830 1582
rect 9882 1530 9883 1582
rect 9583 1518 9883 1530
rect 9583 1466 9584 1518
rect 9636 1466 9666 1518
rect 9718 1466 9748 1518
rect 9800 1466 9830 1518
rect 9882 1466 9883 1518
rect 9583 1454 9883 1466
rect 9583 1402 9584 1454
rect 9636 1402 9666 1454
rect 9718 1402 9748 1454
rect 9800 1402 9830 1454
rect 9882 1402 9883 1454
rect 9583 1390 9883 1402
rect 9583 1338 9584 1390
rect 9636 1338 9666 1390
rect 9718 1338 9748 1390
rect 9800 1338 9830 1390
rect 9882 1338 9883 1390
rect 9583 1326 9883 1338
rect 9583 1274 9584 1326
rect 9636 1274 9666 1326
rect 9718 1274 9748 1326
rect 9800 1274 9830 1326
rect 9882 1274 9883 1326
rect 9583 1262 9883 1274
rect 9583 1210 9584 1262
rect 9636 1210 9666 1262
rect 9718 1210 9748 1262
rect 9800 1210 9830 1262
rect 9882 1210 9883 1262
rect 9583 1198 9883 1210
rect 9583 1146 9584 1198
rect 9636 1146 9666 1198
rect 9718 1146 9748 1198
rect 9800 1146 9830 1198
rect 9882 1146 9883 1198
rect 9583 1134 9883 1146
rect 9583 1082 9584 1134
rect 9636 1082 9666 1134
rect 9718 1082 9748 1134
rect 9800 1082 9830 1134
rect 9882 1082 9883 1134
rect 9583 1070 9883 1082
rect 9583 1018 9584 1070
rect 9636 1018 9666 1070
rect 9718 1018 9748 1070
rect 9800 1018 9830 1070
rect 9882 1018 9883 1070
rect 9583 1006 9883 1018
rect 9583 954 9584 1006
rect 9636 954 9666 1006
rect 9718 954 9748 1006
rect 9800 954 9830 1006
rect 9882 954 9883 1006
rect 9583 942 9883 954
rect 9583 890 9584 942
rect 9636 890 9666 942
rect 9718 890 9748 942
rect 9800 890 9830 942
rect 9882 890 9883 942
rect 9583 878 9883 890
rect 9583 826 9584 878
rect 9636 826 9666 878
rect 9718 826 9748 878
rect 9800 826 9830 878
rect 9882 826 9883 878
rect 9583 814 9883 826
rect 9583 762 9584 814
rect 9636 762 9666 814
rect 9718 762 9748 814
rect 9800 762 9830 814
rect 9882 762 9883 814
rect 9583 750 9883 762
rect 9583 698 9584 750
rect 9636 698 9666 750
rect 9718 698 9748 750
rect 9800 698 9830 750
rect 9882 698 9883 750
rect 9583 685 9883 698
rect 9583 633 9584 685
rect 9636 633 9666 685
rect 9718 633 9748 685
rect 9800 633 9830 685
rect 9882 633 9883 685
rect 9583 620 9883 633
rect 9583 568 9584 620
rect 9636 568 9666 620
rect 9718 568 9748 620
rect 9800 568 9830 620
rect 9882 568 9883 620
rect 9583 555 9883 568
rect 9583 503 9584 555
rect 9636 503 9666 555
rect 9718 503 9748 555
rect 9800 503 9830 555
rect 9882 503 9883 555
rect 9583 490 9883 503
rect 9583 438 9584 490
rect 9636 438 9666 490
rect 9718 438 9748 490
rect 9800 438 9830 490
rect 9882 438 9883 490
rect 9583 425 9883 438
rect 9583 373 9584 425
rect 9636 373 9666 425
rect 9718 373 9748 425
rect 9800 373 9830 425
rect 9882 373 9883 425
rect 9583 367 9883 373
rect 10407 1902 10707 1908
rect 10407 1850 10408 1902
rect 10460 1850 10490 1902
rect 10542 1850 10572 1902
rect 10624 1850 10654 1902
rect 10706 1850 10707 1902
rect 10407 1838 10707 1850
rect 10407 1786 10408 1838
rect 10460 1786 10490 1838
rect 10542 1786 10572 1838
rect 10624 1786 10654 1838
rect 10706 1786 10707 1838
rect 10407 1774 10707 1786
rect 10407 1722 10408 1774
rect 10460 1722 10490 1774
rect 10542 1722 10572 1774
rect 10624 1722 10654 1774
rect 10706 1722 10707 1774
rect 10407 1710 10707 1722
rect 10407 1658 10408 1710
rect 10460 1658 10490 1710
rect 10542 1658 10572 1710
rect 10624 1658 10654 1710
rect 10706 1658 10707 1710
rect 10407 1646 10707 1658
rect 10407 1594 10408 1646
rect 10460 1594 10490 1646
rect 10542 1594 10572 1646
rect 10624 1594 10654 1646
rect 10706 1594 10707 1646
rect 10407 1582 10707 1594
rect 10407 1530 10408 1582
rect 10460 1530 10490 1582
rect 10542 1530 10572 1582
rect 10624 1530 10654 1582
rect 10706 1530 10707 1582
rect 10407 1518 10707 1530
rect 10407 1466 10408 1518
rect 10460 1466 10490 1518
rect 10542 1466 10572 1518
rect 10624 1466 10654 1518
rect 10706 1466 10707 1518
rect 10407 1454 10707 1466
rect 10407 1402 10408 1454
rect 10460 1402 10490 1454
rect 10542 1402 10572 1454
rect 10624 1402 10654 1454
rect 10706 1402 10707 1454
rect 10407 1390 10707 1402
rect 10407 1338 10408 1390
rect 10460 1338 10490 1390
rect 10542 1338 10572 1390
rect 10624 1338 10654 1390
rect 10706 1338 10707 1390
rect 10407 1326 10707 1338
rect 10407 1274 10408 1326
rect 10460 1274 10490 1326
rect 10542 1274 10572 1326
rect 10624 1274 10654 1326
rect 10706 1274 10707 1326
rect 10407 1262 10707 1274
rect 10407 1210 10408 1262
rect 10460 1210 10490 1262
rect 10542 1210 10572 1262
rect 10624 1210 10654 1262
rect 10706 1210 10707 1262
rect 10407 1198 10707 1210
rect 10407 1146 10408 1198
rect 10460 1146 10490 1198
rect 10542 1146 10572 1198
rect 10624 1146 10654 1198
rect 10706 1146 10707 1198
rect 10407 1134 10707 1146
rect 10407 1082 10408 1134
rect 10460 1082 10490 1134
rect 10542 1082 10572 1134
rect 10624 1082 10654 1134
rect 10706 1082 10707 1134
rect 10407 1070 10707 1082
rect 10407 1018 10408 1070
rect 10460 1018 10490 1070
rect 10542 1018 10572 1070
rect 10624 1018 10654 1070
rect 10706 1018 10707 1070
rect 10407 1006 10707 1018
rect 10407 954 10408 1006
rect 10460 954 10490 1006
rect 10542 954 10572 1006
rect 10624 954 10654 1006
rect 10706 954 10707 1006
rect 10407 942 10707 954
rect 10407 890 10408 942
rect 10460 890 10490 942
rect 10542 890 10572 942
rect 10624 890 10654 942
rect 10706 890 10707 942
rect 10407 878 10707 890
rect 10407 826 10408 878
rect 10460 826 10490 878
rect 10542 826 10572 878
rect 10624 826 10654 878
rect 10706 826 10707 878
rect 10407 814 10707 826
rect 10407 762 10408 814
rect 10460 762 10490 814
rect 10542 762 10572 814
rect 10624 762 10654 814
rect 10706 762 10707 814
rect 10407 750 10707 762
rect 10407 698 10408 750
rect 10460 698 10490 750
rect 10542 698 10572 750
rect 10624 698 10654 750
rect 10706 698 10707 750
rect 10407 685 10707 698
rect 10407 633 10408 685
rect 10460 633 10490 685
rect 10542 633 10572 685
rect 10624 633 10654 685
rect 10706 633 10707 685
rect 10407 620 10707 633
rect 10407 568 10408 620
rect 10460 568 10490 620
rect 10542 568 10572 620
rect 10624 568 10654 620
rect 10706 568 10707 620
rect 10407 555 10707 568
rect 10407 503 10408 555
rect 10460 503 10490 555
rect 10542 503 10572 555
rect 10624 503 10654 555
rect 10706 503 10707 555
rect 10407 490 10707 503
rect 10407 438 10408 490
rect 10460 438 10490 490
rect 10542 438 10572 490
rect 10624 438 10654 490
rect 10706 438 10707 490
rect 10407 425 10707 438
rect 10407 373 10408 425
rect 10460 373 10490 425
rect 10542 373 10572 425
rect 10624 373 10654 425
rect 10706 373 10707 425
rect 10407 367 10707 373
rect 12895 374 12975 3936
rect 13064 728 13246 4072
rect 13517 3592 13699 4577
tri 13699 4464 13812 4577 nw
rect 13894 3922 14225 3928
rect 13894 3888 13906 3922
rect 13940 3888 14019 3922
rect 14053 3888 14225 3922
rect 13894 3836 14225 3888
rect 13894 3802 13906 3836
rect 13940 3802 14019 3836
rect 14053 3802 14225 3836
rect 13894 3796 14225 3802
tri 14000 3762 14034 3796 ne
rect 14034 3739 14225 3796
rect 14034 3705 14099 3739
rect 14133 3705 14185 3739
rect 14219 3705 14225 3739
rect 14034 3626 14225 3705
tri 13699 3592 13726 3619 sw
rect 14034 3592 14099 3626
rect 14133 3592 14185 3626
rect 14219 3592 14225 3626
rect 13517 3580 13726 3592
tri 13726 3580 13738 3592 sw
rect 14034 3580 14225 3592
rect 13517 3460 13738 3580
tri 13738 3460 13858 3580 sw
rect 13517 3454 14681 3460
rect 13517 3420 13623 3454
rect 13657 3420 13747 3454
rect 13781 3420 13821 3454
rect 13855 3420 13895 3454
rect 13929 3420 13969 3454
rect 14003 3420 14044 3454
rect 14078 3420 14119 3454
rect 14153 3420 14194 3454
rect 14228 3420 14269 3454
rect 14303 3420 14344 3454
rect 14378 3420 14419 3454
rect 14453 3420 14494 3454
rect 14528 3420 14569 3454
rect 14603 3420 14681 3454
rect 13517 3382 14681 3420
rect 13517 3348 13523 3382
rect 13557 3348 14641 3382
rect 14675 3348 14681 3382
rect 13517 3334 14681 3348
rect 13517 3309 13622 3334
rect 13517 3275 13523 3309
rect 13557 3300 13622 3309
rect 13656 3300 13806 3334
rect 13840 3300 13990 3334
rect 14024 3300 14174 3334
rect 14208 3300 14358 3334
rect 14392 3300 14542 3334
rect 14576 3310 14681 3334
rect 14576 3300 14641 3310
rect 13557 3276 14641 3300
rect 14675 3276 14681 3310
rect 13557 3275 14681 3276
rect 13517 3260 14681 3275
rect 13517 3236 13622 3260
rect 13517 3202 13523 3236
rect 13557 3226 13622 3236
rect 13656 3226 13806 3260
rect 13840 3226 13990 3260
rect 14024 3226 14174 3260
rect 14208 3226 14358 3260
rect 14392 3226 14542 3260
rect 14576 3238 14681 3260
rect 14576 3226 14641 3238
rect 13557 3204 14641 3226
rect 14675 3204 14681 3238
rect 13557 3202 14681 3204
rect 13517 3198 14681 3202
rect 13517 3186 13684 3198
tri 13684 3186 13696 3198 nw
tri 13766 3186 13778 3198 ne
rect 13778 3186 13868 3198
tri 13868 3186 13880 3198 nw
tri 13950 3186 13962 3198 ne
rect 13962 3186 14052 3198
tri 14052 3186 14064 3198 nw
tri 14134 3186 14146 3198 ne
rect 14146 3186 14236 3198
tri 14236 3186 14248 3198 nw
tri 14318 3186 14330 3198 ne
rect 14330 3186 14420 3198
tri 14420 3186 14432 3198 nw
tri 14502 3186 14514 3198 ne
rect 14514 3186 14681 3198
rect 13517 3163 13622 3186
rect 13517 3129 13523 3163
rect 13557 3152 13622 3163
rect 13656 3152 13662 3186
tri 13662 3164 13684 3186 nw
tri 13778 3164 13800 3186 ne
rect 13557 3129 13662 3152
rect 13800 3152 13806 3186
rect 13840 3152 13846 3186
tri 13846 3164 13868 3186 nw
tri 13962 3164 13984 3186 ne
rect 13517 3112 13662 3129
rect 13517 3090 13622 3112
rect 13517 3056 13523 3090
rect 13557 3078 13622 3090
rect 13656 3078 13662 3112
rect 13557 3056 13662 3078
rect 13517 3038 13662 3056
rect 13517 3017 13622 3038
rect 13517 2983 13523 3017
rect 13557 3004 13622 3017
rect 13656 3004 13662 3038
rect 13557 2983 13662 3004
rect 13517 2963 13662 2983
rect 13517 2944 13622 2963
rect 13517 2910 13523 2944
rect 13557 2929 13622 2944
rect 13656 2929 13662 2963
rect 13557 2910 13662 2929
rect 13517 2888 13662 2910
rect 13517 2871 13622 2888
rect 13517 2837 13523 2871
rect 13557 2854 13622 2871
rect 13656 2854 13662 2888
rect 13557 2837 13662 2854
rect 13517 2813 13662 2837
rect 13517 2798 13622 2813
rect 13517 2764 13523 2798
rect 13557 2779 13622 2798
rect 13656 2779 13662 2813
rect 13557 2764 13662 2779
rect 13517 2738 13662 2764
rect 13517 2725 13622 2738
rect 13517 2691 13523 2725
rect 13557 2704 13622 2725
rect 13656 2704 13662 2738
rect 13557 2691 13662 2704
rect 13517 2663 13662 2691
rect 13517 2652 13622 2663
rect 13517 2618 13523 2652
rect 13557 2629 13622 2652
rect 13656 2629 13662 2663
rect 13557 2618 13662 2629
rect 13517 2588 13662 2618
rect 13517 2579 13622 2588
rect 13517 2545 13523 2579
rect 13557 2554 13622 2579
rect 13656 2554 13662 2588
rect 13557 2545 13662 2554
rect 13517 2513 13662 2545
rect 13517 2506 13622 2513
rect 13517 2472 13523 2506
rect 13557 2479 13622 2506
rect 13656 2479 13662 2513
rect 13557 2472 13662 2479
rect 13517 2438 13662 2472
rect 13517 2433 13622 2438
rect 13517 2399 13523 2433
rect 13557 2404 13622 2433
rect 13656 2404 13662 2438
rect 13557 2399 13662 2404
rect 13517 2363 13662 2399
rect 13517 2360 13622 2363
rect 13517 2326 13523 2360
rect 13557 2329 13622 2360
rect 13656 2329 13662 2363
rect 13557 2326 13662 2329
rect 13517 2288 13662 2326
rect 13517 2287 13622 2288
rect 13517 2253 13523 2287
rect 13557 2254 13622 2287
rect 13656 2254 13662 2288
rect 13557 2253 13662 2254
rect 13517 2214 13662 2253
rect 13517 2180 13523 2214
rect 13557 2213 13662 2214
rect 13557 2180 13622 2213
rect 13517 2179 13622 2180
rect 13656 2179 13662 2213
rect 13517 2141 13662 2179
rect 13517 2107 13523 2141
rect 13557 2138 13662 2141
rect 13557 2107 13622 2138
rect 13517 2104 13622 2107
rect 13656 2104 13662 2138
rect 13517 2068 13662 2104
rect 13517 2034 13523 2068
rect 13557 2063 13662 2068
rect 13557 2034 13622 2063
rect 13517 2029 13622 2034
rect 13656 2029 13662 2063
rect 13517 1995 13662 2029
rect 13517 1961 13523 1995
rect 13557 1988 13662 1995
rect 13557 1961 13622 1988
rect 13517 1954 13622 1961
rect 13656 1954 13662 1988
rect 13517 1922 13662 1954
rect 13517 1888 13523 1922
rect 13557 1888 13662 1922
rect 13517 1849 13662 1888
rect 13517 1815 13523 1849
rect 13557 1815 13662 1849
rect 13517 1804 13662 1815
rect 13517 1776 13622 1804
rect 13517 1742 13523 1776
rect 13557 1770 13622 1776
rect 13656 1770 13662 1804
rect 13557 1742 13662 1770
rect 13517 1730 13662 1742
rect 13517 1703 13622 1730
rect 13517 1669 13523 1703
rect 13557 1696 13622 1703
rect 13656 1696 13662 1730
rect 13557 1669 13662 1696
rect 13517 1656 13662 1669
rect 13517 1630 13622 1656
rect 13517 1596 13523 1630
rect 13557 1622 13622 1630
rect 13656 1622 13662 1656
rect 13557 1596 13662 1622
rect 13517 1582 13662 1596
rect 13517 1557 13622 1582
rect 13517 1523 13523 1557
rect 13557 1548 13622 1557
rect 13656 1548 13662 1582
rect 13557 1523 13662 1548
rect 13517 1508 13662 1523
rect 13517 1484 13622 1508
rect 13517 1450 13523 1484
rect 13557 1474 13622 1484
rect 13656 1474 13662 1508
rect 13557 1450 13662 1474
rect 13517 1434 13662 1450
rect 13517 1411 13622 1434
rect 13517 1377 13523 1411
rect 13557 1400 13622 1411
rect 13656 1400 13662 1434
rect 13557 1377 13662 1400
rect 13517 1360 13662 1377
rect 13517 1338 13622 1360
rect 13517 1304 13523 1338
rect 13557 1326 13622 1338
rect 13656 1326 13662 1360
rect 13557 1304 13662 1326
rect 13517 1286 13662 1304
rect 13517 1266 13622 1286
rect 13517 1232 13523 1266
rect 13557 1252 13622 1266
rect 13656 1252 13662 1286
rect 13557 1232 13662 1252
rect 13517 1212 13662 1232
rect 13517 1194 13622 1212
rect 13517 1160 13523 1194
rect 13557 1178 13622 1194
rect 13656 1178 13662 1212
rect 13557 1160 13662 1178
rect 13517 1138 13662 1160
rect 13517 1122 13622 1138
rect 13517 1088 13523 1122
rect 13557 1104 13622 1122
rect 13656 1104 13662 1138
rect 13557 1088 13662 1104
rect 13517 1064 13662 1088
rect 13517 1050 13622 1064
rect 13517 1016 13523 1050
rect 13557 1030 13622 1050
rect 13656 1030 13662 1064
rect 13557 1016 13662 1030
rect 13517 990 13662 1016
rect 13517 978 13622 990
rect 13517 944 13523 978
rect 13557 956 13622 978
rect 13656 956 13662 990
rect 13557 944 13662 956
rect 13517 915 13662 944
rect 13517 906 13622 915
rect 13517 872 13523 906
rect 13557 881 13622 906
rect 13656 881 13662 915
rect 13557 872 13662 881
rect 13517 840 13662 872
rect 13517 834 13622 840
rect 13517 800 13523 834
rect 13557 806 13622 834
rect 13656 806 13662 840
rect 13557 800 13662 806
rect 13517 765 13662 800
rect 13517 762 13622 765
tri 13246 728 13251 733 sw
rect 13517 728 13523 762
rect 13557 731 13622 762
rect 13656 731 13662 765
rect 13557 728 13662 731
rect 13064 724 13251 728
tri 13251 724 13255 728 sw
rect 13064 694 13255 724
tri 13255 694 13285 724 sw
rect 13064 690 13285 694
tri 13285 690 13289 694 sw
rect 13517 690 13662 728
rect 13064 656 13289 690
tri 13289 656 13323 690 sw
rect 13517 656 13523 690
rect 13557 656 13622 690
rect 13656 656 13662 690
rect 13064 649 13323 656
tri 13323 649 13330 656 sw
rect 13064 644 13330 649
tri 13330 644 13335 649 sw
rect 13517 644 13662 656
rect 13708 3132 13754 3144
rect 13708 3098 13714 3132
rect 13748 3098 13754 3132
rect 13708 3057 13754 3098
rect 13708 3023 13714 3057
rect 13748 3023 13754 3057
rect 13708 2982 13754 3023
rect 13708 2948 13714 2982
rect 13748 2948 13754 2982
rect 13708 2907 13754 2948
rect 13708 2873 13714 2907
rect 13748 2873 13754 2907
rect 13708 2832 13754 2873
rect 13708 2798 13714 2832
rect 13748 2798 13754 2832
rect 13708 2757 13754 2798
rect 13708 2723 13714 2757
rect 13748 2723 13754 2757
rect 13708 2682 13754 2723
rect 13708 2648 13714 2682
rect 13748 2648 13754 2682
rect 13708 2606 13754 2648
rect 13708 2572 13714 2606
rect 13748 2572 13754 2606
rect 13708 2530 13754 2572
rect 13708 2496 13714 2530
rect 13748 2496 13754 2530
rect 13708 2454 13754 2496
rect 13708 2420 13714 2454
rect 13748 2420 13754 2454
rect 13708 2378 13754 2420
rect 13708 2344 13714 2378
rect 13748 2344 13754 2378
rect 13708 2302 13754 2344
rect 13708 2268 13714 2302
rect 13748 2268 13754 2302
rect 13708 2226 13754 2268
rect 13708 2192 13714 2226
rect 13748 2192 13754 2226
rect 13708 2150 13754 2192
rect 13708 2116 13714 2150
rect 13748 2116 13754 2150
rect 13708 2074 13754 2116
rect 13708 2040 13714 2074
rect 13748 2040 13754 2074
rect 13708 1804 13754 2040
rect 13708 1770 13714 1804
rect 13748 1770 13754 1804
rect 13708 1730 13754 1770
rect 13708 1696 13714 1730
rect 13748 1696 13754 1730
rect 13708 1656 13754 1696
rect 13708 1622 13714 1656
rect 13748 1622 13754 1656
rect 13708 1582 13754 1622
rect 13708 1548 13714 1582
rect 13748 1548 13754 1582
rect 13708 1508 13754 1548
rect 13708 1474 13714 1508
rect 13748 1474 13754 1508
rect 13708 1434 13754 1474
rect 13708 1400 13714 1434
rect 13748 1400 13754 1434
rect 13708 1360 13754 1400
rect 13708 1326 13714 1360
rect 13748 1326 13754 1360
rect 13708 1286 13754 1326
rect 13708 1252 13714 1286
rect 13748 1252 13754 1286
rect 13708 1212 13754 1252
rect 13708 1178 13714 1212
rect 13748 1178 13754 1212
rect 13708 1138 13754 1178
rect 13708 1104 13714 1138
rect 13748 1104 13754 1138
rect 13708 1064 13754 1104
rect 13708 1030 13714 1064
rect 13748 1030 13754 1064
rect 13708 990 13754 1030
rect 13708 956 13714 990
rect 13748 956 13754 990
rect 13708 916 13754 956
rect 13708 882 13714 916
rect 13748 882 13754 916
rect 13708 842 13754 882
rect 13708 808 13714 842
rect 13748 808 13754 842
rect 13708 768 13754 808
rect 13708 734 13714 768
rect 13748 734 13754 768
rect 13708 694 13754 734
rect 13708 660 13714 694
rect 13748 660 13754 694
rect 13064 642 13335 644
tri 13335 642 13337 644 sw
rect 13064 619 13337 642
tri 13337 619 13360 642 sw
tri 13685 619 13708 642 se
rect 13708 619 13754 660
rect 13800 3112 13846 3152
rect 13984 3152 13990 3186
rect 14024 3152 14030 3186
tri 14030 3164 14052 3186 nw
tri 14146 3164 14168 3186 ne
rect 13800 3078 13806 3112
rect 13840 3078 13846 3112
rect 13800 3038 13846 3078
rect 13800 3004 13806 3038
rect 13840 3004 13846 3038
rect 13800 2963 13846 3004
rect 13800 2929 13806 2963
rect 13840 2929 13846 2963
rect 13800 2888 13846 2929
rect 13800 2854 13806 2888
rect 13840 2854 13846 2888
rect 13800 2813 13846 2854
rect 13800 2779 13806 2813
rect 13840 2779 13846 2813
rect 13800 2738 13846 2779
rect 13800 2704 13806 2738
rect 13840 2704 13846 2738
rect 13800 2663 13846 2704
rect 13800 2629 13806 2663
rect 13840 2629 13846 2663
rect 13800 2588 13846 2629
rect 13800 2554 13806 2588
rect 13840 2554 13846 2588
rect 13800 2513 13846 2554
rect 13800 2479 13806 2513
rect 13840 2479 13846 2513
rect 13800 2438 13846 2479
rect 13800 2404 13806 2438
rect 13840 2404 13846 2438
rect 13800 2363 13846 2404
rect 13800 2329 13806 2363
rect 13840 2329 13846 2363
rect 13800 2288 13846 2329
rect 13800 2254 13806 2288
rect 13840 2254 13846 2288
rect 13800 2213 13846 2254
rect 13800 2179 13806 2213
rect 13840 2179 13846 2213
rect 13800 2138 13846 2179
rect 13800 2104 13806 2138
rect 13840 2104 13846 2138
rect 13800 2063 13846 2104
rect 13800 2029 13806 2063
rect 13840 2029 13846 2063
rect 13800 1988 13846 2029
rect 13800 1954 13806 1988
rect 13840 1954 13846 1988
rect 13800 1804 13846 1954
rect 13800 1770 13806 1804
rect 13840 1770 13846 1804
rect 13800 1730 13846 1770
rect 13800 1696 13806 1730
rect 13840 1696 13846 1730
rect 13800 1656 13846 1696
rect 13800 1622 13806 1656
rect 13840 1622 13846 1656
rect 13800 1582 13846 1622
rect 13800 1548 13806 1582
rect 13840 1548 13846 1582
rect 13800 1508 13846 1548
rect 13800 1474 13806 1508
rect 13840 1474 13846 1508
rect 13800 1434 13846 1474
rect 13800 1400 13806 1434
rect 13840 1400 13846 1434
rect 13800 1360 13846 1400
rect 13800 1326 13806 1360
rect 13840 1326 13846 1360
rect 13800 1286 13846 1326
rect 13800 1252 13806 1286
rect 13840 1252 13846 1286
rect 13800 1212 13846 1252
rect 13800 1178 13806 1212
rect 13840 1178 13846 1212
rect 13800 1138 13846 1178
rect 13800 1104 13806 1138
rect 13840 1104 13846 1138
rect 13800 1064 13846 1104
rect 13800 1030 13806 1064
rect 13840 1030 13846 1064
rect 13800 990 13846 1030
rect 13800 956 13806 990
rect 13840 956 13846 990
rect 13800 915 13846 956
rect 13800 881 13806 915
rect 13840 881 13846 915
rect 13800 840 13846 881
rect 13800 806 13806 840
rect 13840 806 13846 840
rect 13800 765 13846 806
rect 13800 731 13806 765
rect 13840 731 13846 765
rect 13800 690 13846 731
rect 13800 656 13806 690
rect 13840 656 13846 690
rect 13800 644 13846 656
rect 13892 3132 13938 3144
rect 13892 3098 13898 3132
rect 13932 3098 13938 3132
rect 13892 3057 13938 3098
rect 13892 3023 13898 3057
rect 13932 3023 13938 3057
rect 13892 2982 13938 3023
rect 13892 2948 13898 2982
rect 13932 2948 13938 2982
rect 13892 2907 13938 2948
rect 13892 2873 13898 2907
rect 13932 2873 13938 2907
rect 13892 2832 13938 2873
rect 13892 2798 13898 2832
rect 13932 2798 13938 2832
rect 13892 2757 13938 2798
rect 13892 2723 13898 2757
rect 13932 2723 13938 2757
rect 13892 2682 13938 2723
rect 13892 2648 13898 2682
rect 13932 2648 13938 2682
rect 13892 2606 13938 2648
rect 13892 2572 13898 2606
rect 13932 2572 13938 2606
rect 13892 2530 13938 2572
rect 13892 2496 13898 2530
rect 13932 2496 13938 2530
rect 13892 2454 13938 2496
rect 13892 2420 13898 2454
rect 13932 2420 13938 2454
rect 13892 2378 13938 2420
rect 13892 2344 13898 2378
rect 13932 2344 13938 2378
rect 13892 2302 13938 2344
rect 13892 2268 13898 2302
rect 13932 2268 13938 2302
rect 13892 2226 13938 2268
rect 13892 2192 13898 2226
rect 13932 2192 13938 2226
rect 13892 2150 13938 2192
rect 13892 2116 13898 2150
rect 13932 2116 13938 2150
rect 13892 2074 13938 2116
rect 13892 2040 13898 2074
rect 13932 2040 13938 2074
rect 13892 1804 13938 2040
rect 13892 1770 13898 1804
rect 13932 1770 13938 1804
rect 13892 1730 13938 1770
rect 13892 1696 13898 1730
rect 13932 1696 13938 1730
rect 13892 1656 13938 1696
rect 13892 1622 13898 1656
rect 13932 1622 13938 1656
rect 13892 1582 13938 1622
rect 13892 1548 13898 1582
rect 13932 1548 13938 1582
rect 13892 1508 13938 1548
rect 13892 1474 13898 1508
rect 13932 1474 13938 1508
rect 13892 1434 13938 1474
rect 13892 1400 13898 1434
rect 13932 1400 13938 1434
rect 13892 1360 13938 1400
rect 13892 1326 13898 1360
rect 13932 1326 13938 1360
rect 13892 1286 13938 1326
rect 13892 1252 13898 1286
rect 13932 1252 13938 1286
rect 13892 1212 13938 1252
rect 13892 1178 13898 1212
rect 13932 1178 13938 1212
rect 13892 1138 13938 1178
rect 13892 1104 13898 1138
rect 13932 1104 13938 1138
rect 13892 1064 13938 1104
rect 13892 1030 13898 1064
rect 13932 1030 13938 1064
rect 13892 990 13938 1030
rect 13892 956 13898 990
rect 13932 956 13938 990
rect 13892 916 13938 956
rect 13892 882 13898 916
rect 13932 882 13938 916
rect 13892 842 13938 882
rect 13892 808 13898 842
rect 13932 808 13938 842
rect 13892 768 13938 808
rect 13892 734 13898 768
rect 13932 734 13938 768
rect 13892 694 13938 734
rect 13892 660 13898 694
rect 13932 660 13938 694
tri 13754 619 13777 642 sw
tri 13869 619 13892 642 se
rect 13892 619 13938 660
rect 13984 3112 14030 3152
rect 14168 3152 14174 3186
rect 14208 3152 14214 3186
tri 14214 3164 14236 3186 nw
tri 14330 3164 14352 3186 ne
rect 13984 3078 13990 3112
rect 14024 3078 14030 3112
rect 13984 3038 14030 3078
rect 13984 3004 13990 3038
rect 14024 3004 14030 3038
rect 13984 2963 14030 3004
rect 13984 2929 13990 2963
rect 14024 2929 14030 2963
rect 13984 2888 14030 2929
rect 13984 2854 13990 2888
rect 14024 2854 14030 2888
rect 13984 2813 14030 2854
rect 13984 2779 13990 2813
rect 14024 2779 14030 2813
rect 13984 2738 14030 2779
rect 13984 2704 13990 2738
rect 14024 2704 14030 2738
rect 13984 2663 14030 2704
rect 13984 2629 13990 2663
rect 14024 2629 14030 2663
rect 13984 2588 14030 2629
rect 13984 2554 13990 2588
rect 14024 2554 14030 2588
rect 13984 2513 14030 2554
rect 13984 2479 13990 2513
rect 14024 2479 14030 2513
rect 13984 2438 14030 2479
rect 13984 2404 13990 2438
rect 14024 2404 14030 2438
rect 13984 2363 14030 2404
rect 13984 2329 13990 2363
rect 14024 2329 14030 2363
rect 13984 2288 14030 2329
rect 13984 2254 13990 2288
rect 14024 2254 14030 2288
rect 13984 2213 14030 2254
rect 13984 2179 13990 2213
rect 14024 2179 14030 2213
rect 13984 2138 14030 2179
rect 13984 2104 13990 2138
rect 14024 2104 14030 2138
rect 13984 2063 14030 2104
rect 13984 2029 13990 2063
rect 14024 2029 14030 2063
rect 13984 1988 14030 2029
rect 13984 1954 13990 1988
rect 14024 1954 14030 1988
rect 13984 1804 14030 1954
rect 13984 1770 13990 1804
rect 14024 1770 14030 1804
rect 13984 1730 14030 1770
rect 13984 1696 13990 1730
rect 14024 1696 14030 1730
rect 13984 1656 14030 1696
rect 13984 1622 13990 1656
rect 14024 1622 14030 1656
rect 13984 1582 14030 1622
rect 13984 1548 13990 1582
rect 14024 1548 14030 1582
rect 13984 1508 14030 1548
rect 13984 1474 13990 1508
rect 14024 1474 14030 1508
rect 13984 1434 14030 1474
rect 13984 1400 13990 1434
rect 14024 1400 14030 1434
rect 13984 1360 14030 1400
rect 13984 1326 13990 1360
rect 14024 1326 14030 1360
rect 13984 1286 14030 1326
rect 13984 1252 13990 1286
rect 14024 1252 14030 1286
rect 13984 1212 14030 1252
rect 13984 1178 13990 1212
rect 14024 1178 14030 1212
rect 13984 1138 14030 1178
rect 13984 1104 13990 1138
rect 14024 1104 14030 1138
rect 13984 1064 14030 1104
rect 13984 1030 13990 1064
rect 14024 1030 14030 1064
rect 13984 990 14030 1030
rect 13984 956 13990 990
rect 14024 956 14030 990
rect 13984 915 14030 956
rect 13984 881 13990 915
rect 14024 881 14030 915
rect 13984 840 14030 881
rect 13984 806 13990 840
rect 14024 806 14030 840
rect 13984 765 14030 806
rect 13984 731 13990 765
rect 14024 731 14030 765
rect 13984 690 14030 731
rect 13984 656 13990 690
rect 14024 656 14030 690
rect 13984 644 14030 656
rect 14076 3132 14122 3144
rect 14076 3098 14082 3132
rect 14116 3098 14122 3132
rect 14076 3057 14122 3098
rect 14076 3023 14082 3057
rect 14116 3023 14122 3057
rect 14076 2982 14122 3023
rect 14076 2948 14082 2982
rect 14116 2948 14122 2982
rect 14076 2907 14122 2948
rect 14076 2873 14082 2907
rect 14116 2873 14122 2907
rect 14076 2832 14122 2873
rect 14076 2798 14082 2832
rect 14116 2798 14122 2832
rect 14076 2757 14122 2798
rect 14076 2723 14082 2757
rect 14116 2723 14122 2757
rect 14076 2682 14122 2723
rect 14076 2648 14082 2682
rect 14116 2648 14122 2682
rect 14076 2606 14122 2648
rect 14076 2572 14082 2606
rect 14116 2572 14122 2606
rect 14076 2530 14122 2572
rect 14076 2496 14082 2530
rect 14116 2496 14122 2530
rect 14076 2454 14122 2496
rect 14076 2420 14082 2454
rect 14116 2420 14122 2454
rect 14076 2378 14122 2420
rect 14076 2344 14082 2378
rect 14116 2344 14122 2378
rect 14076 2302 14122 2344
rect 14076 2268 14082 2302
rect 14116 2268 14122 2302
rect 14076 2226 14122 2268
rect 14076 2192 14082 2226
rect 14116 2192 14122 2226
rect 14076 2150 14122 2192
rect 14076 2116 14082 2150
rect 14116 2116 14122 2150
rect 14076 2074 14122 2116
rect 14076 2040 14082 2074
rect 14116 2040 14122 2074
rect 14076 1804 14122 2040
rect 14076 1770 14082 1804
rect 14116 1770 14122 1804
rect 14076 1730 14122 1770
rect 14076 1696 14082 1730
rect 14116 1696 14122 1730
rect 14076 1656 14122 1696
rect 14076 1622 14082 1656
rect 14116 1622 14122 1656
rect 14076 1582 14122 1622
rect 14076 1548 14082 1582
rect 14116 1548 14122 1582
rect 14076 1508 14122 1548
rect 14076 1474 14082 1508
rect 14116 1474 14122 1508
rect 14076 1434 14122 1474
rect 14076 1400 14082 1434
rect 14116 1400 14122 1434
rect 14076 1360 14122 1400
rect 14076 1326 14082 1360
rect 14116 1326 14122 1360
rect 14076 1286 14122 1326
rect 14076 1252 14082 1286
rect 14116 1252 14122 1286
rect 14076 1212 14122 1252
rect 14076 1178 14082 1212
rect 14116 1178 14122 1212
rect 14076 1138 14122 1178
rect 14076 1104 14082 1138
rect 14116 1104 14122 1138
rect 14076 1064 14122 1104
rect 14076 1030 14082 1064
rect 14116 1030 14122 1064
rect 14076 990 14122 1030
rect 14076 956 14082 990
rect 14116 956 14122 990
rect 14076 916 14122 956
rect 14076 882 14082 916
rect 14116 882 14122 916
rect 14076 842 14122 882
rect 14076 808 14082 842
rect 14116 808 14122 842
rect 14076 768 14122 808
rect 14076 734 14082 768
rect 14116 734 14122 768
rect 14076 694 14122 734
rect 14076 660 14082 694
rect 14116 660 14122 694
tri 13938 619 13961 642 sw
tri 14053 619 14076 642 se
rect 14076 619 14122 660
rect 14168 3112 14214 3152
rect 14352 3152 14358 3186
rect 14392 3152 14398 3186
tri 14398 3164 14420 3186 nw
tri 14514 3164 14536 3186 ne
rect 14168 3078 14174 3112
rect 14208 3078 14214 3112
rect 14168 3038 14214 3078
rect 14168 3004 14174 3038
rect 14208 3004 14214 3038
rect 14168 2963 14214 3004
rect 14168 2929 14174 2963
rect 14208 2929 14214 2963
rect 14168 2888 14214 2929
rect 14168 2854 14174 2888
rect 14208 2854 14214 2888
rect 14168 2813 14214 2854
rect 14168 2779 14174 2813
rect 14208 2779 14214 2813
rect 14168 2738 14214 2779
rect 14168 2704 14174 2738
rect 14208 2704 14214 2738
rect 14168 2663 14214 2704
rect 14168 2629 14174 2663
rect 14208 2629 14214 2663
rect 14168 2588 14214 2629
rect 14168 2554 14174 2588
rect 14208 2554 14214 2588
rect 14168 2513 14214 2554
rect 14168 2479 14174 2513
rect 14208 2479 14214 2513
rect 14168 2438 14214 2479
rect 14168 2404 14174 2438
rect 14208 2404 14214 2438
rect 14168 2363 14214 2404
rect 14168 2329 14174 2363
rect 14208 2329 14214 2363
rect 14168 2288 14214 2329
rect 14168 2254 14174 2288
rect 14208 2254 14214 2288
rect 14168 2213 14214 2254
rect 14168 2179 14174 2213
rect 14208 2179 14214 2213
rect 14168 2138 14214 2179
rect 14168 2104 14174 2138
rect 14208 2104 14214 2138
rect 14168 2063 14214 2104
rect 14168 2029 14174 2063
rect 14208 2029 14214 2063
rect 14168 1988 14214 2029
rect 14168 1954 14174 1988
rect 14208 1954 14214 1988
rect 14168 1804 14214 1954
rect 14168 1770 14174 1804
rect 14208 1770 14214 1804
rect 14168 1730 14214 1770
rect 14168 1696 14174 1730
rect 14208 1696 14214 1730
rect 14168 1656 14214 1696
rect 14168 1622 14174 1656
rect 14208 1622 14214 1656
rect 14168 1582 14214 1622
rect 14168 1548 14174 1582
rect 14208 1548 14214 1582
rect 14168 1508 14214 1548
rect 14168 1474 14174 1508
rect 14208 1474 14214 1508
rect 14168 1434 14214 1474
rect 14168 1400 14174 1434
rect 14208 1400 14214 1434
rect 14168 1360 14214 1400
rect 14168 1326 14174 1360
rect 14208 1326 14214 1360
rect 14168 1286 14214 1326
rect 14168 1252 14174 1286
rect 14208 1252 14214 1286
rect 14168 1212 14214 1252
rect 14168 1178 14174 1212
rect 14208 1178 14214 1212
rect 14168 1138 14214 1178
rect 14168 1104 14174 1138
rect 14208 1104 14214 1138
rect 14168 1064 14214 1104
rect 14168 1030 14174 1064
rect 14208 1030 14214 1064
rect 14168 990 14214 1030
rect 14168 956 14174 990
rect 14208 956 14214 990
rect 14168 915 14214 956
rect 14168 881 14174 915
rect 14208 881 14214 915
rect 14168 840 14214 881
rect 14168 806 14174 840
rect 14208 806 14214 840
rect 14168 765 14214 806
rect 14168 731 14174 765
rect 14208 731 14214 765
rect 14168 690 14214 731
rect 14168 656 14174 690
rect 14208 656 14214 690
rect 14168 644 14214 656
rect 14260 3132 14306 3144
rect 14260 3098 14266 3132
rect 14300 3098 14306 3132
rect 14260 3057 14306 3098
rect 14260 3023 14266 3057
rect 14300 3023 14306 3057
rect 14260 2982 14306 3023
rect 14260 2948 14266 2982
rect 14300 2948 14306 2982
rect 14260 2907 14306 2948
rect 14260 2873 14266 2907
rect 14300 2873 14306 2907
rect 14260 2832 14306 2873
rect 14260 2798 14266 2832
rect 14300 2798 14306 2832
rect 14260 2757 14306 2798
rect 14260 2723 14266 2757
rect 14300 2723 14306 2757
rect 14260 2682 14306 2723
rect 14260 2648 14266 2682
rect 14300 2648 14306 2682
rect 14260 2606 14306 2648
rect 14260 2572 14266 2606
rect 14300 2572 14306 2606
rect 14260 2530 14306 2572
rect 14260 2496 14266 2530
rect 14300 2496 14306 2530
rect 14260 2454 14306 2496
rect 14260 2420 14266 2454
rect 14300 2420 14306 2454
rect 14260 2378 14306 2420
rect 14260 2344 14266 2378
rect 14300 2344 14306 2378
rect 14260 2302 14306 2344
rect 14260 2268 14266 2302
rect 14300 2268 14306 2302
rect 14260 2226 14306 2268
rect 14260 2192 14266 2226
rect 14300 2192 14306 2226
rect 14260 2150 14306 2192
rect 14260 2116 14266 2150
rect 14300 2116 14306 2150
rect 14260 2074 14306 2116
rect 14260 2040 14266 2074
rect 14300 2040 14306 2074
rect 14260 1804 14306 2040
rect 14260 1770 14266 1804
rect 14300 1770 14306 1804
rect 14260 1730 14306 1770
rect 14260 1696 14266 1730
rect 14300 1696 14306 1730
rect 14260 1656 14306 1696
rect 14260 1622 14266 1656
rect 14300 1622 14306 1656
rect 14260 1582 14306 1622
rect 14260 1548 14266 1582
rect 14300 1548 14306 1582
rect 14260 1508 14306 1548
rect 14260 1474 14266 1508
rect 14300 1474 14306 1508
rect 14260 1434 14306 1474
rect 14260 1400 14266 1434
rect 14300 1400 14306 1434
rect 14260 1360 14306 1400
rect 14260 1326 14266 1360
rect 14300 1326 14306 1360
rect 14260 1286 14306 1326
rect 14260 1252 14266 1286
rect 14300 1252 14306 1286
rect 14260 1212 14306 1252
rect 14260 1178 14266 1212
rect 14300 1178 14306 1212
rect 14260 1138 14306 1178
rect 14260 1104 14266 1138
rect 14300 1104 14306 1138
rect 14260 1064 14306 1104
rect 14260 1030 14266 1064
rect 14300 1030 14306 1064
rect 14260 990 14306 1030
rect 14260 956 14266 990
rect 14300 956 14306 990
rect 14260 916 14306 956
rect 14260 882 14266 916
rect 14300 882 14306 916
rect 14260 842 14306 882
rect 14260 808 14266 842
rect 14300 808 14306 842
rect 14260 768 14306 808
rect 14260 734 14266 768
rect 14300 734 14306 768
rect 14260 694 14306 734
rect 14260 660 14266 694
rect 14300 660 14306 694
tri 14122 619 14145 642 sw
tri 14237 619 14260 642 se
rect 14260 619 14306 660
rect 14352 3112 14398 3152
rect 14536 3152 14542 3186
rect 14576 3166 14681 3186
rect 14576 3152 14641 3166
rect 14352 3078 14358 3112
rect 14392 3078 14398 3112
rect 14352 3038 14398 3078
rect 14352 3004 14358 3038
rect 14392 3004 14398 3038
rect 14352 2963 14398 3004
rect 14352 2929 14358 2963
rect 14392 2929 14398 2963
rect 14352 2888 14398 2929
rect 14352 2854 14358 2888
rect 14392 2854 14398 2888
rect 14352 2813 14398 2854
rect 14352 2779 14358 2813
rect 14392 2779 14398 2813
rect 14352 2738 14398 2779
rect 14352 2704 14358 2738
rect 14392 2704 14398 2738
rect 14352 2663 14398 2704
rect 14352 2629 14358 2663
rect 14392 2629 14398 2663
rect 14352 2588 14398 2629
rect 14352 2554 14358 2588
rect 14392 2554 14398 2588
rect 14352 2513 14398 2554
rect 14352 2479 14358 2513
rect 14392 2479 14398 2513
rect 14352 2438 14398 2479
rect 14352 2404 14358 2438
rect 14392 2404 14398 2438
rect 14352 2363 14398 2404
rect 14352 2329 14358 2363
rect 14392 2329 14398 2363
rect 14352 2288 14398 2329
rect 14352 2254 14358 2288
rect 14392 2254 14398 2288
rect 14352 2213 14398 2254
rect 14352 2179 14358 2213
rect 14392 2179 14398 2213
rect 14352 2138 14398 2179
rect 14352 2104 14358 2138
rect 14392 2104 14398 2138
rect 14352 2063 14398 2104
rect 14352 2029 14358 2063
rect 14392 2029 14398 2063
rect 14352 1988 14398 2029
rect 14352 1954 14358 1988
rect 14392 1954 14398 1988
rect 14352 1804 14398 1954
rect 14352 1770 14358 1804
rect 14392 1770 14398 1804
rect 14352 1730 14398 1770
rect 14352 1696 14358 1730
rect 14392 1696 14398 1730
rect 14352 1656 14398 1696
rect 14352 1622 14358 1656
rect 14392 1622 14398 1656
rect 14352 1582 14398 1622
rect 14352 1548 14358 1582
rect 14392 1548 14398 1582
rect 14352 1508 14398 1548
rect 14352 1474 14358 1508
rect 14392 1474 14398 1508
rect 14352 1434 14398 1474
rect 14352 1400 14358 1434
rect 14392 1400 14398 1434
rect 14352 1360 14398 1400
rect 14352 1326 14358 1360
rect 14392 1326 14398 1360
rect 14352 1286 14398 1326
rect 14352 1252 14358 1286
rect 14392 1252 14398 1286
rect 14352 1212 14398 1252
rect 14352 1178 14358 1212
rect 14392 1178 14398 1212
rect 14352 1138 14398 1178
rect 14352 1104 14358 1138
rect 14392 1104 14398 1138
rect 14352 1064 14398 1104
rect 14352 1030 14358 1064
rect 14392 1030 14398 1064
rect 14352 990 14398 1030
rect 14352 956 14358 990
rect 14392 956 14398 990
rect 14352 915 14398 956
rect 14352 881 14358 915
rect 14392 881 14398 915
rect 14352 840 14398 881
rect 14352 806 14358 840
rect 14392 806 14398 840
rect 14352 765 14398 806
rect 14352 731 14358 765
rect 14392 731 14398 765
rect 14352 690 14398 731
rect 14352 656 14358 690
rect 14392 656 14398 690
rect 14352 644 14398 656
rect 14444 3132 14490 3144
rect 14444 3098 14450 3132
rect 14484 3098 14490 3132
rect 14444 3057 14490 3098
rect 14444 3023 14450 3057
rect 14484 3023 14490 3057
rect 14444 2982 14490 3023
rect 14444 2948 14450 2982
rect 14484 2948 14490 2982
rect 14444 2907 14490 2948
rect 14444 2873 14450 2907
rect 14484 2873 14490 2907
rect 14444 2832 14490 2873
rect 14444 2798 14450 2832
rect 14484 2798 14490 2832
rect 14444 2757 14490 2798
rect 14444 2723 14450 2757
rect 14484 2723 14490 2757
rect 14444 2682 14490 2723
rect 14444 2648 14450 2682
rect 14484 2648 14490 2682
rect 14444 2606 14490 2648
rect 14444 2572 14450 2606
rect 14484 2572 14490 2606
rect 14444 2530 14490 2572
rect 14444 2496 14450 2530
rect 14484 2496 14490 2530
rect 14444 2454 14490 2496
rect 14444 2420 14450 2454
rect 14484 2420 14490 2454
rect 14444 2378 14490 2420
rect 14444 2344 14450 2378
rect 14484 2344 14490 2378
rect 14444 2302 14490 2344
rect 14444 2268 14450 2302
rect 14484 2268 14490 2302
rect 14444 2226 14490 2268
rect 14444 2192 14450 2226
rect 14484 2192 14490 2226
rect 14444 2150 14490 2192
rect 14444 2116 14450 2150
rect 14484 2116 14490 2150
rect 14444 2074 14490 2116
rect 14444 2040 14450 2074
rect 14484 2040 14490 2074
rect 14444 1804 14490 2040
rect 14444 1770 14450 1804
rect 14484 1770 14490 1804
rect 14444 1730 14490 1770
rect 14444 1696 14450 1730
rect 14484 1696 14490 1730
rect 14444 1656 14490 1696
rect 14444 1622 14450 1656
rect 14484 1622 14490 1656
rect 14444 1582 14490 1622
rect 14444 1548 14450 1582
rect 14484 1548 14490 1582
rect 14444 1508 14490 1548
rect 14444 1474 14450 1508
rect 14484 1474 14490 1508
rect 14444 1434 14490 1474
rect 14444 1400 14450 1434
rect 14484 1400 14490 1434
rect 14444 1360 14490 1400
rect 14444 1326 14450 1360
rect 14484 1326 14490 1360
rect 14444 1286 14490 1326
rect 14444 1252 14450 1286
rect 14484 1252 14490 1286
rect 14444 1212 14490 1252
rect 14444 1178 14450 1212
rect 14484 1178 14490 1212
rect 14444 1138 14490 1178
rect 14444 1104 14450 1138
rect 14484 1104 14490 1138
rect 14444 1064 14490 1104
rect 14444 1030 14450 1064
rect 14484 1030 14490 1064
rect 14444 990 14490 1030
rect 14444 956 14450 990
rect 14484 956 14490 990
rect 14444 916 14490 956
rect 14444 882 14450 916
rect 14484 882 14490 916
rect 14444 842 14490 882
rect 14444 808 14450 842
rect 14484 808 14490 842
rect 14444 768 14490 808
rect 14444 734 14450 768
rect 14484 734 14490 768
rect 14444 694 14490 734
rect 14444 660 14450 694
rect 14484 660 14490 694
tri 14306 619 14329 642 sw
tri 14421 619 14444 642 se
rect 14444 619 14490 660
rect 13064 608 13360 619
tri 13360 608 13371 619 sw
tri 13674 608 13685 619 se
rect 13685 608 13714 619
rect 13064 585 13714 608
rect 13748 608 13777 619
tri 13777 608 13788 619 sw
tri 13858 608 13869 619 se
rect 13869 608 13898 619
rect 13748 585 13898 608
rect 13932 608 13961 619
tri 13961 608 13972 619 sw
tri 14042 608 14053 619 se
rect 14053 608 14082 619
rect 13932 585 14082 608
rect 14116 608 14145 619
tri 14145 608 14156 619 sw
tri 14226 608 14237 619 se
rect 14237 608 14266 619
rect 14116 585 14266 608
rect 14300 608 14329 619
tri 14329 608 14340 619 sw
tri 14410 608 14421 619 se
rect 14421 608 14450 619
rect 14300 585 14450 608
rect 14484 585 14490 619
rect 13064 544 14490 585
rect 13064 537 13714 544
tri 13064 510 13091 537 ne
rect 13091 510 13714 537
rect 13748 510 13898 544
rect 13932 510 14082 544
rect 14116 510 14266 544
rect 14300 510 14450 544
rect 14484 510 14490 544
tri 13091 499 13102 510 ne
rect 13102 499 14490 510
tri 13102 468 13133 499 ne
rect 13133 468 14490 499
tri 13133 458 13143 468 ne
rect 13143 458 14490 468
tri 13143 424 13177 458 ne
rect 13177 424 14490 458
tri 13177 408 13193 424 ne
rect 13193 408 14490 424
rect 14536 3132 14641 3152
rect 14675 3132 14681 3166
rect 14536 3112 14681 3132
rect 14536 3078 14542 3112
rect 14576 3094 14681 3112
rect 14576 3078 14641 3094
rect 14536 3060 14641 3078
rect 14675 3060 14681 3094
rect 14536 3038 14681 3060
rect 14536 3004 14542 3038
rect 14576 3022 14681 3038
rect 14576 3004 14641 3022
rect 14536 2988 14641 3004
rect 14675 2988 14681 3022
rect 14536 2963 14681 2988
rect 14536 2929 14542 2963
rect 14576 2950 14681 2963
rect 14576 2929 14641 2950
rect 14536 2916 14641 2929
rect 14675 2916 14681 2950
rect 14536 2888 14681 2916
rect 14536 2854 14542 2888
rect 14576 2877 14681 2888
rect 14576 2854 14641 2877
rect 14536 2843 14641 2854
rect 14675 2843 14681 2877
rect 14536 2813 14681 2843
rect 14536 2779 14542 2813
rect 14576 2804 14681 2813
rect 14576 2779 14641 2804
rect 14536 2770 14641 2779
rect 14675 2770 14681 2804
rect 14536 2738 14681 2770
rect 14536 2704 14542 2738
rect 14576 2731 14681 2738
rect 14576 2704 14641 2731
rect 14536 2697 14641 2704
rect 14675 2697 14681 2731
rect 14536 2663 14681 2697
rect 14536 2629 14542 2663
rect 14576 2658 14681 2663
rect 14576 2629 14641 2658
rect 14536 2624 14641 2629
rect 14675 2624 14681 2658
rect 14536 2588 14681 2624
rect 14536 2554 14542 2588
rect 14576 2585 14681 2588
rect 14576 2554 14641 2585
rect 14536 2551 14641 2554
rect 14675 2551 14681 2585
rect 14536 2513 14681 2551
rect 14536 2479 14542 2513
rect 14576 2512 14681 2513
rect 14576 2479 14641 2512
rect 14536 2478 14641 2479
rect 14675 2478 14681 2512
rect 14536 2439 14681 2478
rect 14536 2438 14641 2439
rect 14536 2404 14542 2438
rect 14576 2405 14641 2438
rect 14675 2405 14681 2439
rect 14576 2404 14681 2405
rect 14536 2366 14681 2404
rect 14536 2363 14641 2366
rect 14536 2329 14542 2363
rect 14576 2332 14641 2363
rect 14675 2332 14681 2366
rect 14576 2329 14681 2332
rect 14536 2293 14681 2329
rect 14536 2288 14641 2293
rect 14536 2254 14542 2288
rect 14576 2259 14641 2288
rect 14675 2259 14681 2293
rect 14576 2254 14681 2259
rect 14536 2220 14681 2254
rect 14536 2213 14641 2220
rect 14536 2179 14542 2213
rect 14576 2186 14641 2213
rect 14675 2186 14681 2220
rect 14576 2179 14681 2186
rect 14536 2147 14681 2179
rect 14536 2138 14641 2147
rect 14536 2104 14542 2138
rect 14576 2113 14641 2138
rect 14675 2113 14681 2147
rect 14576 2104 14681 2113
rect 14536 2074 14681 2104
rect 14536 2063 14641 2074
rect 14536 2029 14542 2063
rect 14576 2040 14641 2063
rect 14675 2040 14681 2074
rect 14576 2029 14681 2040
rect 14536 2001 14681 2029
rect 14536 1988 14641 2001
rect 14536 1954 14542 1988
rect 14576 1967 14641 1988
rect 14675 1967 14681 2001
rect 14576 1954 14681 1967
rect 14536 1928 14681 1954
rect 14536 1894 14641 1928
rect 14675 1894 14681 1928
rect 14536 1855 14681 1894
rect 14536 1821 14641 1855
rect 14675 1821 14681 1855
rect 14536 1804 14681 1821
rect 14536 1770 14542 1804
rect 14576 1782 14681 1804
rect 14576 1770 14641 1782
rect 14536 1748 14641 1770
rect 14675 1748 14681 1782
rect 14536 1730 14681 1748
rect 14536 1696 14542 1730
rect 14576 1709 14681 1730
rect 14576 1696 14641 1709
rect 14536 1675 14641 1696
rect 14675 1675 14681 1709
rect 14536 1656 14681 1675
rect 14536 1622 14542 1656
rect 14576 1636 14681 1656
rect 14576 1622 14641 1636
rect 14536 1602 14641 1622
rect 14675 1602 14681 1636
rect 14536 1582 14681 1602
rect 14536 1548 14542 1582
rect 14576 1563 14681 1582
rect 14576 1548 14641 1563
rect 14536 1529 14641 1548
rect 14675 1529 14681 1563
rect 14536 1508 14681 1529
rect 14536 1474 14542 1508
rect 14576 1490 14681 1508
rect 14576 1474 14641 1490
rect 14536 1456 14641 1474
rect 14675 1456 14681 1490
rect 14536 1433 14681 1456
rect 14536 1399 14542 1433
rect 14576 1417 14681 1433
rect 14576 1399 14641 1417
rect 14536 1383 14641 1399
rect 14675 1383 14681 1417
rect 14536 1358 14681 1383
rect 14536 1324 14542 1358
rect 14576 1344 14681 1358
rect 14576 1324 14641 1344
rect 14536 1310 14641 1324
rect 14675 1310 14681 1344
rect 14536 1283 14681 1310
rect 14536 1249 14542 1283
rect 14576 1271 14681 1283
rect 14576 1249 14641 1271
rect 14536 1237 14641 1249
rect 14675 1237 14681 1271
rect 14536 1208 14681 1237
rect 14536 1174 14542 1208
rect 14576 1198 14681 1208
rect 14576 1174 14641 1198
rect 14536 1164 14641 1174
rect 14675 1164 14681 1198
rect 14536 1133 14681 1164
rect 14536 1099 14542 1133
rect 14576 1125 14681 1133
rect 14576 1099 14641 1125
rect 14536 1091 14641 1099
rect 14675 1091 14681 1125
rect 14536 1058 14681 1091
rect 14536 1024 14542 1058
rect 14576 1052 14681 1058
rect 14576 1024 14641 1052
rect 14536 1018 14641 1024
rect 14675 1018 14681 1052
rect 14536 983 14681 1018
rect 14536 949 14542 983
rect 14576 979 14681 983
rect 14576 949 14641 979
rect 14536 945 14641 949
rect 14675 945 14681 979
rect 14536 908 14681 945
rect 14536 874 14542 908
rect 14576 906 14681 908
rect 14576 874 14641 906
rect 14536 872 14641 874
rect 14675 872 14681 906
rect 14536 833 14681 872
rect 14536 799 14542 833
rect 14576 799 14641 833
rect 14675 799 14681 833
rect 14536 760 14681 799
rect 14536 758 14641 760
rect 14536 724 14542 758
rect 14576 726 14641 758
rect 14675 726 14681 760
rect 14576 724 14681 726
rect 14536 687 14681 724
rect 14536 683 14641 687
rect 14536 649 14542 683
rect 14576 653 14641 683
rect 14675 653 14681 687
rect 14576 649 14681 653
rect 14536 614 14681 649
rect 14536 608 14641 614
rect 14536 574 14542 608
rect 14576 580 14641 608
rect 14675 580 14681 614
rect 14576 574 14681 580
rect 14536 541 14681 574
rect 14536 533 14641 541
rect 14536 499 14542 533
rect 14576 507 14641 533
rect 14675 507 14681 541
rect 14576 499 14681 507
rect 14536 468 14681 499
rect 14536 458 14641 468
rect 14536 424 14542 458
rect 14576 434 14641 458
rect 14675 434 14681 468
rect 14576 424 14681 434
rect 14536 412 14681 424
tri 14536 408 14540 412 ne
rect 14540 408 14681 412
tri 14540 395 14553 408 ne
rect 14553 395 14681 408
tri 14553 387 14561 395 ne
rect 14561 387 14641 395
tri 12975 374 12988 387 sw
tri 14561 384 14564 387 ne
rect 12895 368 12988 374
tri 12988 368 12994 374 sw
tri 13661 368 13667 374 se
rect 13667 368 14531 374
rect 1671 322 3276 360
rect 1671 288 1750 322
rect 1784 288 1823 322
rect 1857 288 1896 322
rect 1930 288 1969 322
rect 2003 288 2042 322
rect 2076 288 2115 322
rect 2149 288 2188 322
rect 2222 288 2261 322
rect 2295 288 2334 322
rect 2368 288 2407 322
rect 2441 288 2480 322
rect 2514 288 2553 322
rect 2587 288 2626 322
rect 2660 288 2699 322
rect 2733 288 2772 322
rect 2806 288 2845 322
rect 2879 288 2918 322
rect 2952 288 2991 322
rect 3025 288 3064 322
rect 3098 288 3137 322
rect 3171 288 3210 322
rect 3244 288 3276 322
rect 1671 282 3276 288
rect 3331 357 11313 364
rect 3331 356 5149 357
rect 3331 304 4191 356
rect 4243 304 4259 356
rect 4311 304 4327 356
rect 4379 304 4395 356
rect 4447 304 4463 356
rect 4515 304 4531 356
rect 4583 304 4599 356
rect 4651 304 4666 356
rect 4718 304 4733 356
rect 4785 304 4800 356
rect 4852 304 4867 356
rect 4919 304 4934 356
rect 4986 304 5001 356
rect 5053 304 5068 356
rect 5120 305 5149 356
rect 5201 305 5221 357
rect 5273 305 5293 357
rect 5345 305 5365 357
rect 5417 305 5436 357
rect 5488 305 5507 357
rect 5559 305 5578 357
rect 5630 356 11313 357
rect 5630 305 5659 356
rect 5120 304 5659 305
rect 5711 304 5724 356
rect 5776 304 5789 356
rect 5841 304 5854 356
rect 5906 304 5919 356
rect 5971 304 5984 356
rect 6036 304 6049 356
rect 6101 304 6114 356
rect 6166 304 6179 356
rect 6231 304 6244 356
rect 6296 304 6309 356
rect 6361 304 6374 356
rect 6426 304 6439 356
rect 6491 304 6504 356
rect 6556 304 6569 356
rect 6621 304 6634 356
rect 6686 304 6699 356
rect 6751 304 6764 356
rect 6816 304 6829 356
rect 6881 304 6894 356
rect 6946 304 6959 356
rect 7011 304 7024 356
rect 7076 304 7089 356
rect 7141 304 7154 356
rect 7206 304 7219 356
rect 7271 304 7284 356
rect 7336 304 7349 356
rect 7401 304 7414 356
rect 7466 304 7479 356
rect 7531 304 7544 356
rect 7596 304 7609 356
rect 7661 304 7674 356
rect 7726 304 7739 356
rect 7791 304 7804 356
rect 7856 304 7869 356
rect 7921 304 7934 356
rect 7986 304 7999 356
rect 8051 304 8064 356
rect 8116 304 8129 356
rect 8181 304 8194 356
rect 8246 304 8259 356
rect 8311 304 8324 356
rect 8376 304 8389 356
rect 8441 304 8454 356
rect 8506 304 8519 356
rect 8571 304 8584 356
rect 8636 304 8649 356
rect 8701 304 8714 356
rect 8766 304 8779 356
rect 8831 304 8844 356
rect 8896 304 8909 356
rect 8961 304 8974 356
rect 9026 304 9039 356
rect 9091 304 9104 356
rect 9156 304 9169 356
rect 9221 304 9234 356
rect 9286 304 9299 356
rect 9351 304 9364 356
rect 9416 304 9429 356
rect 9481 304 9494 356
rect 9546 304 9559 356
rect 9611 304 9624 356
rect 9676 304 9689 356
rect 9741 304 9753 356
rect 9805 304 9817 356
rect 9869 304 9881 356
rect 9933 304 9945 356
rect 9997 304 10009 356
rect 10061 304 10073 356
rect 10125 304 10137 356
rect 10189 304 10201 356
rect 10253 304 10265 356
rect 10317 304 10329 356
rect 10381 304 10393 356
rect 10445 304 10457 356
rect 10509 304 10521 356
rect 10573 304 10585 356
rect 10637 304 10649 356
rect 10701 304 11313 356
rect 12895 353 12994 368
tri 12994 353 13009 368 sw
tri 13646 353 13661 368 se
rect 13661 353 13679 368
rect 12895 347 13679 353
rect 12895 307 13340 347
rect 3331 282 11313 304
rect 3331 230 4191 282
rect 4243 230 4259 282
rect 4311 230 4327 282
rect 4379 230 4395 282
rect 4447 230 4463 282
rect 4515 230 4531 282
rect 4583 230 4599 282
rect 4651 230 4666 282
rect 4718 230 4733 282
rect 4785 230 4800 282
rect 4852 230 4867 282
rect 4919 230 4934 282
rect 4986 230 5001 282
rect 5053 230 5068 282
rect 5120 277 5659 282
rect 5120 230 5149 277
rect 3331 225 5149 230
rect 5201 225 5221 277
rect 5273 225 5293 277
rect 5345 225 5365 277
rect 5417 225 5436 277
rect 5488 225 5507 277
rect 5559 225 5578 277
rect 5630 230 5659 277
rect 5711 230 5724 282
rect 5776 230 5789 282
rect 5841 230 5854 282
rect 5906 230 5919 282
rect 5971 230 5984 282
rect 6036 230 6049 282
rect 6101 230 6114 282
rect 6166 230 6179 282
rect 6231 230 6244 282
rect 6296 230 6309 282
rect 6361 230 6374 282
rect 6426 230 6439 282
rect 6491 230 6504 282
rect 6556 230 6569 282
rect 6621 230 6634 282
rect 6686 230 6699 282
rect 6751 230 6764 282
rect 6816 230 6829 282
rect 6881 230 6894 282
rect 6946 230 6959 282
rect 7011 230 7024 282
rect 7076 230 7089 282
rect 7141 230 7154 282
rect 7206 230 7219 282
rect 7271 230 7284 282
rect 7336 230 7349 282
rect 7401 230 7414 282
rect 7466 230 7479 282
rect 7531 230 7544 282
rect 7596 230 7609 282
rect 7661 230 7674 282
rect 7726 230 7739 282
rect 7791 230 7804 282
rect 7856 230 7869 282
rect 7921 230 7934 282
rect 7986 230 7999 282
rect 8051 230 8064 282
rect 8116 230 8129 282
rect 8181 230 8194 282
rect 8246 230 8259 282
rect 8311 230 8324 282
rect 8376 230 8389 282
rect 8441 230 8454 282
rect 8506 230 8519 282
rect 8571 230 8584 282
rect 8636 230 8649 282
rect 8701 230 8714 282
rect 8766 230 8779 282
rect 8831 230 8844 282
rect 8896 230 8909 282
rect 8961 230 8974 282
rect 9026 230 9039 282
rect 9091 230 9104 282
rect 9156 230 9169 282
rect 9221 230 9234 282
rect 9286 230 9299 282
rect 9351 230 9364 282
rect 9416 230 9429 282
rect 9481 230 9494 282
rect 9546 230 9559 282
rect 9611 230 9624 282
rect 9676 230 9689 282
rect 9741 230 9753 282
rect 9805 230 9817 282
rect 9869 230 9881 282
rect 9933 230 9945 282
rect 9997 230 10009 282
rect 10061 230 10073 282
rect 10125 230 10137 282
rect 10189 230 10201 282
rect 10253 230 10265 282
rect 10317 230 10329 282
rect 10381 230 10393 282
rect 10445 230 10457 282
rect 10509 230 10521 282
rect 10573 230 10585 282
rect 10637 230 10649 282
rect 10701 230 11313 282
tri 13256 241 13322 307 ne
rect 13322 241 13340 307
rect 13446 334 13679 347
rect 13713 334 13753 368
rect 13787 334 13827 368
rect 13861 334 13901 368
rect 13935 334 13974 368
rect 14008 334 14047 368
rect 14081 334 14120 368
rect 14154 334 14193 368
rect 14227 334 14266 368
rect 14300 334 14339 368
rect 14373 334 14412 368
rect 14446 334 14485 368
rect 14519 334 14531 368
rect 13446 307 14531 334
rect 14564 361 14641 387
rect 14675 361 14681 395
rect 14564 322 14681 361
rect 13446 291 13480 307
tri 13480 291 13496 307 nw
rect 13446 288 13477 291
tri 13477 288 13480 291 nw
tri 14561 288 14564 291 se
rect 14564 288 14641 322
rect 14675 288 14681 322
rect 13446 241 13458 288
tri 13458 269 13477 288 nw
tri 14542 269 14561 288 se
rect 14561 269 14681 288
tri 14529 256 14542 269 se
rect 14542 256 14681 269
tri 13322 235 13328 241 ne
rect 13328 235 13458 241
rect 13510 250 14681 256
rect 5630 225 11313 230
rect 3331 208 11313 225
rect 13510 216 13522 250
rect 13556 216 13597 250
rect 13631 216 13672 250
rect 13706 216 13747 250
rect 13781 216 13822 250
rect 13856 216 13897 250
rect 13931 216 13972 250
rect 14006 216 14047 250
rect 14081 216 14122 250
rect 14156 216 14197 250
rect 14231 216 14271 250
rect 14305 216 14345 250
rect 14379 216 14419 250
rect 14453 216 14493 250
rect 14527 216 14567 250
rect 14601 216 14681 250
rect 13510 210 14681 216
rect 3331 156 4191 208
rect 4243 156 4259 208
rect 4311 156 4327 208
rect 4379 156 4395 208
rect 4447 156 4463 208
rect 4515 156 4531 208
rect 4583 156 4599 208
rect 4651 156 4666 208
rect 4718 156 4733 208
rect 4785 156 4800 208
rect 4852 156 4867 208
rect 4919 156 4934 208
rect 4986 156 5001 208
rect 5053 156 5068 208
rect 5120 197 5659 208
rect 5120 156 5149 197
rect 3331 145 5149 156
rect 5201 145 5221 197
rect 5273 145 5293 197
rect 5345 145 5365 197
rect 5417 145 5436 197
rect 5488 145 5507 197
rect 5559 145 5578 197
rect 5630 156 5659 197
rect 5711 156 5724 208
rect 5776 156 5789 208
rect 5841 156 5854 208
rect 5906 156 5919 208
rect 5971 156 5984 208
rect 6036 156 6049 208
rect 6101 156 6114 208
rect 6166 156 6179 208
rect 6231 156 6244 208
rect 6296 156 6309 208
rect 6361 156 6374 208
rect 6426 156 6439 208
rect 6491 156 6504 208
rect 6556 156 6569 208
rect 6621 156 6634 208
rect 6686 156 6699 208
rect 6751 156 6764 208
rect 6816 156 6829 208
rect 6881 156 6894 208
rect 6946 156 6959 208
rect 7011 156 7024 208
rect 7076 156 7089 208
rect 7141 156 7154 208
rect 7206 156 7219 208
rect 7271 156 7284 208
rect 7336 156 7349 208
rect 7401 156 7414 208
rect 7466 156 7479 208
rect 7531 156 7544 208
rect 7596 156 7609 208
rect 7661 156 7674 208
rect 7726 156 7739 208
rect 7791 156 7804 208
rect 7856 156 7869 208
rect 7921 156 7934 208
rect 7986 156 7999 208
rect 8051 156 8064 208
rect 8116 156 8129 208
rect 8181 156 8194 208
rect 8246 156 8259 208
rect 8311 156 8324 208
rect 8376 156 8389 208
rect 8441 156 8454 208
rect 8506 156 8519 208
rect 8571 156 8584 208
rect 8636 156 8649 208
rect 8701 156 8714 208
rect 8766 156 8779 208
rect 8831 156 8844 208
rect 8896 156 8909 208
rect 8961 156 8974 208
rect 9026 156 9039 208
rect 9091 156 9104 208
rect 9156 156 9169 208
rect 9221 156 9234 208
rect 9286 156 9299 208
rect 9351 156 9364 208
rect 9416 156 9429 208
rect 9481 156 9494 208
rect 9546 156 9559 208
rect 9611 156 9624 208
rect 9676 156 9689 208
rect 9741 156 9753 208
rect 9805 156 9817 208
rect 9869 156 9881 208
rect 9933 156 9945 208
rect 9997 156 10009 208
rect 10061 156 10073 208
rect 10125 156 10137 208
rect 10189 156 10201 208
rect 10253 156 10265 208
rect 10317 156 10329 208
rect 10381 156 10393 208
rect 10445 156 10457 208
rect 10509 156 10521 208
rect 10573 156 10585 208
rect 10637 156 10649 208
rect 10701 156 11313 208
rect 5630 145 11313 156
rect 3331 134 11313 145
rect 3331 82 4191 134
rect 4243 82 4259 134
rect 4311 82 4327 134
rect 4379 82 4395 134
rect 4447 82 4463 134
rect 4515 82 4531 134
rect 4583 82 4599 134
rect 4651 82 4666 134
rect 4718 82 4733 134
rect 4785 82 4800 134
rect 4852 82 4867 134
rect 4919 82 4934 134
rect 4986 82 5001 134
rect 5053 82 5068 134
rect 5120 117 5659 134
rect 5120 82 5149 117
rect 3331 65 5149 82
rect 5201 65 5221 117
rect 5273 65 5293 117
rect 5345 65 5365 117
rect 5417 65 5436 117
rect 5488 65 5507 117
rect 5559 65 5578 117
rect 5630 82 5659 117
rect 5711 82 5724 134
rect 5776 82 5789 134
rect 5841 82 5854 134
rect 5906 82 5919 134
rect 5971 82 5984 134
rect 6036 82 6049 134
rect 6101 82 6114 134
rect 6166 82 6179 134
rect 6231 82 6244 134
rect 6296 82 6309 134
rect 6361 82 6374 134
rect 6426 82 6439 134
rect 6491 82 6504 134
rect 6556 82 6569 134
rect 6621 82 6634 134
rect 6686 82 6699 134
rect 6751 82 6764 134
rect 6816 82 6829 134
rect 6881 82 6894 134
rect 6946 82 6959 134
rect 7011 82 7024 134
rect 7076 82 7089 134
rect 7141 82 7154 134
rect 7206 82 7219 134
rect 7271 82 7284 134
rect 7336 82 7349 134
rect 7401 82 7414 134
rect 7466 82 7479 134
rect 7531 82 7544 134
rect 7596 82 7609 134
rect 7661 82 7674 134
rect 7726 82 7739 134
rect 7791 82 7804 134
rect 7856 82 7869 134
rect 7921 82 7934 134
rect 7986 82 7999 134
rect 8051 82 8064 134
rect 8116 82 8129 134
rect 8181 82 8194 134
rect 8246 82 8259 134
rect 8311 82 8324 134
rect 8376 82 8389 134
rect 8441 82 8454 134
rect 8506 82 8519 134
rect 8571 82 8584 134
rect 8636 82 8649 134
rect 8701 82 8714 134
rect 8766 82 8779 134
rect 8831 82 8844 134
rect 8896 82 8909 134
rect 8961 82 8974 134
rect 9026 82 9039 134
rect 9091 82 9104 134
rect 9156 82 9169 134
rect 9221 82 9234 134
rect 9286 82 9299 134
rect 9351 82 9364 134
rect 9416 82 9429 134
rect 9481 82 9494 134
rect 9546 82 9559 134
rect 9611 82 9624 134
rect 9676 82 9689 134
rect 9741 82 9753 134
rect 9805 82 9817 134
rect 9869 82 9881 134
rect 9933 82 9945 134
rect 9997 82 10009 134
rect 10061 82 10073 134
rect 10125 82 10137 134
rect 10189 82 10201 134
rect 10253 82 10265 134
rect 10317 82 10329 134
rect 10381 82 10393 134
rect 10445 82 10457 134
rect 10509 82 10521 134
rect 10573 82 10585 134
rect 10637 82 10649 134
rect 10701 82 11313 134
rect 5630 65 11313 82
rect 3331 60 5161 65
rect 3331 8 4191 60
rect 4243 8 4259 60
rect 4311 8 4327 60
rect 4379 8 4395 60
rect 4447 8 4463 60
rect 4515 8 4531 60
rect 4583 8 4599 60
rect 4651 8 4666 60
rect 4718 8 4733 60
rect 4785 8 4800 60
rect 4852 8 4867 60
rect 4919 8 4934 60
rect 4986 8 5001 60
rect 5053 8 5068 60
rect 5120 34 5161 60
tri 5161 34 5192 65 nw
rect 5590 64 11313 65
tri 5590 34 5620 64 ne
rect 5620 60 11313 64
rect 5620 34 5659 60
rect 5120 8 5134 34
rect 3331 7 5134 8
tri 5134 7 5161 34 nw
rect 3331 0 5127 7
tri 5127 0 5134 7 nw
rect 5242 0 5540 34
tri 5620 7 5647 34 ne
rect 5647 8 5659 34
rect 5711 8 5724 60
rect 5776 8 5789 60
rect 5841 8 5854 60
rect 5906 8 5919 60
rect 5971 8 5984 60
rect 6036 8 6049 60
rect 6101 8 6114 60
rect 6166 8 6179 60
rect 6231 8 6244 60
rect 6296 8 6309 60
rect 6361 8 6374 60
rect 6426 8 6439 60
rect 6491 8 6504 60
rect 6556 8 6569 60
rect 6621 8 6634 60
rect 6686 8 6699 60
rect 6751 8 6764 60
rect 6816 8 6829 60
rect 6881 8 6894 60
rect 6946 8 6959 60
rect 7011 8 7024 60
rect 7076 8 7089 60
rect 7141 8 7154 60
rect 7206 8 7219 60
rect 7271 8 7284 60
rect 7336 8 7349 60
rect 7401 8 7414 60
rect 7466 8 7479 60
rect 7531 8 7544 60
rect 7596 8 7609 60
rect 7661 8 7674 60
rect 7726 8 7739 60
rect 7791 8 7804 60
rect 7856 8 7869 60
rect 7921 8 7934 60
rect 7986 8 7999 60
rect 8051 8 8064 60
rect 8116 8 8129 60
rect 8181 8 8194 60
rect 8246 8 8259 60
rect 8311 8 8324 60
rect 8376 8 8389 60
rect 8441 8 8454 60
rect 8506 8 8519 60
rect 8571 8 8584 60
rect 8636 8 8649 60
rect 8701 8 8714 60
rect 8766 8 8779 60
rect 8831 8 8844 60
rect 8896 8 8909 60
rect 8961 8 8974 60
rect 9026 8 9039 60
rect 9091 8 9104 60
rect 9156 8 9169 60
rect 9221 8 9234 60
rect 9286 8 9299 60
rect 9351 8 9364 60
rect 9416 8 9429 60
rect 9481 8 9494 60
rect 9546 8 9559 60
rect 9611 8 9624 60
rect 9676 8 9689 60
rect 9741 8 9753 60
rect 9805 8 9817 60
rect 9869 8 9881 60
rect 9933 8 9945 60
rect 9997 8 10009 60
rect 10061 8 10073 60
rect 10125 8 10137 60
rect 10189 8 10201 60
rect 10253 8 10265 60
rect 10317 8 10329 60
rect 10381 8 10393 60
rect 10445 8 10457 60
rect 10509 8 10521 60
rect 10573 8 10585 60
rect 10637 8 10649 60
rect 10701 8 11313 60
rect 5647 7 11313 8
tri 5647 0 5654 7 ne
rect 5654 0 11313 7
<< via1 >>
rect 2249 38700 2253 38720
rect 2253 38700 2291 38720
rect 2291 38700 2301 38720
rect 2315 38700 2325 38720
rect 2325 38701 2363 38720
rect 2363 38701 2367 38720
rect 2325 38700 2367 38701
rect 2249 38668 2301 38700
rect 2315 38668 2367 38700
rect 2249 38627 2253 38656
rect 2253 38627 2291 38656
rect 2291 38627 2301 38656
rect 2315 38627 2325 38656
rect 2325 38628 2363 38656
rect 2363 38628 2367 38656
rect 2325 38627 2367 38628
rect 2249 38604 2301 38627
rect 2315 38604 2367 38627
rect 2249 38588 2301 38592
rect 2315 38589 2367 38592
rect 2315 38588 2363 38589
rect 2249 38554 2253 38588
rect 2253 38554 2291 38588
rect 2291 38554 2301 38588
rect 2315 38554 2325 38588
rect 2325 38555 2363 38588
rect 2363 38555 2367 38589
rect 2325 38554 2367 38555
rect 2249 38540 2301 38554
rect 2315 38540 2367 38554
rect 2249 38515 2301 38528
rect 2315 38516 2367 38528
rect 2315 38515 2363 38516
rect 2249 38481 2253 38515
rect 2253 38481 2291 38515
rect 2291 38481 2301 38515
rect 2315 38481 2325 38515
rect 2325 38482 2363 38515
rect 2363 38482 2367 38516
rect 2325 38481 2367 38482
rect 2249 38476 2301 38481
rect 2315 38476 2367 38481
rect 2249 38442 2301 38464
rect 2315 38443 2367 38464
rect 2315 38442 2363 38443
rect 2249 38412 2253 38442
rect 2253 38412 2291 38442
rect 2291 38412 2301 38442
rect 2315 38412 2325 38442
rect 2325 38412 2363 38442
rect 2363 38412 2367 38443
rect 2249 38369 2301 38400
rect 2315 38370 2367 38400
rect 2315 38369 2363 38370
rect 2249 38348 2253 38369
rect 2253 38348 2291 38369
rect 2291 38348 2301 38369
rect 2315 38348 2325 38369
rect 2325 38348 2363 38369
rect 2363 38348 2367 38370
rect 2249 38335 2253 38336
rect 2253 38335 2291 38336
rect 2291 38335 2301 38336
rect 2315 38335 2325 38336
rect 2325 38335 2367 38336
rect 2249 38296 2301 38335
rect 2315 38297 2367 38335
rect 2315 38296 2363 38297
rect 2249 38284 2253 38296
rect 2253 38284 2291 38296
rect 2291 38284 2301 38296
rect 2315 38284 2325 38296
rect 2325 38284 2363 38296
rect 2363 38284 2367 38297
rect 2249 38262 2253 38272
rect 2253 38262 2291 38272
rect 2291 38262 2301 38272
rect 2315 38262 2325 38272
rect 2325 38263 2363 38272
rect 2363 38263 2367 38272
rect 2325 38262 2367 38263
rect 2249 38223 2301 38262
rect 2315 38224 2367 38262
rect 2315 38223 2363 38224
rect 2249 38220 2253 38223
rect 2253 38220 2291 38223
rect 2291 38220 2301 38223
rect 2315 38220 2325 38223
rect 2325 38220 2363 38223
rect 2363 38220 2367 38224
rect 2249 38189 2253 38208
rect 2253 38189 2291 38208
rect 2291 38189 2301 38208
rect 2315 38189 2325 38208
rect 2325 38190 2363 38208
rect 2363 38190 2367 38208
rect 2325 38189 2367 38190
rect 2249 38156 2301 38189
rect 2315 38156 2367 38189
rect 2249 38116 2253 38144
rect 2253 38116 2291 38144
rect 2291 38116 2301 38144
rect 2315 38116 2325 38144
rect 2325 38117 2363 38144
rect 2363 38117 2367 38144
rect 2325 38116 2367 38117
rect 2249 38092 2301 38116
rect 2315 38092 2367 38116
rect 2249 38077 2301 38080
rect 2315 38078 2367 38080
rect 2315 38077 2363 38078
rect 2249 38043 2253 38077
rect 2253 38043 2291 38077
rect 2291 38043 2301 38077
rect 2315 38043 2325 38077
rect 2325 38044 2363 38077
rect 2363 38044 2367 38078
rect 2325 38043 2367 38044
rect 2249 38028 2301 38043
rect 2315 38028 2367 38043
rect 2249 38004 2301 38016
rect 2315 38005 2367 38016
rect 2315 38004 2363 38005
rect 2249 37970 2253 38004
rect 2253 37970 2291 38004
rect 2291 37970 2301 38004
rect 2315 37970 2325 38004
rect 2325 37971 2363 38004
rect 2363 37971 2367 38005
rect 2325 37970 2367 37971
rect 2249 37964 2301 37970
rect 2315 37964 2367 37970
rect 2249 37931 2301 37952
rect 2315 37932 2367 37952
rect 2315 37931 2363 37932
rect 2249 37900 2253 37931
rect 2253 37900 2291 37931
rect 2291 37900 2301 37931
rect 2315 37900 2325 37931
rect 2325 37900 2363 37931
rect 2363 37900 2367 37932
rect 2249 37858 2301 37888
rect 2315 37859 2367 37888
rect 2315 37858 2363 37859
rect 2249 37836 2253 37858
rect 2253 37836 2291 37858
rect 2291 37836 2301 37858
rect 2315 37836 2325 37858
rect 2325 37836 2363 37858
rect 2363 37836 2367 37859
rect 2249 37785 2301 37824
rect 2315 37786 2367 37824
rect 2315 37785 2363 37786
rect 2249 37772 2253 37785
rect 2253 37772 2291 37785
rect 2291 37772 2301 37785
rect 2315 37772 2325 37785
rect 2325 37772 2363 37785
rect 2363 37772 2367 37786
rect 2249 37751 2253 37760
rect 2253 37751 2291 37760
rect 2291 37751 2301 37760
rect 2315 37751 2325 37760
rect 2325 37752 2363 37760
rect 2363 37752 2367 37760
rect 2325 37751 2367 37752
rect 2249 37712 2301 37751
rect 2315 37713 2367 37751
rect 2315 37712 2363 37713
rect 2249 37708 2253 37712
rect 2253 37708 2291 37712
rect 2291 37708 2301 37712
rect 2315 37708 2325 37712
rect 2325 37708 2363 37712
rect 2363 37708 2367 37713
rect 2249 37678 2253 37696
rect 2253 37678 2291 37696
rect 2291 37678 2301 37696
rect 2315 37678 2325 37696
rect 2325 37679 2363 37696
rect 2363 37679 2367 37696
rect 2325 37678 2367 37679
rect 2249 37644 2301 37678
rect 2315 37644 2367 37678
rect 2249 37605 2253 37632
rect 2253 37605 2291 37632
rect 2291 37605 2301 37632
rect 2315 37605 2325 37632
rect 2325 37606 2363 37632
rect 2363 37606 2367 37632
rect 2325 37605 2367 37606
rect 2249 37580 2301 37605
rect 2315 37580 2367 37605
rect 2249 37566 2301 37568
rect 2315 37567 2367 37568
rect 2315 37566 2363 37567
rect 2249 37532 2253 37566
rect 2253 37532 2291 37566
rect 2291 37532 2301 37566
rect 2315 37532 2325 37566
rect 2325 37533 2363 37566
rect 2363 37533 2367 37567
rect 2325 37532 2367 37533
rect 2249 37516 2301 37532
rect 2315 37516 2367 37532
rect 2249 37493 2301 37504
rect 2315 37494 2367 37504
rect 2315 37493 2363 37494
rect 2249 37459 2253 37493
rect 2253 37459 2291 37493
rect 2291 37459 2301 37493
rect 2315 37459 2325 37493
rect 2325 37460 2363 37493
rect 2363 37460 2367 37494
rect 2325 37459 2367 37460
rect 2249 37452 2301 37459
rect 2315 37452 2367 37459
rect 2249 37420 2301 37440
rect 2315 37421 2367 37440
rect 2315 37420 2363 37421
rect 2249 37388 2253 37420
rect 2253 37388 2291 37420
rect 2291 37388 2301 37420
rect 2315 37388 2325 37420
rect 2325 37388 2363 37420
rect 2363 37388 2367 37421
rect 2249 37347 2301 37376
rect 2315 37348 2367 37376
rect 2315 37347 2363 37348
rect 2249 37324 2253 37347
rect 2253 37324 2291 37347
rect 2291 37324 2301 37347
rect 2315 37324 2325 37347
rect 2325 37324 2363 37347
rect 2363 37324 2367 37348
rect 2249 37274 2301 37312
rect 2315 37275 2367 37312
rect 2315 37274 2363 37275
rect 2249 37260 2253 37274
rect 2253 37260 2291 37274
rect 2291 37260 2301 37274
rect 2315 37260 2325 37274
rect 2325 37260 2363 37274
rect 2363 37260 2367 37275
rect 2249 37240 2253 37248
rect 2253 37240 2291 37248
rect 2291 37240 2301 37248
rect 2315 37240 2325 37248
rect 2325 37241 2363 37248
rect 2363 37241 2367 37248
rect 2325 37240 2367 37241
rect 2249 37201 2301 37240
rect 2315 37202 2367 37240
rect 2315 37201 2363 37202
rect 2249 37196 2253 37201
rect 2253 37196 2291 37201
rect 2291 37196 2301 37201
rect 2315 37196 2325 37201
rect 2325 37196 2363 37201
rect 2363 37196 2367 37202
rect 2249 37167 2253 37184
rect 2253 37167 2291 37184
rect 2291 37167 2301 37184
rect 2315 37167 2325 37184
rect 2325 37168 2363 37184
rect 2363 37168 2367 37184
rect 2325 37167 2367 37168
rect 2249 37132 2301 37167
rect 2315 37132 2367 37167
rect 2249 37094 2253 37120
rect 2253 37094 2291 37120
rect 2291 37094 2301 37120
rect 2315 37094 2325 37120
rect 2325 37095 2363 37120
rect 2363 37095 2367 37120
rect 2325 37094 2367 37095
rect 2249 37068 2301 37094
rect 2315 37068 2367 37094
rect 2249 37055 2301 37056
rect 2315 37055 2363 37056
rect 2249 37021 2253 37055
rect 2253 37021 2291 37055
rect 2291 37021 2301 37055
rect 2315 37021 2325 37055
rect 2325 37022 2363 37055
rect 2363 37022 2367 37056
rect 2325 37021 2367 37022
rect 2249 37004 2301 37021
rect 2315 37004 2367 37021
rect 2249 36982 2301 36992
rect 2315 36983 2367 36992
rect 2315 36982 2363 36983
rect 2249 36948 2253 36982
rect 2253 36948 2291 36982
rect 2291 36948 2301 36982
rect 2315 36948 2325 36982
rect 2325 36949 2363 36982
rect 2363 36949 2367 36983
rect 2325 36948 2367 36949
rect 2249 36940 2301 36948
rect 2315 36940 2367 36948
rect 2249 36909 2301 36928
rect 2315 36910 2367 36928
rect 2315 36909 2363 36910
rect 2249 36876 2253 36909
rect 2253 36876 2291 36909
rect 2291 36876 2301 36909
rect 2315 36876 2325 36909
rect 2325 36876 2363 36909
rect 2363 36876 2367 36910
rect 2249 36836 2301 36864
rect 2315 36837 2367 36864
rect 2315 36836 2363 36837
rect 2249 36812 2253 36836
rect 2253 36812 2291 36836
rect 2291 36812 2301 36836
rect 2315 36812 2325 36836
rect 2325 36812 2363 36836
rect 2363 36812 2367 36837
rect 2249 36763 2301 36800
rect 2315 36764 2367 36800
rect 2315 36763 2363 36764
rect 2249 36748 2253 36763
rect 2253 36748 2291 36763
rect 2291 36748 2301 36763
rect 2315 36748 2325 36763
rect 2325 36748 2363 36763
rect 2363 36748 2367 36764
rect 2249 36729 2253 36736
rect 2253 36729 2291 36736
rect 2291 36729 2301 36736
rect 2315 36729 2325 36736
rect 2325 36730 2363 36736
rect 2363 36730 2367 36736
rect 2325 36729 2367 36730
rect 2249 36690 2301 36729
rect 2315 36691 2367 36729
rect 2878 38854 2930 38886
rect 2878 38834 2884 38854
rect 2884 38834 2918 38854
rect 2918 38834 2930 38854
rect 2943 38854 2995 38886
rect 2943 38834 2957 38854
rect 2957 38834 2991 38854
rect 2991 38834 2995 38854
rect 3008 38854 3060 38886
rect 3073 38854 3125 38886
rect 3138 38854 3190 38886
rect 3203 38854 3255 38886
rect 3268 38854 3320 38886
rect 3332 38854 3384 38886
rect 3396 38854 3448 38886
rect 3008 38834 3030 38854
rect 3030 38834 3060 38854
rect 3073 38834 3103 38854
rect 3103 38834 3125 38854
rect 3138 38834 3176 38854
rect 3176 38834 3190 38854
rect 3203 38834 3210 38854
rect 3210 38834 3249 38854
rect 3249 38834 3255 38854
rect 3268 38834 3283 38854
rect 3283 38834 3320 38854
rect 3332 38834 3356 38854
rect 3356 38834 3384 38854
rect 3396 38834 3429 38854
rect 3429 38834 3448 38854
rect 3460 38854 3512 38886
rect 3460 38834 3468 38854
rect 3468 38834 3502 38854
rect 3502 38834 3512 38854
rect 3524 38854 3576 38886
rect 3524 38834 3541 38854
rect 3541 38834 3575 38854
rect 3575 38834 3576 38854
rect 3588 38854 3640 38886
rect 3652 38854 3704 38886
rect 3716 38854 3768 38886
rect 3780 38854 3832 38886
rect 3844 38854 3896 38886
rect 3908 38854 3960 38886
rect 3588 38834 3614 38854
rect 3614 38834 3640 38854
rect 3652 38834 3687 38854
rect 3687 38834 3704 38854
rect 3716 38834 3721 38854
rect 3721 38834 3760 38854
rect 3760 38834 3768 38854
rect 3780 38834 3794 38854
rect 3794 38834 3832 38854
rect 3844 38834 3867 38854
rect 3867 38834 3896 38854
rect 3908 38834 3940 38854
rect 3940 38834 3960 38854
rect 3972 38854 4024 38886
rect 3972 38834 3979 38854
rect 3979 38834 4013 38854
rect 4013 38834 4024 38854
rect 4036 38854 4088 38886
rect 4036 38834 4052 38854
rect 4052 38834 4086 38854
rect 4086 38834 4088 38854
rect 4100 38854 4152 38886
rect 4164 38854 4216 38886
rect 4228 38854 4280 38886
rect 4292 38854 4344 38886
rect 4356 38854 4408 38886
rect 4420 38854 4472 38886
rect 4100 38834 4125 38854
rect 4125 38834 4152 38854
rect 4164 38834 4198 38854
rect 4198 38834 4216 38854
rect 4228 38834 4232 38854
rect 4232 38834 4271 38854
rect 4271 38834 4280 38854
rect 4292 38834 4305 38854
rect 4305 38834 4344 38854
rect 4356 38834 4378 38854
rect 4378 38834 4408 38854
rect 4420 38834 4451 38854
rect 4451 38834 4472 38854
rect 4484 38854 4536 38886
rect 4484 38834 4490 38854
rect 4490 38834 4524 38854
rect 4524 38834 4536 38854
rect 4548 38854 4600 38886
rect 4548 38834 4563 38854
rect 4563 38834 4597 38854
rect 4597 38834 4600 38854
rect 4612 38854 4664 38886
rect 4676 38854 4728 38886
rect 4740 38854 4792 38886
rect 4804 38854 4856 38886
rect 4868 38854 4920 38886
rect 4932 38854 4984 38886
rect 4612 38834 4636 38854
rect 4636 38834 4664 38854
rect 4676 38834 4709 38854
rect 4709 38834 4728 38854
rect 4740 38834 4743 38854
rect 4743 38834 4782 38854
rect 4782 38834 4792 38854
rect 4804 38834 4816 38854
rect 4816 38834 4855 38854
rect 4855 38834 4856 38854
rect 4868 38834 4889 38854
rect 4889 38834 4920 38854
rect 4932 38834 4962 38854
rect 4962 38834 4984 38854
rect 4996 38854 5048 38886
rect 4996 38834 5001 38854
rect 5001 38834 5035 38854
rect 5035 38834 5048 38854
rect 5060 38854 5112 38886
rect 5060 38834 5074 38854
rect 5074 38834 5108 38854
rect 5108 38834 5112 38854
rect 5124 38854 5176 38886
rect 5188 38854 5240 38886
rect 5252 38854 5304 38886
rect 5316 38854 5368 38886
rect 5380 38854 5432 38886
rect 5444 38854 5496 38886
rect 5124 38834 5147 38854
rect 5147 38834 5176 38854
rect 5188 38834 5220 38854
rect 5220 38834 5240 38854
rect 5252 38834 5254 38854
rect 5254 38834 5293 38854
rect 5293 38834 5304 38854
rect 5316 38834 5327 38854
rect 5327 38834 5366 38854
rect 5366 38834 5368 38854
rect 5380 38834 5400 38854
rect 5400 38834 5432 38854
rect 5444 38834 5473 38854
rect 5473 38834 5496 38854
rect 5508 38854 5560 38886
rect 5508 38834 5512 38854
rect 5512 38834 5546 38854
rect 5546 38834 5560 38854
rect 5572 38854 5624 38886
rect 5572 38834 5584 38854
rect 5584 38834 5618 38854
rect 5618 38834 5624 38854
rect 5636 38854 5688 38886
rect 5700 38854 5752 38886
rect 5764 38854 5816 38886
rect 5828 38854 5880 38886
rect 5892 38854 5944 38886
rect 5956 38854 6008 38886
rect 6020 38854 6072 38886
rect 5636 38834 5656 38854
rect 5656 38834 5688 38854
rect 5700 38834 5728 38854
rect 5728 38834 5752 38854
rect 5764 38834 5800 38854
rect 5800 38834 5816 38854
rect 5828 38834 5834 38854
rect 5834 38834 5872 38854
rect 5872 38834 5880 38854
rect 5892 38834 5906 38854
rect 5906 38834 5944 38854
rect 5956 38834 5978 38854
rect 5978 38834 6008 38854
rect 6020 38834 6050 38854
rect 6050 38834 6072 38854
rect 6084 38854 6136 38886
rect 6084 38834 6088 38854
rect 6088 38834 6122 38854
rect 6122 38834 6136 38854
rect 6148 38854 6200 38886
rect 6148 38834 6160 38854
rect 6160 38834 6194 38854
rect 6194 38834 6200 38854
rect 6212 38854 6264 38886
rect 6276 38854 6328 38886
rect 6340 38854 6392 38886
rect 6404 38854 6456 38886
rect 6468 38854 6520 38886
rect 6532 38854 6584 38886
rect 6596 38854 6648 38886
rect 6212 38834 6232 38854
rect 6232 38834 6264 38854
rect 6276 38834 6304 38854
rect 6304 38834 6328 38854
rect 6340 38834 6376 38854
rect 6376 38834 6392 38854
rect 6404 38834 6410 38854
rect 6410 38834 6448 38854
rect 6448 38834 6456 38854
rect 6468 38834 6482 38854
rect 6482 38834 6520 38854
rect 6532 38834 6554 38854
rect 6554 38834 6584 38854
rect 6596 38834 6626 38854
rect 6626 38834 6648 38854
rect 6660 38854 6712 38886
rect 6660 38834 6664 38854
rect 6664 38834 6698 38854
rect 6698 38834 6712 38854
rect 6724 38854 6776 38886
rect 6724 38834 6736 38854
rect 6736 38834 6770 38854
rect 6770 38834 6776 38854
rect 6788 38854 6840 38886
rect 6852 38854 6904 38886
rect 6916 38854 6968 38886
rect 6980 38854 7032 38886
rect 7044 38854 7096 38886
rect 7108 38854 7160 38886
rect 7172 38854 7224 38886
rect 6788 38834 6808 38854
rect 6808 38834 6840 38854
rect 6852 38834 6880 38854
rect 6880 38834 6904 38854
rect 6916 38834 6952 38854
rect 6952 38834 6968 38854
rect 6980 38834 6986 38854
rect 6986 38834 7024 38854
rect 7024 38834 7032 38854
rect 7044 38834 7058 38854
rect 7058 38834 7096 38854
rect 7108 38834 7130 38854
rect 7130 38834 7160 38854
rect 7172 38834 7202 38854
rect 7202 38834 7224 38854
rect 7236 38854 7288 38886
rect 7236 38834 7240 38854
rect 7240 38834 7274 38854
rect 7274 38834 7288 38854
rect 7300 38854 7352 38886
rect 7300 38834 7312 38854
rect 7312 38834 7346 38854
rect 7346 38834 7352 38854
rect 7364 38854 7416 38886
rect 7428 38854 7480 38886
rect 7492 38854 7544 38886
rect 7556 38854 7608 38886
rect 7620 38854 7672 38886
rect 7684 38854 7736 38886
rect 7748 38854 7800 38886
rect 7364 38834 7384 38854
rect 7384 38834 7416 38854
rect 7428 38834 7456 38854
rect 7456 38834 7480 38854
rect 7492 38834 7528 38854
rect 7528 38834 7544 38854
rect 7556 38834 7562 38854
rect 7562 38834 7600 38854
rect 7600 38834 7608 38854
rect 7620 38834 7634 38854
rect 7634 38834 7672 38854
rect 7684 38834 7706 38854
rect 7706 38834 7736 38854
rect 7748 38834 7778 38854
rect 7778 38834 7800 38854
rect 7812 38854 7864 38886
rect 7812 38834 7816 38854
rect 7816 38834 7850 38854
rect 7850 38834 7864 38854
rect 7876 38854 7928 38886
rect 7876 38834 7888 38854
rect 7888 38834 7922 38854
rect 7922 38834 7928 38854
rect 7940 38854 7992 38886
rect 8004 38854 8056 38886
rect 8068 38854 8120 38886
rect 8132 38854 8184 38886
rect 8196 38854 8248 38886
rect 8260 38854 8312 38886
rect 8324 38854 8376 38886
rect 7940 38834 7960 38854
rect 7960 38834 7992 38854
rect 8004 38834 8032 38854
rect 8032 38834 8056 38854
rect 8068 38834 8104 38854
rect 8104 38834 8120 38854
rect 8132 38834 8138 38854
rect 8138 38834 8176 38854
rect 8176 38834 8184 38854
rect 8196 38834 8210 38854
rect 8210 38834 8248 38854
rect 8260 38834 8282 38854
rect 8282 38834 8312 38854
rect 8324 38834 8354 38854
rect 8354 38834 8376 38854
rect 8388 38854 8440 38886
rect 8388 38834 8392 38854
rect 8392 38834 8426 38854
rect 8426 38834 8440 38854
rect 8452 38854 8504 38886
rect 8452 38834 8464 38854
rect 8464 38834 8498 38854
rect 8498 38834 8504 38854
rect 8516 38854 8568 38886
rect 8580 38854 8632 38886
rect 8644 38854 8696 38886
rect 8708 38854 8760 38886
rect 8772 38854 8824 38886
rect 8836 38854 8888 38886
rect 8900 38854 8952 38886
rect 8516 38834 8536 38854
rect 8536 38834 8568 38854
rect 8580 38834 8608 38854
rect 8608 38834 8632 38854
rect 8644 38834 8680 38854
rect 8680 38834 8696 38854
rect 8708 38834 8714 38854
rect 8714 38834 8752 38854
rect 8752 38834 8760 38854
rect 8772 38834 8786 38854
rect 8786 38834 8824 38854
rect 8836 38834 8858 38854
rect 8858 38834 8888 38854
rect 8900 38834 8930 38854
rect 8930 38834 8952 38854
rect 8964 38854 9016 38886
rect 8964 38834 8968 38854
rect 8968 38834 9002 38854
rect 9002 38834 9016 38854
rect 9028 38854 9080 38886
rect 9028 38834 9040 38854
rect 9040 38834 9074 38854
rect 9074 38834 9080 38854
rect 9092 38854 9144 38886
rect 9156 38854 9208 38886
rect 9220 38854 9272 38886
rect 9284 38854 9336 38886
rect 9348 38854 9400 38886
rect 9412 38854 9464 38886
rect 9476 38854 9528 38886
rect 9092 38834 9112 38854
rect 9112 38834 9144 38854
rect 9156 38834 9184 38854
rect 9184 38834 9208 38854
rect 9220 38834 9256 38854
rect 9256 38834 9272 38854
rect 9284 38834 9290 38854
rect 9290 38834 9328 38854
rect 9328 38834 9336 38854
rect 9348 38834 9362 38854
rect 9362 38834 9400 38854
rect 9412 38834 9434 38854
rect 9434 38834 9464 38854
rect 9476 38834 9506 38854
rect 9506 38834 9528 38854
rect 9540 38854 9592 38886
rect 9540 38834 9544 38854
rect 9544 38834 9578 38854
rect 9578 38834 9592 38854
rect 9604 38854 9656 38886
rect 9604 38834 9616 38854
rect 9616 38834 9650 38854
rect 9650 38834 9656 38854
rect 9668 38854 9720 38886
rect 9732 38854 9784 38886
rect 9796 38854 9848 38886
rect 9860 38854 9912 38886
rect 9924 38854 9976 38886
rect 9988 38854 10040 38886
rect 10052 38854 10104 38886
rect 9668 38834 9688 38854
rect 9688 38834 9720 38854
rect 9732 38834 9760 38854
rect 9760 38834 9784 38854
rect 9796 38834 9832 38854
rect 9832 38834 9848 38854
rect 9860 38834 9866 38854
rect 9866 38834 9904 38854
rect 9904 38834 9912 38854
rect 9924 38834 9938 38854
rect 9938 38834 9976 38854
rect 9988 38834 10010 38854
rect 10010 38834 10040 38854
rect 10052 38834 10082 38854
rect 10082 38834 10104 38854
rect 10116 38854 10168 38886
rect 10116 38834 10120 38854
rect 10120 38834 10154 38854
rect 10154 38834 10168 38854
rect 10180 38854 10232 38886
rect 10180 38834 10192 38854
rect 10192 38834 10226 38854
rect 10226 38834 10232 38854
rect 10244 38854 10296 38886
rect 10308 38854 10360 38886
rect 10372 38854 10424 38886
rect 10436 38854 10488 38886
rect 10500 38854 10552 38886
rect 10564 38854 10616 38886
rect 10628 38854 10680 38886
rect 10244 38834 10264 38854
rect 10264 38834 10296 38854
rect 10308 38834 10336 38854
rect 10336 38834 10360 38854
rect 10372 38834 10408 38854
rect 10408 38834 10424 38854
rect 10436 38834 10442 38854
rect 10442 38834 10480 38854
rect 10480 38834 10488 38854
rect 10500 38834 10514 38854
rect 10514 38834 10552 38854
rect 10564 38834 10586 38854
rect 10586 38834 10616 38854
rect 10628 38834 10658 38854
rect 10658 38834 10680 38854
rect 10692 38854 10744 38886
rect 10692 38834 10696 38854
rect 10696 38834 10730 38854
rect 10730 38834 10744 38854
rect 10756 38854 10808 38886
rect 10756 38834 10768 38854
rect 10768 38834 10802 38854
rect 10802 38834 10808 38854
rect 10820 38854 10872 38886
rect 10884 38854 10936 38886
rect 10948 38854 11000 38886
rect 11012 38854 11064 38886
rect 11076 38854 11128 38886
rect 11140 38854 11192 38886
rect 11204 38854 11256 38886
rect 10820 38834 10840 38854
rect 10840 38834 10872 38854
rect 10884 38834 10912 38854
rect 10912 38834 10936 38854
rect 10948 38834 10984 38854
rect 10984 38834 11000 38854
rect 11012 38834 11018 38854
rect 11018 38834 11056 38854
rect 11056 38834 11064 38854
rect 11076 38834 11090 38854
rect 11090 38834 11128 38854
rect 11140 38834 11162 38854
rect 11162 38834 11192 38854
rect 11204 38834 11234 38854
rect 11234 38834 11256 38854
rect 11268 38854 11320 38886
rect 11268 38834 11272 38854
rect 11272 38834 11306 38854
rect 11306 38834 11320 38854
rect 11332 38854 11384 38886
rect 11332 38834 11344 38854
rect 11344 38834 11378 38854
rect 11378 38834 11384 38854
rect 11396 38854 11448 38886
rect 11460 38854 11512 38886
rect 11524 38854 11576 38886
rect 11588 38854 11640 38886
rect 11652 38854 11704 38886
rect 11716 38854 11768 38886
rect 11780 38854 11832 38886
rect 11396 38834 11416 38854
rect 11416 38834 11448 38854
rect 11460 38834 11488 38854
rect 11488 38834 11512 38854
rect 11524 38834 11560 38854
rect 11560 38834 11576 38854
rect 11588 38834 11594 38854
rect 11594 38834 11632 38854
rect 11632 38834 11640 38854
rect 11652 38834 11666 38854
rect 11666 38834 11704 38854
rect 11716 38834 11738 38854
rect 11738 38834 11768 38854
rect 11780 38834 11810 38854
rect 11810 38834 11832 38854
rect 11844 38854 11896 38886
rect 11844 38834 11848 38854
rect 11848 38834 11882 38854
rect 11882 38834 11896 38854
rect 11908 38854 11960 38886
rect 11908 38834 11920 38854
rect 11920 38834 11954 38854
rect 11954 38834 11960 38854
rect 11972 38854 12024 38886
rect 12036 38854 12088 38886
rect 12100 38854 12152 38886
rect 12164 38854 12216 38886
rect 12228 38854 12280 38886
rect 12292 38854 12344 38886
rect 12356 38854 12408 38886
rect 11972 38834 11992 38854
rect 11992 38834 12024 38854
rect 12036 38834 12064 38854
rect 12064 38834 12088 38854
rect 12100 38834 12136 38854
rect 12136 38834 12152 38854
rect 12164 38834 12170 38854
rect 12170 38834 12208 38854
rect 12208 38834 12216 38854
rect 12228 38834 12242 38854
rect 12242 38834 12280 38854
rect 12292 38834 12314 38854
rect 12314 38834 12344 38854
rect 12356 38834 12386 38854
rect 12386 38834 12408 38854
rect 12420 38854 12472 38886
rect 12420 38834 12424 38854
rect 12424 38834 12458 38854
rect 12458 38834 12472 38854
rect 12484 38854 12536 38886
rect 12484 38834 12496 38854
rect 12496 38834 12530 38854
rect 12530 38834 12536 38854
rect 12548 38854 12600 38886
rect 12612 38854 12664 38886
rect 12676 38854 12728 38886
rect 12740 38854 12792 38886
rect 12804 38854 12856 38886
rect 12868 38854 12920 38886
rect 12932 38854 12984 38886
rect 12548 38834 12568 38854
rect 12568 38834 12600 38854
rect 12612 38834 12640 38854
rect 12640 38834 12664 38854
rect 12676 38834 12712 38854
rect 12712 38834 12728 38854
rect 12740 38834 12746 38854
rect 12746 38834 12784 38854
rect 12784 38834 12792 38854
rect 12804 38834 12818 38854
rect 12818 38834 12856 38854
rect 12868 38834 12890 38854
rect 12890 38834 12920 38854
rect 12932 38834 12962 38854
rect 12962 38834 12984 38854
rect 12996 38854 13048 38886
rect 12996 38834 13000 38854
rect 13000 38834 13034 38854
rect 13034 38834 13048 38854
rect 13060 38854 13112 38886
rect 13060 38834 13072 38854
rect 13072 38834 13106 38854
rect 13106 38834 13112 38854
rect 2673 38714 2725 38720
rect 2673 38680 2679 38714
rect 2679 38680 2713 38714
rect 2713 38680 2725 38714
rect 2673 38668 2725 38680
rect 2739 38714 2791 38720
rect 2739 38680 2751 38714
rect 2751 38680 2785 38714
rect 2785 38680 2791 38714
rect 2739 38668 2791 38680
rect 2673 38641 2725 38656
rect 2673 38607 2679 38641
rect 2679 38607 2713 38641
rect 2713 38607 2725 38641
rect 2673 38604 2725 38607
rect 2739 38641 2791 38656
rect 2739 38607 2751 38641
rect 2751 38607 2785 38641
rect 2785 38607 2791 38641
rect 2739 38604 2791 38607
rect 2673 38568 2725 38592
rect 2673 38540 2679 38568
rect 2679 38540 2713 38568
rect 2713 38540 2725 38568
rect 2739 38568 2791 38592
rect 2739 38540 2751 38568
rect 2751 38540 2785 38568
rect 2785 38540 2791 38568
rect 2673 38495 2725 38528
rect 2673 38476 2679 38495
rect 2679 38476 2713 38495
rect 2713 38476 2725 38495
rect 2739 38495 2791 38528
rect 2739 38476 2751 38495
rect 2751 38476 2785 38495
rect 2785 38476 2791 38495
rect 2673 38461 2679 38464
rect 2679 38461 2713 38464
rect 2713 38461 2725 38464
rect 2673 38422 2725 38461
rect 2739 38461 2751 38464
rect 2751 38461 2785 38464
rect 2785 38461 2791 38464
rect 2739 38422 2791 38461
rect 2673 38412 2679 38422
rect 2679 38412 2725 38422
rect 2739 38412 2785 38422
rect 2785 38412 2791 38422
rect 2673 38348 2679 38400
rect 2679 38348 2725 38400
rect 2739 38348 2785 38400
rect 2785 38348 2791 38400
rect 2673 38284 2679 38336
rect 2679 38284 2725 38336
rect 2739 38284 2785 38336
rect 2785 38284 2791 38336
rect 2673 38219 2679 38271
rect 2679 38219 2725 38271
rect 2739 38219 2785 38271
rect 2785 38219 2791 38271
rect 2673 38154 2679 38206
rect 2679 38154 2725 38206
rect 2739 38154 2785 38206
rect 2785 38154 2791 38206
rect 2673 38089 2679 38141
rect 2679 38089 2725 38141
rect 2739 38089 2785 38141
rect 2785 38089 2791 38141
rect 2673 38024 2679 38076
rect 2679 38024 2725 38076
rect 2739 38024 2785 38076
rect 2785 38024 2791 38076
rect 2673 37959 2679 38011
rect 2679 37959 2725 38011
rect 2739 37959 2785 38011
rect 2785 37959 2791 38011
rect 2673 37894 2679 37946
rect 2679 37894 2725 37946
rect 2739 37894 2785 37946
rect 2785 37894 2791 37946
rect 2673 37829 2679 37881
rect 2679 37829 2725 37881
rect 2739 37829 2785 37881
rect 2785 37829 2791 37881
rect 2673 37764 2679 37816
rect 2679 37764 2725 37816
rect 2739 37764 2785 37816
rect 2785 37764 2791 37816
rect 2673 37699 2679 37751
rect 2679 37699 2725 37751
rect 2739 37699 2785 37751
rect 2785 37699 2791 37751
rect 2673 37634 2679 37686
rect 2679 37634 2725 37686
rect 2739 37634 2785 37686
rect 2785 37634 2791 37686
rect 2673 37569 2679 37621
rect 2679 37569 2725 37621
rect 2739 37569 2785 37621
rect 2785 37569 2791 37621
rect 2673 37504 2679 37556
rect 2679 37504 2725 37556
rect 2739 37504 2785 37556
rect 2785 37504 2791 37556
rect 2673 37439 2679 37491
rect 2679 37439 2725 37491
rect 2739 37439 2785 37491
rect 2785 37439 2791 37491
rect 2673 37380 2679 37426
rect 2679 37380 2725 37426
rect 2739 37380 2785 37426
rect 2785 37380 2791 37426
rect 2673 37374 2725 37380
rect 2739 37374 2791 37380
rect 2950 37840 2956 37892
rect 2956 37840 3002 37892
rect 3016 37840 3062 37892
rect 3062 37840 3068 37892
rect 2950 37773 2956 37825
rect 2956 37773 3002 37825
rect 3016 37773 3062 37825
rect 3062 37773 3068 37825
rect 2950 37706 2956 37758
rect 2956 37706 3002 37758
rect 3016 37706 3062 37758
rect 3062 37706 3068 37758
rect 2950 37639 2956 37691
rect 2956 37639 3002 37691
rect 3016 37639 3062 37691
rect 3062 37639 3068 37691
rect 2950 37572 2956 37624
rect 2956 37572 3002 37624
rect 3016 37572 3062 37624
rect 3062 37572 3068 37624
rect 2950 37505 2956 37557
rect 2956 37505 3002 37557
rect 3016 37505 3062 37557
rect 3062 37505 3068 37557
rect 2950 37438 2956 37490
rect 2956 37438 3002 37490
rect 3016 37438 3062 37490
rect 3062 37438 3068 37490
rect 2950 37380 2956 37423
rect 2956 37380 3002 37423
rect 3016 37380 3062 37423
rect 3062 37380 3068 37423
rect 2950 37371 3002 37380
rect 3016 37371 3068 37380
rect 2950 37304 3002 37356
rect 3016 37304 3068 37356
rect 2950 37237 3002 37289
rect 3016 37237 3068 37289
rect 2950 37170 3002 37222
rect 3016 37170 3068 37222
rect 2950 37103 3002 37155
rect 3016 37103 3068 37155
rect 2950 37036 3002 37088
rect 3016 37036 3068 37088
rect 3227 38714 3279 38720
rect 3227 38680 3233 38714
rect 3233 38680 3267 38714
rect 3267 38680 3279 38714
rect 3227 38668 3279 38680
rect 3293 38714 3345 38720
rect 3293 38680 3305 38714
rect 3305 38680 3339 38714
rect 3339 38680 3345 38714
rect 3293 38668 3345 38680
rect 3227 38641 3279 38654
rect 3227 38607 3233 38641
rect 3233 38607 3267 38641
rect 3267 38607 3279 38641
rect 3227 38602 3279 38607
rect 3293 38641 3345 38654
rect 3293 38607 3305 38641
rect 3305 38607 3339 38641
rect 3339 38607 3345 38641
rect 3293 38602 3345 38607
rect 3227 38568 3279 38588
rect 3227 38536 3233 38568
rect 3233 38536 3267 38568
rect 3267 38536 3279 38568
rect 3293 38568 3345 38588
rect 3293 38536 3305 38568
rect 3305 38536 3339 38568
rect 3339 38536 3345 38568
rect 3227 38495 3279 38522
rect 3227 38470 3233 38495
rect 3233 38470 3267 38495
rect 3267 38470 3279 38495
rect 3293 38495 3345 38522
rect 3293 38470 3305 38495
rect 3305 38470 3339 38495
rect 3339 38470 3345 38495
rect 3227 38422 3279 38456
rect 3293 38422 3345 38456
rect 3227 38404 3233 38422
rect 3233 38404 3279 38422
rect 3293 38404 3339 38422
rect 3339 38404 3345 38422
rect 3227 38338 3233 38390
rect 3233 38338 3279 38390
rect 3293 38338 3339 38390
rect 3339 38338 3345 38390
rect 3227 38271 3233 38323
rect 3233 38271 3279 38323
rect 3293 38271 3339 38323
rect 3339 38271 3345 38323
rect 3227 38204 3233 38256
rect 3233 38204 3279 38256
rect 3293 38204 3339 38256
rect 3339 38204 3345 38256
rect 2315 36690 2363 36691
rect 2249 36684 2253 36690
rect 2253 36684 2291 36690
rect 2291 36684 2301 36690
rect 2315 36684 2325 36690
rect 2325 36684 2363 36690
rect 2363 36684 2367 36691
rect 2249 36656 2253 36672
rect 2253 36656 2291 36672
rect 2291 36656 2301 36672
rect 2315 36656 2325 36672
rect 2325 36657 2363 36672
rect 2363 36657 2367 36672
rect 2325 36656 2367 36657
rect 2249 36620 2301 36656
rect 2315 36620 2367 36656
rect 2249 36583 2253 36608
rect 2253 36583 2291 36608
rect 2291 36583 2301 36608
rect 2315 36583 2325 36608
rect 2325 36584 2363 36608
rect 2363 36584 2367 36608
rect 2325 36583 2367 36584
rect 2249 36556 2301 36583
rect 2315 36556 2367 36583
rect 2249 36510 2253 36544
rect 2253 36510 2291 36544
rect 2291 36510 2301 36544
rect 2315 36510 2325 36544
rect 2325 36511 2363 36544
rect 2363 36511 2367 36544
rect 2325 36510 2367 36511
rect 2249 36492 2301 36510
rect 2315 36492 2367 36510
rect 2249 36471 2301 36480
rect 2315 36472 2367 36480
rect 2315 36471 2363 36472
rect 2249 36437 2253 36471
rect 2253 36437 2291 36471
rect 2291 36437 2301 36471
rect 2315 36437 2325 36471
rect 2325 36438 2363 36471
rect 2363 36438 2367 36472
rect 2325 36437 2367 36438
rect 2249 36428 2301 36437
rect 2315 36428 2367 36437
rect 2249 36398 2301 36416
rect 2315 36399 2367 36416
rect 2315 36398 2363 36399
rect 2249 36364 2253 36398
rect 2253 36364 2291 36398
rect 2291 36364 2301 36398
rect 2315 36364 2325 36398
rect 2325 36365 2363 36398
rect 2363 36365 2367 36399
rect 2325 36364 2367 36365
rect 2249 36325 2301 36352
rect 2315 36326 2367 36352
rect 2315 36325 2363 36326
rect 2249 36300 2253 36325
rect 2253 36300 2291 36325
rect 2291 36300 2301 36325
rect 2315 36300 2325 36325
rect 2325 36300 2363 36325
rect 2363 36300 2367 36326
rect 2249 36252 2301 36288
rect 2315 36253 2367 36288
rect 2315 36252 2363 36253
rect 2249 36236 2253 36252
rect 2253 36236 2291 36252
rect 2291 36236 2301 36252
rect 2315 36236 2325 36252
rect 2325 36236 2363 36252
rect 2363 36236 2367 36253
rect 2249 36218 2253 36224
rect 2253 36218 2291 36224
rect 2291 36218 2301 36224
rect 2315 36218 2325 36224
rect 2325 36219 2363 36224
rect 2363 36219 2367 36224
rect 2325 36218 2367 36219
rect 2249 36179 2301 36218
rect 2315 36180 2367 36218
rect 2315 36179 2363 36180
rect 2249 36172 2253 36179
rect 2253 36172 2291 36179
rect 2291 36172 2301 36179
rect 2315 36172 2325 36179
rect 2325 36172 2363 36179
rect 2363 36172 2367 36180
rect 2249 36145 2253 36160
rect 2253 36145 2291 36160
rect 2291 36145 2301 36160
rect 2315 36145 2325 36160
rect 2325 36146 2363 36160
rect 2363 36146 2367 36160
rect 2325 36145 2367 36146
rect 2249 36108 2301 36145
rect 2315 36108 2367 36145
rect 2249 36072 2253 36096
rect 2253 36072 2291 36096
rect 2291 36072 2301 36096
rect 2315 36072 2325 36096
rect 2325 36073 2363 36096
rect 2363 36073 2367 36096
rect 2325 36072 2367 36073
rect 2249 36044 2301 36072
rect 2315 36044 2367 36072
rect 2249 35999 2253 36032
rect 2253 35999 2291 36032
rect 2291 35999 2301 36032
rect 2315 35999 2325 36032
rect 2325 36000 2363 36032
rect 2363 36000 2367 36032
rect 2325 35999 2367 36000
rect 2249 35980 2301 35999
rect 2315 35980 2367 35999
rect 2249 35960 2301 35968
rect 2315 35961 2367 35968
rect 2315 35960 2363 35961
rect 2249 35926 2253 35960
rect 2253 35926 2291 35960
rect 2291 35926 2301 35960
rect 2315 35926 2325 35960
rect 2325 35927 2363 35960
rect 2363 35927 2367 35961
rect 2325 35926 2367 35927
rect 2249 35916 2301 35926
rect 2315 35916 2367 35926
rect 2249 35887 2301 35904
rect 2315 35888 2367 35904
rect 2315 35887 2363 35888
rect 2249 35853 2253 35887
rect 2253 35853 2291 35887
rect 2291 35853 2301 35887
rect 2315 35853 2325 35887
rect 2325 35854 2363 35887
rect 2363 35854 2367 35888
rect 2325 35853 2367 35854
rect 2249 35852 2301 35853
rect 2315 35852 2367 35853
rect 2249 35814 2301 35840
rect 2315 35815 2367 35840
rect 2315 35814 2363 35815
rect 2249 35788 2253 35814
rect 2253 35788 2291 35814
rect 2291 35788 2301 35814
rect 2315 35788 2325 35814
rect 2325 35788 2363 35814
rect 2363 35788 2367 35815
rect 2249 35741 2301 35776
rect 2315 35742 2367 35776
rect 2315 35741 2363 35742
rect 2249 35724 2253 35741
rect 2253 35724 2291 35741
rect 2291 35724 2301 35741
rect 2315 35724 2325 35741
rect 2325 35724 2363 35741
rect 2363 35724 2367 35742
rect 2249 35707 2253 35712
rect 2253 35707 2291 35712
rect 2291 35707 2301 35712
rect 2315 35707 2325 35712
rect 2325 35708 2363 35712
rect 2363 35708 2367 35712
rect 2325 35707 2367 35708
rect 2249 35668 2301 35707
rect 2315 35669 2367 35707
rect 2315 35668 2363 35669
rect 2249 35660 2253 35668
rect 2253 35660 2291 35668
rect 2291 35660 2301 35668
rect 2315 35660 2325 35668
rect 2325 35660 2363 35668
rect 2363 35660 2367 35669
rect 2249 35634 2253 35648
rect 2253 35634 2291 35648
rect 2291 35634 2301 35648
rect 2315 35634 2325 35648
rect 2325 35635 2363 35648
rect 2363 35635 2367 35648
rect 2325 35634 2367 35635
rect 2249 35596 2301 35634
rect 2315 35596 2367 35634
rect 2249 35561 2253 35584
rect 2253 35561 2291 35584
rect 2291 35561 2301 35584
rect 2315 35561 2325 35584
rect 2325 35562 2363 35584
rect 2363 35562 2367 35584
rect 2325 35561 2367 35562
rect 2249 35532 2301 35561
rect 2315 35532 2367 35561
rect 2249 35468 2301 35520
rect 2315 35468 2325 35520
rect 2325 35489 2363 35520
rect 2363 35489 2367 35520
rect 2325 35468 2367 35489
rect 2249 35404 2301 35456
rect 2315 35450 2325 35456
rect 2325 35450 2367 35456
rect 2315 35404 2367 35450
rect 2249 35340 2301 35392
rect 2315 35340 2367 35392
rect 2249 35276 2301 35328
rect 2315 35276 2367 35328
rect 2249 35212 2301 35264
rect 2315 35212 2367 35264
rect 2249 35148 2301 35200
rect 2315 35148 2367 35200
rect 2249 35084 2301 35136
rect 2315 35084 2367 35136
rect 2249 35020 2301 35072
rect 2315 35020 2367 35072
rect 2249 34956 2301 35008
rect 2315 34956 2367 35008
rect 2249 34892 2301 34944
rect 2315 34892 2367 34944
rect 2249 34828 2301 34880
rect 2315 34828 2367 34880
rect 2249 34764 2301 34816
rect 2315 34764 2367 34816
rect 2249 34700 2301 34752
rect 2315 34700 2367 34752
rect 2249 34636 2301 34688
rect 2315 34636 2367 34688
rect 2249 34572 2301 34624
rect 2315 34572 2367 34624
rect 2249 34508 2301 34560
rect 2315 34508 2367 34560
rect 2249 34444 2301 34496
rect 2315 34444 2367 34496
rect 2249 34380 2301 34432
rect 2315 34380 2367 34432
rect 2249 34316 2301 34368
rect 2315 34316 2367 34368
rect 2249 34252 2301 34304
rect 2315 34252 2367 34304
rect 2249 34188 2301 34240
rect 2315 34188 2367 34240
rect 2249 34124 2301 34176
rect 2315 34124 2367 34176
rect 2249 34060 2301 34112
rect 2315 34060 2367 34112
rect 2249 33996 2301 34048
rect 2315 33996 2367 34048
rect 2249 33932 2301 33984
rect 2315 33932 2367 33984
rect 2249 33868 2301 33920
rect 2315 33868 2367 33920
rect 2249 33804 2301 33856
rect 2315 33804 2367 33856
rect 2249 33740 2301 33792
rect 2315 33740 2367 33792
rect 2249 33688 2301 33728
rect 2315 33688 2367 33728
rect 2249 33676 2301 33688
rect 2315 33676 2367 33688
rect 2249 33644 2301 33664
rect 2249 33612 2253 33644
rect 2253 33612 2301 33644
rect 2315 33644 2367 33664
rect 2315 33612 2325 33644
rect 2325 33612 2359 33644
rect 2359 33612 2367 33644
rect 3227 36714 3279 36720
rect 3227 36680 3233 36714
rect 3233 36680 3267 36714
rect 3267 36680 3279 36714
rect 3227 36668 3279 36680
rect 3293 36714 3345 36720
rect 3293 36680 3305 36714
rect 3305 36680 3339 36714
rect 3339 36680 3345 36714
rect 3293 36668 3345 36680
rect 3227 36641 3279 36654
rect 3227 36607 3233 36641
rect 3233 36607 3267 36641
rect 3267 36607 3279 36641
rect 3227 36602 3279 36607
rect 3293 36641 3345 36654
rect 3293 36607 3305 36641
rect 3305 36607 3339 36641
rect 3339 36607 3345 36641
rect 3293 36602 3345 36607
rect 3227 36568 3279 36588
rect 3227 36536 3233 36568
rect 3233 36536 3267 36568
rect 3267 36536 3279 36568
rect 3293 36568 3345 36588
rect 3293 36536 3305 36568
rect 3305 36536 3339 36568
rect 3339 36536 3345 36568
rect 3227 36495 3279 36522
rect 3227 36470 3233 36495
rect 3233 36470 3267 36495
rect 3267 36470 3279 36495
rect 3293 36495 3345 36522
rect 3293 36470 3305 36495
rect 3305 36470 3339 36495
rect 3339 36470 3345 36495
rect 3227 36422 3279 36456
rect 3293 36422 3345 36456
rect 3227 36404 3233 36422
rect 3233 36404 3279 36422
rect 3293 36404 3339 36422
rect 3339 36404 3345 36422
rect 3227 36338 3233 36390
rect 3233 36338 3279 36390
rect 3293 36338 3339 36390
rect 3339 36338 3345 36390
rect 3227 36271 3233 36323
rect 3233 36271 3279 36323
rect 3293 36271 3339 36323
rect 3339 36271 3345 36323
rect 3227 36204 3233 36256
rect 3233 36204 3279 36256
rect 3293 36204 3339 36256
rect 3339 36204 3345 36256
rect 3504 37840 3510 37892
rect 3510 37840 3556 37892
rect 3570 37840 3616 37892
rect 3616 37840 3622 37892
rect 3504 37773 3510 37825
rect 3510 37773 3556 37825
rect 3570 37773 3616 37825
rect 3616 37773 3622 37825
rect 3504 37706 3510 37758
rect 3510 37706 3556 37758
rect 3570 37706 3616 37758
rect 3616 37706 3622 37758
rect 3504 37639 3510 37691
rect 3510 37639 3556 37691
rect 3570 37639 3616 37691
rect 3616 37639 3622 37691
rect 3504 37572 3510 37624
rect 3510 37572 3556 37624
rect 3570 37572 3616 37624
rect 3616 37572 3622 37624
rect 3504 37505 3510 37557
rect 3510 37505 3556 37557
rect 3570 37505 3616 37557
rect 3616 37505 3622 37557
rect 3504 37438 3510 37490
rect 3510 37438 3556 37490
rect 3570 37438 3616 37490
rect 3616 37438 3622 37490
rect 3504 37380 3510 37423
rect 3510 37380 3556 37423
rect 3570 37380 3616 37423
rect 3616 37380 3622 37423
rect 3504 37371 3556 37380
rect 3570 37371 3622 37380
rect 3504 37304 3556 37356
rect 3570 37304 3622 37356
rect 3504 37237 3556 37289
rect 3570 37237 3622 37289
rect 3504 37170 3556 37222
rect 3570 37170 3622 37222
rect 3504 37103 3556 37155
rect 3570 37103 3622 37155
rect 3504 37036 3556 37088
rect 3570 37036 3622 37088
rect 3504 35840 3510 35892
rect 3510 35840 3556 35892
rect 3570 35840 3616 35892
rect 3616 35840 3622 35892
rect 3504 35774 3510 35826
rect 3510 35774 3556 35826
rect 3570 35774 3616 35826
rect 3616 35774 3622 35826
rect 3504 35708 3510 35760
rect 3510 35708 3556 35760
rect 3570 35708 3616 35760
rect 3616 35708 3622 35760
rect 3504 35642 3510 35694
rect 3510 35642 3556 35694
rect 3570 35642 3616 35694
rect 3616 35642 3622 35694
rect 3504 35575 3510 35627
rect 3510 35575 3556 35627
rect 3570 35575 3616 35627
rect 3616 35575 3622 35627
rect 3504 35508 3510 35560
rect 3510 35508 3556 35560
rect 3570 35508 3616 35560
rect 3616 35508 3622 35560
rect 3504 35441 3510 35493
rect 3510 35441 3556 35493
rect 3570 35441 3616 35493
rect 3616 35441 3622 35493
rect 3504 35380 3510 35426
rect 3510 35380 3556 35426
rect 3570 35380 3616 35426
rect 3616 35380 3622 35426
rect 3504 35374 3556 35380
rect 3570 35374 3622 35380
rect 2249 33571 2301 33600
rect 2249 33548 2253 33571
rect 2253 33548 2301 33571
rect 2315 33571 2367 33600
rect 2315 33548 2325 33571
rect 2325 33548 2359 33571
rect 2359 33548 2367 33571
rect 2249 33498 2301 33536
rect 2249 33484 2253 33498
rect 2253 33484 2301 33498
rect 2315 33498 2367 33536
rect 2315 33484 2325 33498
rect 2325 33484 2359 33498
rect 2359 33484 2367 33498
rect 2249 33464 2253 33472
rect 2253 33464 2301 33472
rect 2249 33425 2301 33464
rect 2249 33420 2253 33425
rect 2253 33420 2301 33425
rect 2315 33464 2325 33472
rect 2325 33464 2359 33472
rect 2359 33464 2367 33472
rect 2315 33425 2367 33464
rect 2315 33420 2325 33425
rect 2325 33420 2359 33425
rect 2359 33420 2367 33425
rect 2249 33391 2253 33408
rect 2253 33391 2301 33408
rect 2249 33356 2301 33391
rect 2315 33391 2325 33408
rect 2325 33391 2359 33408
rect 2359 33391 2367 33408
rect 2315 33356 2367 33391
rect 2249 33318 2253 33344
rect 2253 33318 2301 33344
rect 2249 33292 2301 33318
rect 2315 33318 2325 33344
rect 2325 33318 2359 33344
rect 2359 33318 2367 33344
rect 2315 33292 2367 33318
rect 2249 33279 2301 33280
rect 2249 33245 2253 33279
rect 2253 33245 2301 33279
rect 2249 33228 2301 33245
rect 2315 33279 2367 33280
rect 2315 33245 2325 33279
rect 2325 33245 2359 33279
rect 2359 33245 2367 33279
rect 2315 33228 2367 33245
rect 2249 33206 2301 33216
rect 2249 33172 2253 33206
rect 2253 33172 2301 33206
rect 2249 33164 2301 33172
rect 2315 33206 2367 33216
rect 2315 33172 2325 33206
rect 2325 33172 2359 33206
rect 2359 33172 2367 33206
rect 2315 33164 2367 33172
rect 2249 33133 2301 33152
rect 2249 33100 2253 33133
rect 2253 33100 2301 33133
rect 2315 33133 2367 33152
rect 2315 33100 2325 33133
rect 2325 33100 2359 33133
rect 2359 33100 2367 33133
rect 2249 33060 2301 33088
rect 2249 33036 2253 33060
rect 2253 33036 2301 33060
rect 2315 33060 2367 33088
rect 2315 33036 2325 33060
rect 2325 33036 2359 33060
rect 2359 33036 2367 33060
rect 2249 32987 2301 33024
rect 2249 32972 2253 32987
rect 2253 32972 2301 32987
rect 2315 32987 2367 33024
rect 2315 32972 2325 32987
rect 2325 32972 2359 32987
rect 2359 32972 2367 32987
rect 2249 32953 2253 32960
rect 2253 32953 2301 32960
rect 2249 32914 2301 32953
rect 2249 32908 2253 32914
rect 2253 32908 2301 32914
rect 2315 32953 2325 32960
rect 2325 32953 2359 32960
rect 2359 32953 2367 32960
rect 2315 32914 2367 32953
rect 2315 32908 2325 32914
rect 2325 32908 2359 32914
rect 2359 32908 2367 32914
rect 2249 32880 2253 32896
rect 2253 32880 2301 32896
rect 2249 32844 2301 32880
rect 2315 32880 2325 32896
rect 2325 32880 2359 32896
rect 2359 32880 2367 32896
rect 2315 32844 2367 32880
rect 2249 32807 2253 32832
rect 2253 32807 2301 32832
rect 2249 32780 2301 32807
rect 2315 32807 2325 32832
rect 2325 32807 2359 32832
rect 2359 32807 2367 32832
rect 2315 32780 2367 32807
rect 2249 32734 2253 32768
rect 2253 32734 2301 32768
rect 2249 32716 2301 32734
rect 2315 32734 2325 32768
rect 2325 32734 2359 32768
rect 2359 32734 2367 32768
rect 2315 32716 2367 32734
rect 2249 32695 2301 32704
rect 2249 32661 2253 32695
rect 2253 32661 2301 32695
rect 2249 32652 2301 32661
rect 2315 32695 2367 32704
rect 2315 32661 2325 32695
rect 2325 32661 2359 32695
rect 2359 32661 2367 32695
rect 2315 32652 2367 32661
rect 2249 32622 2301 32640
rect 2249 32588 2253 32622
rect 2253 32588 2301 32622
rect 2315 32622 2367 32640
rect 2315 32588 2325 32622
rect 2325 32588 2359 32622
rect 2359 32588 2367 32622
rect 2249 32549 2301 32576
rect 2249 32524 2253 32549
rect 2253 32524 2301 32549
rect 2315 32549 2367 32576
rect 2315 32524 2325 32549
rect 2325 32524 2359 32549
rect 2359 32524 2367 32549
rect 2249 32476 2301 32512
rect 2249 32460 2253 32476
rect 2253 32460 2301 32476
rect 2315 32476 2367 32512
rect 2315 32460 2325 32476
rect 2325 32460 2359 32476
rect 2359 32460 2367 32476
rect 2249 32442 2253 32448
rect 2253 32442 2301 32448
rect 2249 32403 2301 32442
rect 2249 32396 2253 32403
rect 2253 32396 2301 32403
rect 2315 32442 2325 32448
rect 2325 32442 2359 32448
rect 2359 32442 2367 32448
rect 2315 32403 2367 32442
rect 2315 32396 2325 32403
rect 2325 32396 2359 32403
rect 2359 32396 2367 32403
rect 2249 32369 2253 32384
rect 2253 32369 2301 32384
rect 2249 32332 2301 32369
rect 2315 32369 2325 32384
rect 2325 32369 2359 32384
rect 2359 32369 2367 32384
rect 2315 32332 2367 32369
rect 2249 32296 2253 32319
rect 2253 32296 2301 32319
rect 2249 32267 2301 32296
rect 2315 32296 2325 32319
rect 2325 32296 2359 32319
rect 2359 32296 2367 32319
rect 2315 32267 2367 32296
rect 2249 32223 2253 32254
rect 2253 32223 2301 32254
rect 2249 32202 2301 32223
rect 2315 32223 2325 32254
rect 2325 32223 2359 32254
rect 2359 32223 2367 32254
rect 2315 32202 2367 32223
rect 2249 32184 2301 32189
rect 2249 32150 2253 32184
rect 2253 32150 2301 32184
rect 2249 32137 2301 32150
rect 2315 32184 2367 32189
rect 2315 32150 2325 32184
rect 2325 32150 2359 32184
rect 2359 32150 2367 32184
rect 2315 32137 2367 32150
rect 2249 32111 2301 32124
rect 2249 32077 2253 32111
rect 2253 32077 2301 32111
rect 2249 32072 2301 32077
rect 2315 32111 2367 32124
rect 2315 32077 2325 32111
rect 2325 32077 2359 32111
rect 2359 32077 2367 32111
rect 2315 32072 2367 32077
rect 2249 32038 2301 32059
rect 2249 32007 2253 32038
rect 2253 32007 2301 32038
rect 2315 32038 2367 32059
rect 2315 32007 2325 32038
rect 2325 32007 2359 32038
rect 2359 32007 2367 32038
rect 2249 31965 2301 31994
rect 2249 31942 2253 31965
rect 2253 31942 2301 31965
rect 2315 31965 2367 31994
rect 2315 31942 2325 31965
rect 2325 31942 2359 31965
rect 2359 31942 2367 31965
rect 2249 31892 2301 31929
rect 2249 31877 2253 31892
rect 2253 31877 2301 31892
rect 2315 31892 2367 31929
rect 2315 31877 2325 31892
rect 2325 31877 2359 31892
rect 2359 31877 2367 31892
rect 2249 31858 2253 31864
rect 2253 31858 2301 31864
rect 2249 31819 2301 31858
rect 2249 31812 2253 31819
rect 2253 31812 2301 31819
rect 2315 31858 2325 31864
rect 2325 31858 2359 31864
rect 2359 31858 2367 31864
rect 2315 31819 2367 31858
rect 2315 31812 2325 31819
rect 2325 31812 2359 31819
rect 2359 31812 2367 31819
rect 2249 31785 2253 31799
rect 2253 31785 2301 31799
rect 2249 31747 2301 31785
rect 2315 31785 2325 31799
rect 2325 31785 2359 31799
rect 2359 31785 2367 31799
rect 2315 31747 2367 31785
rect 2249 31712 2253 31734
rect 2253 31712 2301 31734
rect 2249 31682 2301 31712
rect 2315 31712 2325 31734
rect 2325 31712 2359 31734
rect 2359 31712 2367 31734
rect 2315 31682 2367 31712
rect 2249 31639 2253 31669
rect 2253 31639 2301 31669
rect 2249 31617 2301 31639
rect 2315 31639 2325 31669
rect 2325 31639 2359 31669
rect 2359 31639 2367 31669
rect 2315 31617 2367 31639
rect 2249 31600 2301 31604
rect 2249 31566 2253 31600
rect 2253 31566 2301 31600
rect 2249 31552 2301 31566
rect 2315 31600 2367 31604
rect 2315 31566 2325 31600
rect 2325 31566 2359 31600
rect 2359 31566 2367 31600
rect 2315 31552 2367 31566
rect 2249 31527 2301 31539
rect 2249 31493 2253 31527
rect 2253 31493 2301 31527
rect 2249 31487 2301 31493
rect 2315 31527 2367 31539
rect 2315 31493 2325 31527
rect 2325 31493 2359 31527
rect 2359 31493 2367 31527
rect 2315 31487 2367 31493
rect 2249 31454 2301 31474
rect 2249 31422 2253 31454
rect 2253 31422 2301 31454
rect 2315 31454 2367 31474
rect 2315 31422 2325 31454
rect 2325 31422 2359 31454
rect 2359 31422 2367 31454
rect 2249 31381 2301 31409
rect 2249 31357 2253 31381
rect 2253 31357 2301 31381
rect 2315 31381 2367 31409
rect 2315 31357 2325 31381
rect 2325 31357 2359 31381
rect 2359 31357 2367 31381
rect 2249 31308 2301 31344
rect 2249 31292 2253 31308
rect 2253 31292 2301 31308
rect 2315 31308 2367 31344
rect 2315 31292 2325 31308
rect 2325 31292 2359 31308
rect 2359 31292 2367 31308
rect 2249 31274 2253 31279
rect 2253 31274 2301 31279
rect 2249 31235 2301 31274
rect 2249 31227 2253 31235
rect 2253 31227 2301 31235
rect 2315 31274 2325 31279
rect 2325 31274 2359 31279
rect 2359 31274 2367 31279
rect 2315 31235 2367 31274
rect 2315 31227 2325 31235
rect 2325 31227 2359 31235
rect 2359 31227 2367 31235
rect 2249 31201 2253 31214
rect 2253 31201 2301 31214
rect 2249 31162 2301 31201
rect 2315 31201 2325 31214
rect 2325 31201 2359 31214
rect 2359 31201 2367 31214
rect 2315 31162 2367 31201
rect 2249 31128 2253 31149
rect 2253 31128 2301 31149
rect 2249 31097 2301 31128
rect 2315 31128 2325 31149
rect 2325 31128 2359 31149
rect 2359 31128 2367 31149
rect 2315 31097 2367 31128
rect 2249 31055 2253 31084
rect 2253 31055 2301 31084
rect 2249 31032 2301 31055
rect 2315 31055 2325 31084
rect 2325 31055 2359 31084
rect 2359 31055 2367 31084
rect 2315 31032 2367 31055
rect 2249 31016 2301 31019
rect 2249 30982 2253 31016
rect 2253 30982 2301 31016
rect 2249 30967 2301 30982
rect 2315 31016 2367 31019
rect 2315 30982 2325 31016
rect 2325 30982 2359 31016
rect 2359 30982 2367 31016
rect 2315 30967 2367 30982
rect 2249 30943 2301 30954
rect 2249 30909 2253 30943
rect 2253 30909 2301 30943
rect 2249 30902 2301 30909
rect 2315 30943 2367 30954
rect 2315 30909 2325 30943
rect 2325 30909 2359 30943
rect 2359 30909 2367 30943
rect 2315 30902 2367 30909
rect 2249 30871 2301 30889
rect 2249 30837 2253 30871
rect 2253 30837 2301 30871
rect 2315 30871 2367 30889
rect 2315 30837 2325 30871
rect 2325 30837 2359 30871
rect 2359 30837 2367 30871
rect 2249 30799 2301 30824
rect 2249 30772 2253 30799
rect 2253 30772 2301 30799
rect 2315 30799 2367 30824
rect 2315 30772 2325 30799
rect 2325 30772 2359 30799
rect 2359 30772 2367 30799
rect 2249 30727 2301 30759
rect 2249 30707 2253 30727
rect 2253 30707 2301 30727
rect 2315 30727 2367 30759
rect 2315 30707 2325 30727
rect 2325 30707 2359 30727
rect 2359 30707 2367 30727
rect 2249 30693 2253 30694
rect 2253 30693 2301 30694
rect 2249 30655 2301 30693
rect 2249 30642 2253 30655
rect 2253 30642 2301 30655
rect 2315 30693 2325 30694
rect 2325 30693 2359 30694
rect 2359 30693 2367 30694
rect 2315 30655 2367 30693
rect 2315 30642 2325 30655
rect 2325 30642 2359 30655
rect 2359 30642 2367 30655
rect 2249 30621 2253 30629
rect 2253 30621 2301 30629
rect 2249 30583 2301 30621
rect 2249 30577 2253 30583
rect 2253 30577 2301 30583
rect 2315 30621 2325 30629
rect 2325 30621 2359 30629
rect 2359 30621 2367 30629
rect 2315 30583 2367 30621
rect 2315 30577 2325 30583
rect 2325 30577 2359 30583
rect 2359 30577 2367 30583
rect 2249 30549 2253 30564
rect 2253 30549 2301 30564
rect 2249 30512 2301 30549
rect 2315 30549 2325 30564
rect 2325 30549 2359 30564
rect 2359 30549 2367 30564
rect 2315 30512 2367 30549
rect 2249 30477 2253 30499
rect 2253 30477 2301 30499
rect 2249 30447 2301 30477
rect 2315 30477 2325 30499
rect 2325 30477 2359 30499
rect 2359 30477 2367 30499
rect 2315 30447 2367 30477
rect 2249 30405 2253 30434
rect 2253 30405 2301 30434
rect 2249 30382 2301 30405
rect 2315 30405 2325 30434
rect 2325 30405 2359 30434
rect 2359 30405 2367 30434
rect 2315 30382 2367 30405
rect 2249 30367 2301 30369
rect 2249 30333 2253 30367
rect 2253 30333 2301 30367
rect 2249 30317 2301 30333
rect 2315 30367 2367 30369
rect 2315 30333 2325 30367
rect 2325 30333 2359 30367
rect 2359 30333 2367 30367
rect 2315 30317 2367 30333
rect 2249 30295 2301 30304
rect 2249 30261 2253 30295
rect 2253 30261 2301 30295
rect 2249 30252 2301 30261
rect 2315 30295 2367 30304
rect 2315 30261 2325 30295
rect 2325 30261 2359 30295
rect 2359 30261 2367 30295
rect 2315 30252 2367 30261
rect 2249 30223 2301 30239
rect 2249 30189 2253 30223
rect 2253 30189 2301 30223
rect 2249 30187 2301 30189
rect 2315 30223 2367 30239
rect 2315 30189 2325 30223
rect 2325 30189 2359 30223
rect 2359 30189 2367 30223
rect 2315 30187 2367 30189
rect 2249 30151 2301 30174
rect 2249 30122 2253 30151
rect 2253 30122 2301 30151
rect 2315 30151 2367 30174
rect 2315 30122 2325 30151
rect 2325 30122 2359 30151
rect 2359 30122 2367 30151
rect 2249 30079 2301 30109
rect 2249 30057 2253 30079
rect 2253 30057 2301 30079
rect 2315 30079 2367 30109
rect 2315 30057 2325 30079
rect 2325 30057 2359 30079
rect 2359 30057 2367 30079
rect 2249 30007 2301 30044
rect 2249 29992 2253 30007
rect 2253 29992 2301 30007
rect 2315 30007 2367 30044
rect 2315 29992 2325 30007
rect 2325 29992 2359 30007
rect 2359 29992 2367 30007
rect 2249 29973 2253 29979
rect 2253 29973 2301 29979
rect 2249 29935 2301 29973
rect 2249 29927 2253 29935
rect 2253 29927 2301 29935
rect 2315 29973 2325 29979
rect 2325 29973 2359 29979
rect 2359 29973 2367 29979
rect 2315 29935 2367 29973
rect 2315 29927 2325 29935
rect 2325 29927 2359 29935
rect 2359 29927 2367 29935
rect 2249 29901 2253 29914
rect 2253 29901 2301 29914
rect 2249 29863 2301 29901
rect 2249 29862 2253 29863
rect 2253 29862 2301 29863
rect 2315 29901 2325 29914
rect 2325 29901 2359 29914
rect 2359 29901 2367 29914
rect 2315 29863 2367 29901
rect 2315 29862 2325 29863
rect 2325 29862 2359 29863
rect 2359 29862 2367 29863
rect 2249 29829 2253 29849
rect 2253 29829 2301 29849
rect 2249 29797 2301 29829
rect 2315 29829 2325 29849
rect 2325 29829 2359 29849
rect 2359 29829 2367 29849
rect 2315 29797 2367 29829
rect 2249 29757 2253 29784
rect 2253 29757 2301 29784
rect 2249 29732 2301 29757
rect 2315 29757 2325 29784
rect 2325 29757 2359 29784
rect 2359 29757 2367 29784
rect 2315 29732 2367 29757
rect 2249 29685 2253 29719
rect 2253 29685 2301 29719
rect 2249 29667 2301 29685
rect 2315 29685 2325 29719
rect 2325 29685 2359 29719
rect 2359 29685 2367 29719
rect 2315 29667 2367 29685
rect 2249 29647 2301 29654
rect 2249 29613 2253 29647
rect 2253 29613 2301 29647
rect 2249 29602 2301 29613
rect 2315 29647 2367 29654
rect 2315 29613 2325 29647
rect 2325 29613 2359 29647
rect 2359 29613 2367 29647
rect 2315 29602 2367 29613
rect 2249 29575 2301 29589
rect 2249 29541 2253 29575
rect 2253 29541 2301 29575
rect 2249 29537 2301 29541
rect 2315 29575 2367 29589
rect 2315 29541 2325 29575
rect 2325 29541 2359 29575
rect 2359 29541 2367 29575
rect 2315 29537 2367 29541
rect 2249 29503 2301 29524
rect 2249 29472 2253 29503
rect 2253 29472 2301 29503
rect 2315 29503 2367 29524
rect 2315 29472 2325 29503
rect 2325 29472 2359 29503
rect 2359 29472 2367 29503
rect 2249 29431 2301 29459
rect 2249 29407 2253 29431
rect 2253 29407 2301 29431
rect 2315 29431 2367 29459
rect 2315 29407 2325 29431
rect 2325 29407 2359 29431
rect 2359 29407 2367 29431
rect 2249 29359 2301 29394
rect 2249 29342 2253 29359
rect 2253 29342 2301 29359
rect 2315 29359 2367 29394
rect 2315 29342 2325 29359
rect 2325 29342 2359 29359
rect 2359 29342 2367 29359
rect 2249 29325 2253 29329
rect 2253 29325 2301 29329
rect 2249 29287 2301 29325
rect 2249 29277 2253 29287
rect 2253 29277 2301 29287
rect 2315 29325 2325 29329
rect 2325 29325 2359 29329
rect 2359 29325 2367 29329
rect 2315 29287 2367 29325
rect 2315 29277 2325 29287
rect 2325 29277 2359 29287
rect 2359 29277 2367 29287
rect 2249 29253 2253 29264
rect 2253 29253 2301 29264
rect 2249 29215 2301 29253
rect 2249 29212 2253 29215
rect 2253 29212 2301 29215
rect 2315 29253 2325 29264
rect 2325 29253 2359 29264
rect 2359 29253 2367 29264
rect 2315 29215 2367 29253
rect 2315 29212 2325 29215
rect 2325 29212 2359 29215
rect 2359 29212 2367 29215
rect 2249 29181 2253 29199
rect 2253 29181 2301 29199
rect 2249 29147 2301 29181
rect 2315 29181 2325 29199
rect 2325 29181 2359 29199
rect 2359 29181 2367 29199
rect 2315 29147 2367 29181
rect 2249 29109 2253 29134
rect 2253 29109 2301 29134
rect 2249 29082 2301 29109
rect 2315 29109 2325 29134
rect 2325 29109 2359 29134
rect 2359 29109 2367 29134
rect 2315 29082 2367 29109
rect 2249 29037 2253 29069
rect 2253 29037 2301 29069
rect 2249 29017 2301 29037
rect 2315 29037 2325 29069
rect 2325 29037 2359 29069
rect 2359 29037 2367 29069
rect 2315 29017 2367 29037
rect 2249 28999 2301 29004
rect 2249 28965 2253 28999
rect 2253 28965 2301 28999
rect 2249 28952 2301 28965
rect 2315 28999 2367 29004
rect 2315 28965 2325 28999
rect 2325 28965 2359 28999
rect 2359 28965 2367 28999
rect 2315 28952 2367 28965
rect 2249 28927 2301 28939
rect 2249 28893 2253 28927
rect 2253 28893 2301 28927
rect 2249 28887 2301 28893
rect 2315 28927 2367 28939
rect 2315 28893 2325 28927
rect 2325 28893 2359 28927
rect 2359 28893 2367 28927
rect 2315 28887 2367 28893
rect 3781 38714 3833 38720
rect 3781 38680 3787 38714
rect 3787 38680 3821 38714
rect 3821 38680 3833 38714
rect 3781 38668 3833 38680
rect 3847 38714 3899 38720
rect 3847 38680 3859 38714
rect 3859 38680 3893 38714
rect 3893 38680 3899 38714
rect 3847 38668 3899 38680
rect 3781 38641 3833 38654
rect 3781 38607 3787 38641
rect 3787 38607 3821 38641
rect 3821 38607 3833 38641
rect 3781 38602 3833 38607
rect 3847 38641 3899 38654
rect 3847 38607 3859 38641
rect 3859 38607 3893 38641
rect 3893 38607 3899 38641
rect 3847 38602 3899 38607
rect 3781 38568 3833 38588
rect 3781 38536 3787 38568
rect 3787 38536 3821 38568
rect 3821 38536 3833 38568
rect 3847 38568 3899 38588
rect 3847 38536 3859 38568
rect 3859 38536 3893 38568
rect 3893 38536 3899 38568
rect 3781 38495 3833 38522
rect 3781 38470 3787 38495
rect 3787 38470 3821 38495
rect 3821 38470 3833 38495
rect 3847 38495 3899 38522
rect 3847 38470 3859 38495
rect 3859 38470 3893 38495
rect 3893 38470 3899 38495
rect 3781 38422 3833 38456
rect 3847 38422 3899 38456
rect 3781 38404 3787 38422
rect 3787 38404 3833 38422
rect 3847 38404 3893 38422
rect 3893 38404 3899 38422
rect 3781 38338 3787 38390
rect 3787 38338 3833 38390
rect 3847 38338 3893 38390
rect 3893 38338 3899 38390
rect 3781 38271 3787 38323
rect 3787 38271 3833 38323
rect 3847 38271 3893 38323
rect 3893 38271 3899 38323
rect 3781 38204 3787 38256
rect 3787 38204 3833 38256
rect 3847 38204 3893 38256
rect 3893 38204 3899 38256
rect 3781 36714 3833 36720
rect 3781 36680 3787 36714
rect 3787 36680 3821 36714
rect 3821 36680 3833 36714
rect 3781 36668 3833 36680
rect 3847 36714 3899 36720
rect 3847 36680 3859 36714
rect 3859 36680 3893 36714
rect 3893 36680 3899 36714
rect 3847 36668 3899 36680
rect 3781 36641 3833 36654
rect 3781 36607 3787 36641
rect 3787 36607 3821 36641
rect 3821 36607 3833 36641
rect 3781 36602 3833 36607
rect 3847 36641 3899 36654
rect 3847 36607 3859 36641
rect 3859 36607 3893 36641
rect 3893 36607 3899 36641
rect 3847 36602 3899 36607
rect 3781 36568 3833 36588
rect 3781 36536 3787 36568
rect 3787 36536 3821 36568
rect 3821 36536 3833 36568
rect 3847 36568 3899 36588
rect 3847 36536 3859 36568
rect 3859 36536 3893 36568
rect 3893 36536 3899 36568
rect 3781 36495 3833 36522
rect 3781 36470 3787 36495
rect 3787 36470 3821 36495
rect 3821 36470 3833 36495
rect 3847 36495 3899 36522
rect 3847 36470 3859 36495
rect 3859 36470 3893 36495
rect 3893 36470 3899 36495
rect 3781 36422 3833 36456
rect 3847 36422 3899 36456
rect 3781 36404 3787 36422
rect 3787 36404 3833 36422
rect 3847 36404 3893 36422
rect 3893 36404 3899 36422
rect 3781 36338 3787 36390
rect 3787 36338 3833 36390
rect 3847 36338 3893 36390
rect 3893 36338 3899 36390
rect 3781 36271 3787 36323
rect 3787 36271 3833 36323
rect 3847 36271 3893 36323
rect 3893 36271 3899 36323
rect 3781 36204 3787 36256
rect 3787 36204 3833 36256
rect 3847 36204 3893 36256
rect 3893 36204 3899 36256
rect 4058 37840 4064 37892
rect 4064 37840 4110 37892
rect 4124 37840 4170 37892
rect 4170 37840 4176 37892
rect 4058 37773 4064 37825
rect 4064 37773 4110 37825
rect 4124 37773 4170 37825
rect 4170 37773 4176 37825
rect 4058 37706 4064 37758
rect 4064 37706 4110 37758
rect 4124 37706 4170 37758
rect 4170 37706 4176 37758
rect 4058 37639 4064 37691
rect 4064 37639 4110 37691
rect 4124 37639 4170 37691
rect 4170 37639 4176 37691
rect 4058 37572 4064 37624
rect 4064 37572 4110 37624
rect 4124 37572 4170 37624
rect 4170 37572 4176 37624
rect 4058 37505 4064 37557
rect 4064 37505 4110 37557
rect 4124 37505 4170 37557
rect 4170 37505 4176 37557
rect 4058 37438 4064 37490
rect 4064 37438 4110 37490
rect 4124 37438 4170 37490
rect 4170 37438 4176 37490
rect 4058 37380 4064 37423
rect 4064 37380 4110 37423
rect 4124 37380 4170 37423
rect 4170 37380 4176 37423
rect 4058 37371 4110 37380
rect 4124 37371 4176 37380
rect 4058 37304 4110 37356
rect 4124 37304 4176 37356
rect 4058 37237 4110 37289
rect 4124 37237 4176 37289
rect 4058 37170 4110 37222
rect 4124 37170 4176 37222
rect 4058 37103 4110 37155
rect 4124 37103 4176 37155
rect 4058 37036 4110 37088
rect 4124 37036 4176 37088
rect 4058 35840 4064 35892
rect 4064 35840 4110 35892
rect 4124 35840 4170 35892
rect 4170 35840 4176 35892
rect 4058 35774 4064 35826
rect 4064 35774 4110 35826
rect 4124 35774 4170 35826
rect 4170 35774 4176 35826
rect 4058 35708 4064 35760
rect 4064 35708 4110 35760
rect 4124 35708 4170 35760
rect 4170 35708 4176 35760
rect 4058 35642 4064 35694
rect 4064 35642 4110 35694
rect 4124 35642 4170 35694
rect 4170 35642 4176 35694
rect 4058 35575 4064 35627
rect 4064 35575 4110 35627
rect 4124 35575 4170 35627
rect 4170 35575 4176 35627
rect 4058 35508 4064 35560
rect 4064 35508 4110 35560
rect 4124 35508 4170 35560
rect 4170 35508 4176 35560
rect 4058 35441 4064 35493
rect 4064 35441 4110 35493
rect 4124 35441 4170 35493
rect 4170 35441 4176 35493
rect 4058 35380 4064 35426
rect 4064 35380 4110 35426
rect 4124 35380 4170 35426
rect 4170 35380 4176 35426
rect 4058 35374 4110 35380
rect 4124 35374 4176 35380
rect 4335 38714 4387 38720
rect 4335 38680 4341 38714
rect 4341 38680 4375 38714
rect 4375 38680 4387 38714
rect 4335 38668 4387 38680
rect 4401 38714 4453 38720
rect 4401 38680 4413 38714
rect 4413 38680 4447 38714
rect 4447 38680 4453 38714
rect 4401 38668 4453 38680
rect 4335 38641 4387 38654
rect 4335 38607 4341 38641
rect 4341 38607 4375 38641
rect 4375 38607 4387 38641
rect 4335 38602 4387 38607
rect 4401 38641 4453 38654
rect 4401 38607 4413 38641
rect 4413 38607 4447 38641
rect 4447 38607 4453 38641
rect 4401 38602 4453 38607
rect 4335 38568 4387 38588
rect 4335 38536 4341 38568
rect 4341 38536 4375 38568
rect 4375 38536 4387 38568
rect 4401 38568 4453 38588
rect 4401 38536 4413 38568
rect 4413 38536 4447 38568
rect 4447 38536 4453 38568
rect 4335 38495 4387 38522
rect 4335 38470 4341 38495
rect 4341 38470 4375 38495
rect 4375 38470 4387 38495
rect 4401 38495 4453 38522
rect 4401 38470 4413 38495
rect 4413 38470 4447 38495
rect 4447 38470 4453 38495
rect 4335 38422 4387 38456
rect 4401 38422 4453 38456
rect 4335 38404 4341 38422
rect 4341 38404 4387 38422
rect 4401 38404 4447 38422
rect 4447 38404 4453 38422
rect 4335 38338 4341 38390
rect 4341 38338 4387 38390
rect 4401 38338 4447 38390
rect 4447 38338 4453 38390
rect 4335 38271 4341 38323
rect 4341 38271 4387 38323
rect 4401 38271 4447 38323
rect 4447 38271 4453 38323
rect 4335 38204 4341 38256
rect 4341 38204 4387 38256
rect 4401 38204 4447 38256
rect 4447 38204 4453 38256
rect 4335 36714 4387 36720
rect 4335 36680 4341 36714
rect 4341 36680 4375 36714
rect 4375 36680 4387 36714
rect 4335 36668 4387 36680
rect 4401 36714 4453 36720
rect 4401 36680 4413 36714
rect 4413 36680 4447 36714
rect 4447 36680 4453 36714
rect 4401 36668 4453 36680
rect 4335 36641 4387 36654
rect 4335 36607 4341 36641
rect 4341 36607 4375 36641
rect 4375 36607 4387 36641
rect 4335 36602 4387 36607
rect 4401 36641 4453 36654
rect 4401 36607 4413 36641
rect 4413 36607 4447 36641
rect 4447 36607 4453 36641
rect 4401 36602 4453 36607
rect 4335 36568 4387 36588
rect 4335 36536 4341 36568
rect 4341 36536 4375 36568
rect 4375 36536 4387 36568
rect 4401 36568 4453 36588
rect 4401 36536 4413 36568
rect 4413 36536 4447 36568
rect 4447 36536 4453 36568
rect 4335 36495 4387 36522
rect 4335 36470 4341 36495
rect 4341 36470 4375 36495
rect 4375 36470 4387 36495
rect 4401 36495 4453 36522
rect 4401 36470 4413 36495
rect 4413 36470 4447 36495
rect 4447 36470 4453 36495
rect 4335 36422 4387 36456
rect 4401 36422 4453 36456
rect 4335 36404 4341 36422
rect 4341 36404 4387 36422
rect 4401 36404 4447 36422
rect 4447 36404 4453 36422
rect 4335 36338 4341 36390
rect 4341 36338 4387 36390
rect 4401 36338 4447 36390
rect 4447 36338 4453 36390
rect 4335 36271 4341 36323
rect 4341 36271 4387 36323
rect 4401 36271 4447 36323
rect 4447 36271 4453 36323
rect 4335 36204 4341 36256
rect 4341 36204 4387 36256
rect 4401 36204 4447 36256
rect 4447 36204 4453 36256
rect 4612 37840 4618 37892
rect 4618 37840 4664 37892
rect 4678 37840 4724 37892
rect 4724 37840 4730 37892
rect 4612 37773 4618 37825
rect 4618 37773 4664 37825
rect 4678 37773 4724 37825
rect 4724 37773 4730 37825
rect 4612 37706 4618 37758
rect 4618 37706 4664 37758
rect 4678 37706 4724 37758
rect 4724 37706 4730 37758
rect 4612 37639 4618 37691
rect 4618 37639 4664 37691
rect 4678 37639 4724 37691
rect 4724 37639 4730 37691
rect 4612 37572 4618 37624
rect 4618 37572 4664 37624
rect 4678 37572 4724 37624
rect 4724 37572 4730 37624
rect 4612 37505 4618 37557
rect 4618 37505 4664 37557
rect 4678 37505 4724 37557
rect 4724 37505 4730 37557
rect 4612 37438 4618 37490
rect 4618 37438 4664 37490
rect 4678 37438 4724 37490
rect 4724 37438 4730 37490
rect 4612 37380 4618 37423
rect 4618 37380 4664 37423
rect 4678 37380 4724 37423
rect 4724 37380 4730 37423
rect 4612 37371 4664 37380
rect 4678 37371 4730 37380
rect 4612 37304 4664 37356
rect 4678 37304 4730 37356
rect 4612 37237 4664 37289
rect 4678 37237 4730 37289
rect 4612 37170 4664 37222
rect 4678 37170 4730 37222
rect 4612 37103 4664 37155
rect 4678 37103 4730 37155
rect 4612 37036 4664 37088
rect 4678 37036 4730 37088
rect 4612 35840 4618 35892
rect 4618 35840 4664 35892
rect 4678 35840 4724 35892
rect 4724 35840 4730 35892
rect 4612 35774 4618 35826
rect 4618 35774 4664 35826
rect 4678 35774 4724 35826
rect 4724 35774 4730 35826
rect 4612 35708 4618 35760
rect 4618 35708 4664 35760
rect 4678 35708 4724 35760
rect 4724 35708 4730 35760
rect 4612 35642 4618 35694
rect 4618 35642 4664 35694
rect 4678 35642 4724 35694
rect 4724 35642 4730 35694
rect 4612 35575 4618 35627
rect 4618 35575 4664 35627
rect 4678 35575 4724 35627
rect 4724 35575 4730 35627
rect 4612 35508 4618 35560
rect 4618 35508 4664 35560
rect 4678 35508 4724 35560
rect 4724 35508 4730 35560
rect 4612 35441 4618 35493
rect 4618 35441 4664 35493
rect 4678 35441 4724 35493
rect 4724 35441 4730 35493
rect 4612 35380 4618 35426
rect 4618 35380 4664 35426
rect 4678 35380 4724 35426
rect 4724 35380 4730 35426
rect 4612 35374 4664 35380
rect 4678 35374 4730 35380
rect 4889 38714 4941 38720
rect 4889 38680 4895 38714
rect 4895 38680 4929 38714
rect 4929 38680 4941 38714
rect 4889 38668 4941 38680
rect 4955 38714 5007 38720
rect 4955 38680 4967 38714
rect 4967 38680 5001 38714
rect 5001 38680 5007 38714
rect 4955 38668 5007 38680
rect 4889 38641 4941 38654
rect 4889 38607 4895 38641
rect 4895 38607 4929 38641
rect 4929 38607 4941 38641
rect 4889 38602 4941 38607
rect 4955 38641 5007 38654
rect 4955 38607 4967 38641
rect 4967 38607 5001 38641
rect 5001 38607 5007 38641
rect 4955 38602 5007 38607
rect 4889 38568 4941 38588
rect 4889 38536 4895 38568
rect 4895 38536 4929 38568
rect 4929 38536 4941 38568
rect 4955 38568 5007 38588
rect 4955 38536 4967 38568
rect 4967 38536 5001 38568
rect 5001 38536 5007 38568
rect 4889 38495 4941 38522
rect 4889 38470 4895 38495
rect 4895 38470 4929 38495
rect 4929 38470 4941 38495
rect 4955 38495 5007 38522
rect 4955 38470 4967 38495
rect 4967 38470 5001 38495
rect 5001 38470 5007 38495
rect 4889 38422 4941 38456
rect 4955 38422 5007 38456
rect 4889 38404 4895 38422
rect 4895 38404 4941 38422
rect 4955 38404 5001 38422
rect 5001 38404 5007 38422
rect 4889 38338 4895 38390
rect 4895 38338 4941 38390
rect 4955 38338 5001 38390
rect 5001 38338 5007 38390
rect 4889 38271 4895 38323
rect 4895 38271 4941 38323
rect 4955 38271 5001 38323
rect 5001 38271 5007 38323
rect 4889 38204 4895 38256
rect 4895 38204 4941 38256
rect 4955 38204 5001 38256
rect 5001 38204 5007 38256
rect 4889 36714 4941 36720
rect 4889 36680 4895 36714
rect 4895 36680 4929 36714
rect 4929 36680 4941 36714
rect 4889 36668 4941 36680
rect 4955 36714 5007 36720
rect 4955 36680 4967 36714
rect 4967 36680 5001 36714
rect 5001 36680 5007 36714
rect 4955 36668 5007 36680
rect 4889 36641 4941 36654
rect 4889 36607 4895 36641
rect 4895 36607 4929 36641
rect 4929 36607 4941 36641
rect 4889 36602 4941 36607
rect 4955 36641 5007 36654
rect 4955 36607 4967 36641
rect 4967 36607 5001 36641
rect 5001 36607 5007 36641
rect 4955 36602 5007 36607
rect 4889 36568 4941 36588
rect 4889 36536 4895 36568
rect 4895 36536 4929 36568
rect 4929 36536 4941 36568
rect 4955 36568 5007 36588
rect 4955 36536 4967 36568
rect 4967 36536 5001 36568
rect 5001 36536 5007 36568
rect 4889 36495 4941 36522
rect 4889 36470 4895 36495
rect 4895 36470 4929 36495
rect 4929 36470 4941 36495
rect 4955 36495 5007 36522
rect 4955 36470 4967 36495
rect 4967 36470 5001 36495
rect 5001 36470 5007 36495
rect 4889 36422 4941 36456
rect 4955 36422 5007 36456
rect 4889 36404 4895 36422
rect 4895 36404 4941 36422
rect 4955 36404 5001 36422
rect 5001 36404 5007 36422
rect 4889 36338 4895 36390
rect 4895 36338 4941 36390
rect 4955 36338 5001 36390
rect 5001 36338 5007 36390
rect 4889 36271 4895 36323
rect 4895 36271 4941 36323
rect 4955 36271 5001 36323
rect 5001 36271 5007 36323
rect 4889 36204 4895 36256
rect 4895 36204 4941 36256
rect 4955 36204 5001 36256
rect 5001 36204 5007 36256
rect 5166 37840 5172 37892
rect 5172 37840 5218 37892
rect 5232 37840 5278 37892
rect 5278 37840 5284 37892
rect 5166 37773 5172 37825
rect 5172 37773 5218 37825
rect 5232 37773 5278 37825
rect 5278 37773 5284 37825
rect 5166 37706 5172 37758
rect 5172 37706 5218 37758
rect 5232 37706 5278 37758
rect 5278 37706 5284 37758
rect 5166 37639 5172 37691
rect 5172 37639 5218 37691
rect 5232 37639 5278 37691
rect 5278 37639 5284 37691
rect 5166 37572 5172 37624
rect 5172 37572 5218 37624
rect 5232 37572 5278 37624
rect 5278 37572 5284 37624
rect 5166 37505 5172 37557
rect 5172 37505 5218 37557
rect 5232 37505 5278 37557
rect 5278 37505 5284 37557
rect 5166 37438 5172 37490
rect 5172 37438 5218 37490
rect 5232 37438 5278 37490
rect 5278 37438 5284 37490
rect 5166 37380 5172 37423
rect 5172 37380 5218 37423
rect 5232 37380 5278 37423
rect 5278 37380 5284 37423
rect 5166 37371 5218 37380
rect 5232 37371 5284 37380
rect 5166 37304 5218 37356
rect 5232 37304 5284 37356
rect 5166 37237 5218 37289
rect 5232 37237 5284 37289
rect 5166 37170 5218 37222
rect 5232 37170 5284 37222
rect 5166 37103 5218 37155
rect 5232 37103 5284 37155
rect 5166 37036 5218 37088
rect 5232 37036 5284 37088
rect 5166 35840 5172 35892
rect 5172 35840 5218 35892
rect 5232 35840 5278 35892
rect 5278 35840 5284 35892
rect 5166 35774 5172 35826
rect 5172 35774 5218 35826
rect 5232 35774 5278 35826
rect 5278 35774 5284 35826
rect 5166 35708 5172 35760
rect 5172 35708 5218 35760
rect 5232 35708 5278 35760
rect 5278 35708 5284 35760
rect 5166 35642 5172 35694
rect 5172 35642 5218 35694
rect 5232 35642 5278 35694
rect 5278 35642 5284 35694
rect 5166 35575 5172 35627
rect 5172 35575 5218 35627
rect 5232 35575 5278 35627
rect 5278 35575 5284 35627
rect 5166 35508 5172 35560
rect 5172 35508 5218 35560
rect 5232 35508 5278 35560
rect 5278 35508 5284 35560
rect 5166 35441 5172 35493
rect 5172 35441 5218 35493
rect 5232 35441 5278 35493
rect 5278 35441 5284 35493
rect 5166 35380 5172 35426
rect 5172 35380 5218 35426
rect 5232 35380 5278 35426
rect 5278 35380 5284 35426
rect 5166 35374 5218 35380
rect 5232 35374 5284 35380
rect 5443 38714 5495 38720
rect 5443 38680 5449 38714
rect 5449 38680 5483 38714
rect 5483 38680 5495 38714
rect 5443 38668 5495 38680
rect 5509 38714 5561 38720
rect 5509 38680 5521 38714
rect 5521 38680 5555 38714
rect 5555 38680 5561 38714
rect 5509 38668 5561 38680
rect 5443 38641 5495 38654
rect 5443 38607 5449 38641
rect 5449 38607 5483 38641
rect 5483 38607 5495 38641
rect 5443 38602 5495 38607
rect 5509 38641 5561 38654
rect 5509 38607 5521 38641
rect 5521 38607 5555 38641
rect 5555 38607 5561 38641
rect 5509 38602 5561 38607
rect 5443 38568 5495 38588
rect 5443 38536 5449 38568
rect 5449 38536 5483 38568
rect 5483 38536 5495 38568
rect 5509 38568 5561 38588
rect 5509 38536 5521 38568
rect 5521 38536 5555 38568
rect 5555 38536 5561 38568
rect 5443 38495 5495 38522
rect 5443 38470 5449 38495
rect 5449 38470 5483 38495
rect 5483 38470 5495 38495
rect 5509 38495 5561 38522
rect 5509 38470 5521 38495
rect 5521 38470 5555 38495
rect 5555 38470 5561 38495
rect 5443 38422 5495 38456
rect 5509 38422 5561 38456
rect 5443 38404 5449 38422
rect 5449 38404 5495 38422
rect 5509 38404 5555 38422
rect 5555 38404 5561 38422
rect 5443 38338 5449 38390
rect 5449 38338 5495 38390
rect 5509 38338 5555 38390
rect 5555 38338 5561 38390
rect 5443 38271 5449 38323
rect 5449 38271 5495 38323
rect 5509 38271 5555 38323
rect 5555 38271 5561 38323
rect 5443 38204 5449 38256
rect 5449 38204 5495 38256
rect 5509 38204 5555 38256
rect 5555 38204 5561 38256
rect 5443 36714 5495 36720
rect 5443 36680 5449 36714
rect 5449 36680 5483 36714
rect 5483 36680 5495 36714
rect 5443 36668 5495 36680
rect 5509 36714 5561 36720
rect 5509 36680 5521 36714
rect 5521 36680 5555 36714
rect 5555 36680 5561 36714
rect 5509 36668 5561 36680
rect 5443 36641 5495 36654
rect 5443 36607 5449 36641
rect 5449 36607 5483 36641
rect 5483 36607 5495 36641
rect 5443 36602 5495 36607
rect 5509 36641 5561 36654
rect 5509 36607 5521 36641
rect 5521 36607 5555 36641
rect 5555 36607 5561 36641
rect 5509 36602 5561 36607
rect 5443 36568 5495 36588
rect 5443 36536 5449 36568
rect 5449 36536 5483 36568
rect 5483 36536 5495 36568
rect 5509 36568 5561 36588
rect 5509 36536 5521 36568
rect 5521 36536 5555 36568
rect 5555 36536 5561 36568
rect 5443 36495 5495 36522
rect 5443 36470 5449 36495
rect 5449 36470 5483 36495
rect 5483 36470 5495 36495
rect 5509 36495 5561 36522
rect 5509 36470 5521 36495
rect 5521 36470 5555 36495
rect 5555 36470 5561 36495
rect 5443 36422 5495 36456
rect 5509 36422 5561 36456
rect 5443 36404 5449 36422
rect 5449 36404 5495 36422
rect 5509 36404 5555 36422
rect 5555 36404 5561 36422
rect 5443 36338 5449 36390
rect 5449 36338 5495 36390
rect 5509 36338 5555 36390
rect 5555 36338 5561 36390
rect 5443 36271 5449 36323
rect 5449 36271 5495 36323
rect 5509 36271 5555 36323
rect 5555 36271 5561 36323
rect 5443 36204 5449 36256
rect 5449 36204 5495 36256
rect 5509 36204 5555 36256
rect 5555 36204 5561 36256
rect 5720 37840 5726 37892
rect 5726 37840 5772 37892
rect 5786 37840 5832 37892
rect 5832 37840 5838 37892
rect 5720 37773 5726 37825
rect 5726 37773 5772 37825
rect 5786 37773 5832 37825
rect 5832 37773 5838 37825
rect 5720 37706 5726 37758
rect 5726 37706 5772 37758
rect 5786 37706 5832 37758
rect 5832 37706 5838 37758
rect 5720 37639 5726 37691
rect 5726 37639 5772 37691
rect 5786 37639 5832 37691
rect 5832 37639 5838 37691
rect 5720 37572 5726 37624
rect 5726 37572 5772 37624
rect 5786 37572 5832 37624
rect 5832 37572 5838 37624
rect 5720 37505 5726 37557
rect 5726 37505 5772 37557
rect 5786 37505 5832 37557
rect 5832 37505 5838 37557
rect 5720 37438 5726 37490
rect 5726 37438 5772 37490
rect 5786 37438 5832 37490
rect 5832 37438 5838 37490
rect 5720 37380 5726 37423
rect 5726 37380 5772 37423
rect 5786 37380 5832 37423
rect 5832 37380 5838 37423
rect 5720 37371 5772 37380
rect 5786 37371 5838 37380
rect 5720 37304 5772 37356
rect 5786 37304 5838 37356
rect 5720 37237 5772 37289
rect 5786 37237 5838 37289
rect 5720 37170 5772 37222
rect 5786 37170 5838 37222
rect 5720 37103 5772 37155
rect 5786 37103 5838 37155
rect 5720 37036 5772 37088
rect 5786 37036 5838 37088
rect 5720 35840 5726 35892
rect 5726 35840 5772 35892
rect 5786 35840 5832 35892
rect 5832 35840 5838 35892
rect 5720 35774 5726 35826
rect 5726 35774 5772 35826
rect 5786 35774 5832 35826
rect 5832 35774 5838 35826
rect 5720 35708 5726 35760
rect 5726 35708 5772 35760
rect 5786 35708 5832 35760
rect 5832 35708 5838 35760
rect 5720 35642 5726 35694
rect 5726 35642 5772 35694
rect 5786 35642 5832 35694
rect 5832 35642 5838 35694
rect 5720 35575 5726 35627
rect 5726 35575 5772 35627
rect 5786 35575 5832 35627
rect 5832 35575 5838 35627
rect 5720 35508 5726 35560
rect 5726 35508 5772 35560
rect 5786 35508 5832 35560
rect 5832 35508 5838 35560
rect 5720 35441 5726 35493
rect 5726 35441 5772 35493
rect 5786 35441 5832 35493
rect 5832 35441 5838 35493
rect 5720 35380 5726 35426
rect 5726 35380 5772 35426
rect 5786 35380 5832 35426
rect 5832 35380 5838 35426
rect 5720 35374 5772 35380
rect 5786 35374 5838 35380
rect 5997 38714 6049 38720
rect 5997 38680 6003 38714
rect 6003 38680 6037 38714
rect 6037 38680 6049 38714
rect 5997 38668 6049 38680
rect 6063 38714 6115 38720
rect 6063 38680 6075 38714
rect 6075 38680 6109 38714
rect 6109 38680 6115 38714
rect 6063 38668 6115 38680
rect 5997 38641 6049 38654
rect 5997 38607 6003 38641
rect 6003 38607 6037 38641
rect 6037 38607 6049 38641
rect 5997 38602 6049 38607
rect 6063 38641 6115 38654
rect 6063 38607 6075 38641
rect 6075 38607 6109 38641
rect 6109 38607 6115 38641
rect 6063 38602 6115 38607
rect 5997 38568 6049 38588
rect 5997 38536 6003 38568
rect 6003 38536 6037 38568
rect 6037 38536 6049 38568
rect 6063 38568 6115 38588
rect 6063 38536 6075 38568
rect 6075 38536 6109 38568
rect 6109 38536 6115 38568
rect 5997 38495 6049 38522
rect 5997 38470 6003 38495
rect 6003 38470 6037 38495
rect 6037 38470 6049 38495
rect 6063 38495 6115 38522
rect 6063 38470 6075 38495
rect 6075 38470 6109 38495
rect 6109 38470 6115 38495
rect 5997 38422 6049 38456
rect 6063 38422 6115 38456
rect 5997 38404 6003 38422
rect 6003 38404 6049 38422
rect 6063 38404 6109 38422
rect 6109 38404 6115 38422
rect 5997 38338 6003 38390
rect 6003 38338 6049 38390
rect 6063 38338 6109 38390
rect 6109 38338 6115 38390
rect 5997 38271 6003 38323
rect 6003 38271 6049 38323
rect 6063 38271 6109 38323
rect 6109 38271 6115 38323
rect 5997 38204 6003 38256
rect 6003 38204 6049 38256
rect 6063 38204 6109 38256
rect 6109 38204 6115 38256
rect 5997 36714 6049 36720
rect 5997 36680 6003 36714
rect 6003 36680 6037 36714
rect 6037 36680 6049 36714
rect 5997 36668 6049 36680
rect 6063 36714 6115 36720
rect 6063 36680 6075 36714
rect 6075 36680 6109 36714
rect 6109 36680 6115 36714
rect 6063 36668 6115 36680
rect 5997 36641 6049 36654
rect 5997 36607 6003 36641
rect 6003 36607 6037 36641
rect 6037 36607 6049 36641
rect 5997 36602 6049 36607
rect 6063 36641 6115 36654
rect 6063 36607 6075 36641
rect 6075 36607 6109 36641
rect 6109 36607 6115 36641
rect 6063 36602 6115 36607
rect 5997 36568 6049 36588
rect 5997 36536 6003 36568
rect 6003 36536 6037 36568
rect 6037 36536 6049 36568
rect 6063 36568 6115 36588
rect 6063 36536 6075 36568
rect 6075 36536 6109 36568
rect 6109 36536 6115 36568
rect 5997 36495 6049 36522
rect 5997 36470 6003 36495
rect 6003 36470 6037 36495
rect 6037 36470 6049 36495
rect 6063 36495 6115 36522
rect 6063 36470 6075 36495
rect 6075 36470 6109 36495
rect 6109 36470 6115 36495
rect 5997 36422 6049 36456
rect 6063 36422 6115 36456
rect 5997 36404 6003 36422
rect 6003 36404 6049 36422
rect 6063 36404 6109 36422
rect 6109 36404 6115 36422
rect 5997 36338 6003 36390
rect 6003 36338 6049 36390
rect 6063 36338 6109 36390
rect 6109 36338 6115 36390
rect 5997 36271 6003 36323
rect 6003 36271 6049 36323
rect 6063 36271 6109 36323
rect 6109 36271 6115 36323
rect 5997 36204 6003 36256
rect 6003 36204 6049 36256
rect 6063 36204 6109 36256
rect 6109 36204 6115 36256
rect 6274 37840 6280 37892
rect 6280 37840 6326 37892
rect 6340 37840 6386 37892
rect 6386 37840 6392 37892
rect 6274 37773 6280 37825
rect 6280 37773 6326 37825
rect 6340 37773 6386 37825
rect 6386 37773 6392 37825
rect 6274 37706 6280 37758
rect 6280 37706 6326 37758
rect 6340 37706 6386 37758
rect 6386 37706 6392 37758
rect 6274 37639 6280 37691
rect 6280 37639 6326 37691
rect 6340 37639 6386 37691
rect 6386 37639 6392 37691
rect 6274 37572 6280 37624
rect 6280 37572 6326 37624
rect 6340 37572 6386 37624
rect 6386 37572 6392 37624
rect 6274 37505 6280 37557
rect 6280 37505 6326 37557
rect 6340 37505 6386 37557
rect 6386 37505 6392 37557
rect 6274 37438 6280 37490
rect 6280 37438 6326 37490
rect 6340 37438 6386 37490
rect 6386 37438 6392 37490
rect 6274 37380 6280 37423
rect 6280 37380 6326 37423
rect 6340 37380 6386 37423
rect 6386 37380 6392 37423
rect 6274 37371 6326 37380
rect 6340 37371 6392 37380
rect 6274 37304 6326 37356
rect 6340 37304 6392 37356
rect 6274 37237 6326 37289
rect 6340 37237 6392 37289
rect 6274 37170 6326 37222
rect 6340 37170 6392 37222
rect 6274 37103 6326 37155
rect 6340 37103 6392 37155
rect 6274 37036 6326 37088
rect 6340 37036 6392 37088
rect 6274 35840 6280 35892
rect 6280 35840 6326 35892
rect 6340 35840 6386 35892
rect 6386 35840 6392 35892
rect 6274 35774 6280 35826
rect 6280 35774 6326 35826
rect 6340 35774 6386 35826
rect 6386 35774 6392 35826
rect 6274 35708 6280 35760
rect 6280 35708 6326 35760
rect 6340 35708 6386 35760
rect 6386 35708 6392 35760
rect 6274 35642 6280 35694
rect 6280 35642 6326 35694
rect 6340 35642 6386 35694
rect 6386 35642 6392 35694
rect 6274 35575 6280 35627
rect 6280 35575 6326 35627
rect 6340 35575 6386 35627
rect 6386 35575 6392 35627
rect 6274 35508 6280 35560
rect 6280 35508 6326 35560
rect 6340 35508 6386 35560
rect 6386 35508 6392 35560
rect 6274 35441 6280 35493
rect 6280 35441 6326 35493
rect 6340 35441 6386 35493
rect 6386 35441 6392 35493
rect 6274 35380 6280 35426
rect 6280 35380 6326 35426
rect 6340 35380 6386 35426
rect 6386 35380 6392 35426
rect 6274 35374 6326 35380
rect 6340 35374 6392 35380
rect 6551 38714 6603 38720
rect 6551 38680 6557 38714
rect 6557 38680 6591 38714
rect 6591 38680 6603 38714
rect 6551 38668 6603 38680
rect 6617 38714 6669 38720
rect 6617 38680 6629 38714
rect 6629 38680 6663 38714
rect 6663 38680 6669 38714
rect 6617 38668 6669 38680
rect 6551 38641 6603 38654
rect 6551 38607 6557 38641
rect 6557 38607 6591 38641
rect 6591 38607 6603 38641
rect 6551 38602 6603 38607
rect 6617 38641 6669 38654
rect 6617 38607 6629 38641
rect 6629 38607 6663 38641
rect 6663 38607 6669 38641
rect 6617 38602 6669 38607
rect 6551 38568 6603 38588
rect 6551 38536 6557 38568
rect 6557 38536 6591 38568
rect 6591 38536 6603 38568
rect 6617 38568 6669 38588
rect 6617 38536 6629 38568
rect 6629 38536 6663 38568
rect 6663 38536 6669 38568
rect 6551 38495 6603 38522
rect 6551 38470 6557 38495
rect 6557 38470 6591 38495
rect 6591 38470 6603 38495
rect 6617 38495 6669 38522
rect 6617 38470 6629 38495
rect 6629 38470 6663 38495
rect 6663 38470 6669 38495
rect 6551 38422 6603 38456
rect 6617 38422 6669 38456
rect 6551 38404 6557 38422
rect 6557 38404 6603 38422
rect 6617 38404 6663 38422
rect 6663 38404 6669 38422
rect 6551 38338 6557 38390
rect 6557 38338 6603 38390
rect 6617 38338 6663 38390
rect 6663 38338 6669 38390
rect 6551 38271 6557 38323
rect 6557 38271 6603 38323
rect 6617 38271 6663 38323
rect 6663 38271 6669 38323
rect 6551 38204 6557 38256
rect 6557 38204 6603 38256
rect 6617 38204 6663 38256
rect 6663 38204 6669 38256
rect 6551 36714 6603 36720
rect 6551 36680 6557 36714
rect 6557 36680 6591 36714
rect 6591 36680 6603 36714
rect 6551 36668 6603 36680
rect 6617 36714 6669 36720
rect 6617 36680 6629 36714
rect 6629 36680 6663 36714
rect 6663 36680 6669 36714
rect 6617 36668 6669 36680
rect 6551 36641 6603 36654
rect 6551 36607 6557 36641
rect 6557 36607 6591 36641
rect 6591 36607 6603 36641
rect 6551 36602 6603 36607
rect 6617 36641 6669 36654
rect 6617 36607 6629 36641
rect 6629 36607 6663 36641
rect 6663 36607 6669 36641
rect 6617 36602 6669 36607
rect 6551 36568 6603 36588
rect 6551 36536 6557 36568
rect 6557 36536 6591 36568
rect 6591 36536 6603 36568
rect 6617 36568 6669 36588
rect 6617 36536 6629 36568
rect 6629 36536 6663 36568
rect 6663 36536 6669 36568
rect 6551 36495 6603 36522
rect 6551 36470 6557 36495
rect 6557 36470 6591 36495
rect 6591 36470 6603 36495
rect 6617 36495 6669 36522
rect 6617 36470 6629 36495
rect 6629 36470 6663 36495
rect 6663 36470 6669 36495
rect 6551 36422 6603 36456
rect 6617 36422 6669 36456
rect 6551 36404 6557 36422
rect 6557 36404 6603 36422
rect 6617 36404 6663 36422
rect 6663 36404 6669 36422
rect 6551 36338 6557 36390
rect 6557 36338 6603 36390
rect 6617 36338 6663 36390
rect 6663 36338 6669 36390
rect 6551 36271 6557 36323
rect 6557 36271 6603 36323
rect 6617 36271 6663 36323
rect 6663 36271 6669 36323
rect 6551 36204 6557 36256
rect 6557 36204 6603 36256
rect 6617 36204 6663 36256
rect 6663 36204 6669 36256
rect 6828 37840 6834 37892
rect 6834 37840 6880 37892
rect 6894 37840 6940 37892
rect 6940 37840 6946 37892
rect 6828 37773 6834 37825
rect 6834 37773 6880 37825
rect 6894 37773 6940 37825
rect 6940 37773 6946 37825
rect 6828 37706 6834 37758
rect 6834 37706 6880 37758
rect 6894 37706 6940 37758
rect 6940 37706 6946 37758
rect 6828 37639 6834 37691
rect 6834 37639 6880 37691
rect 6894 37639 6940 37691
rect 6940 37639 6946 37691
rect 6828 37572 6834 37624
rect 6834 37572 6880 37624
rect 6894 37572 6940 37624
rect 6940 37572 6946 37624
rect 6828 37505 6834 37557
rect 6834 37505 6880 37557
rect 6894 37505 6940 37557
rect 6940 37505 6946 37557
rect 6828 37438 6834 37490
rect 6834 37438 6880 37490
rect 6894 37438 6940 37490
rect 6940 37438 6946 37490
rect 6828 37380 6834 37423
rect 6834 37380 6880 37423
rect 6894 37380 6940 37423
rect 6940 37380 6946 37423
rect 6828 37371 6880 37380
rect 6894 37371 6946 37380
rect 6828 37304 6880 37356
rect 6894 37304 6946 37356
rect 6828 37237 6880 37289
rect 6894 37237 6946 37289
rect 6828 37170 6880 37222
rect 6894 37170 6946 37222
rect 6828 37103 6880 37155
rect 6894 37103 6946 37155
rect 6828 37036 6880 37088
rect 6894 37036 6946 37088
rect 6828 35840 6834 35892
rect 6834 35840 6880 35892
rect 6894 35840 6940 35892
rect 6940 35840 6946 35892
rect 6828 35774 6834 35826
rect 6834 35774 6880 35826
rect 6894 35774 6940 35826
rect 6940 35774 6946 35826
rect 6828 35708 6834 35760
rect 6834 35708 6880 35760
rect 6894 35708 6940 35760
rect 6940 35708 6946 35760
rect 6828 35642 6834 35694
rect 6834 35642 6880 35694
rect 6894 35642 6940 35694
rect 6940 35642 6946 35694
rect 6828 35575 6834 35627
rect 6834 35575 6880 35627
rect 6894 35575 6940 35627
rect 6940 35575 6946 35627
rect 6828 35508 6834 35560
rect 6834 35508 6880 35560
rect 6894 35508 6940 35560
rect 6940 35508 6946 35560
rect 6828 35441 6834 35493
rect 6834 35441 6880 35493
rect 6894 35441 6940 35493
rect 6940 35441 6946 35493
rect 6828 35380 6834 35426
rect 6834 35380 6880 35426
rect 6894 35380 6940 35426
rect 6940 35380 6946 35426
rect 6828 35374 6880 35380
rect 6894 35374 6946 35380
rect 7105 38714 7157 38720
rect 7105 38680 7111 38714
rect 7111 38680 7145 38714
rect 7145 38680 7157 38714
rect 7105 38668 7157 38680
rect 7171 38714 7223 38720
rect 7171 38680 7183 38714
rect 7183 38680 7217 38714
rect 7217 38680 7223 38714
rect 7171 38668 7223 38680
rect 7105 38641 7157 38654
rect 7105 38607 7111 38641
rect 7111 38607 7145 38641
rect 7145 38607 7157 38641
rect 7105 38602 7157 38607
rect 7171 38641 7223 38654
rect 7171 38607 7183 38641
rect 7183 38607 7217 38641
rect 7217 38607 7223 38641
rect 7171 38602 7223 38607
rect 7105 38568 7157 38588
rect 7105 38536 7111 38568
rect 7111 38536 7145 38568
rect 7145 38536 7157 38568
rect 7171 38568 7223 38588
rect 7171 38536 7183 38568
rect 7183 38536 7217 38568
rect 7217 38536 7223 38568
rect 7105 38495 7157 38522
rect 7105 38470 7111 38495
rect 7111 38470 7145 38495
rect 7145 38470 7157 38495
rect 7171 38495 7223 38522
rect 7171 38470 7183 38495
rect 7183 38470 7217 38495
rect 7217 38470 7223 38495
rect 7105 38422 7157 38456
rect 7171 38422 7223 38456
rect 7105 38404 7111 38422
rect 7111 38404 7157 38422
rect 7171 38404 7217 38422
rect 7217 38404 7223 38422
rect 7105 38338 7111 38390
rect 7111 38338 7157 38390
rect 7171 38338 7217 38390
rect 7217 38338 7223 38390
rect 7105 38271 7111 38323
rect 7111 38271 7157 38323
rect 7171 38271 7217 38323
rect 7217 38271 7223 38323
rect 7105 38204 7111 38256
rect 7111 38204 7157 38256
rect 7171 38204 7217 38256
rect 7217 38204 7223 38256
rect 7105 36714 7157 36720
rect 7105 36680 7111 36714
rect 7111 36680 7145 36714
rect 7145 36680 7157 36714
rect 7105 36668 7157 36680
rect 7171 36714 7223 36720
rect 7171 36680 7183 36714
rect 7183 36680 7217 36714
rect 7217 36680 7223 36714
rect 7171 36668 7223 36680
rect 7105 36641 7157 36654
rect 7105 36607 7111 36641
rect 7111 36607 7145 36641
rect 7145 36607 7157 36641
rect 7105 36602 7157 36607
rect 7171 36641 7223 36654
rect 7171 36607 7183 36641
rect 7183 36607 7217 36641
rect 7217 36607 7223 36641
rect 7171 36602 7223 36607
rect 7105 36568 7157 36588
rect 7105 36536 7111 36568
rect 7111 36536 7145 36568
rect 7145 36536 7157 36568
rect 7171 36568 7223 36588
rect 7171 36536 7183 36568
rect 7183 36536 7217 36568
rect 7217 36536 7223 36568
rect 7105 36495 7157 36522
rect 7105 36470 7111 36495
rect 7111 36470 7145 36495
rect 7145 36470 7157 36495
rect 7171 36495 7223 36522
rect 7171 36470 7183 36495
rect 7183 36470 7217 36495
rect 7217 36470 7223 36495
rect 7105 36422 7157 36456
rect 7171 36422 7223 36456
rect 7105 36404 7111 36422
rect 7111 36404 7157 36422
rect 7171 36404 7217 36422
rect 7217 36404 7223 36422
rect 7105 36338 7111 36390
rect 7111 36338 7157 36390
rect 7171 36338 7217 36390
rect 7217 36338 7223 36390
rect 7105 36271 7111 36323
rect 7111 36271 7157 36323
rect 7171 36271 7217 36323
rect 7217 36271 7223 36323
rect 7105 36204 7111 36256
rect 7111 36204 7157 36256
rect 7171 36204 7217 36256
rect 7217 36204 7223 36256
rect 7382 37840 7388 37892
rect 7388 37840 7434 37892
rect 7448 37840 7494 37892
rect 7494 37840 7500 37892
rect 7382 37773 7388 37825
rect 7388 37773 7434 37825
rect 7448 37773 7494 37825
rect 7494 37773 7500 37825
rect 7382 37706 7388 37758
rect 7388 37706 7434 37758
rect 7448 37706 7494 37758
rect 7494 37706 7500 37758
rect 7382 37639 7388 37691
rect 7388 37639 7434 37691
rect 7448 37639 7494 37691
rect 7494 37639 7500 37691
rect 7382 37572 7388 37624
rect 7388 37572 7434 37624
rect 7448 37572 7494 37624
rect 7494 37572 7500 37624
rect 7382 37505 7388 37557
rect 7388 37505 7434 37557
rect 7448 37505 7494 37557
rect 7494 37505 7500 37557
rect 7382 37438 7388 37490
rect 7388 37438 7434 37490
rect 7448 37438 7494 37490
rect 7494 37438 7500 37490
rect 7382 37380 7388 37423
rect 7388 37380 7434 37423
rect 7448 37380 7494 37423
rect 7494 37380 7500 37423
rect 7382 37371 7434 37380
rect 7448 37371 7500 37380
rect 7382 37304 7434 37356
rect 7448 37304 7500 37356
rect 7382 37237 7434 37289
rect 7448 37237 7500 37289
rect 7382 37170 7434 37222
rect 7448 37170 7500 37222
rect 7382 37103 7434 37155
rect 7448 37103 7500 37155
rect 7382 37036 7434 37088
rect 7448 37036 7500 37088
rect 7382 35840 7388 35892
rect 7388 35840 7434 35892
rect 7448 35840 7494 35892
rect 7494 35840 7500 35892
rect 7382 35774 7388 35826
rect 7388 35774 7434 35826
rect 7448 35774 7494 35826
rect 7494 35774 7500 35826
rect 7382 35708 7388 35760
rect 7388 35708 7434 35760
rect 7448 35708 7494 35760
rect 7494 35708 7500 35760
rect 7382 35642 7388 35694
rect 7388 35642 7434 35694
rect 7448 35642 7494 35694
rect 7494 35642 7500 35694
rect 7382 35575 7388 35627
rect 7388 35575 7434 35627
rect 7448 35575 7494 35627
rect 7494 35575 7500 35627
rect 7382 35508 7388 35560
rect 7388 35508 7434 35560
rect 7448 35508 7494 35560
rect 7494 35508 7500 35560
rect 7382 35441 7388 35493
rect 7388 35441 7434 35493
rect 7448 35441 7494 35493
rect 7494 35441 7500 35493
rect 7382 35380 7388 35426
rect 7388 35380 7434 35426
rect 7448 35380 7494 35426
rect 7494 35380 7500 35426
rect 7382 35374 7434 35380
rect 7448 35374 7500 35380
rect 7659 38714 7711 38720
rect 7659 38680 7665 38714
rect 7665 38680 7699 38714
rect 7699 38680 7711 38714
rect 7659 38668 7711 38680
rect 7725 38714 7777 38720
rect 7725 38680 7737 38714
rect 7737 38680 7771 38714
rect 7771 38680 7777 38714
rect 7725 38668 7777 38680
rect 7659 38641 7711 38654
rect 7659 38607 7665 38641
rect 7665 38607 7699 38641
rect 7699 38607 7711 38641
rect 7659 38602 7711 38607
rect 7725 38641 7777 38654
rect 7725 38607 7737 38641
rect 7737 38607 7771 38641
rect 7771 38607 7777 38641
rect 7725 38602 7777 38607
rect 7659 38568 7711 38588
rect 7659 38536 7665 38568
rect 7665 38536 7699 38568
rect 7699 38536 7711 38568
rect 7725 38568 7777 38588
rect 7725 38536 7737 38568
rect 7737 38536 7771 38568
rect 7771 38536 7777 38568
rect 7659 38495 7711 38522
rect 7659 38470 7665 38495
rect 7665 38470 7699 38495
rect 7699 38470 7711 38495
rect 7725 38495 7777 38522
rect 7725 38470 7737 38495
rect 7737 38470 7771 38495
rect 7771 38470 7777 38495
rect 7659 38422 7711 38456
rect 7725 38422 7777 38456
rect 7659 38404 7665 38422
rect 7665 38404 7711 38422
rect 7725 38404 7771 38422
rect 7771 38404 7777 38422
rect 7659 38338 7665 38390
rect 7665 38338 7711 38390
rect 7725 38338 7771 38390
rect 7771 38338 7777 38390
rect 7659 38271 7665 38323
rect 7665 38271 7711 38323
rect 7725 38271 7771 38323
rect 7771 38271 7777 38323
rect 7659 38204 7665 38256
rect 7665 38204 7711 38256
rect 7725 38204 7771 38256
rect 7771 38204 7777 38256
rect 7659 36714 7711 36720
rect 7659 36680 7665 36714
rect 7665 36680 7699 36714
rect 7699 36680 7711 36714
rect 7659 36668 7711 36680
rect 7725 36714 7777 36720
rect 7725 36680 7737 36714
rect 7737 36680 7771 36714
rect 7771 36680 7777 36714
rect 7725 36668 7777 36680
rect 7659 36641 7711 36654
rect 7659 36607 7665 36641
rect 7665 36607 7699 36641
rect 7699 36607 7711 36641
rect 7659 36602 7711 36607
rect 7725 36641 7777 36654
rect 7725 36607 7737 36641
rect 7737 36607 7771 36641
rect 7771 36607 7777 36641
rect 7725 36602 7777 36607
rect 7659 36568 7711 36588
rect 7659 36536 7665 36568
rect 7665 36536 7699 36568
rect 7699 36536 7711 36568
rect 7725 36568 7777 36588
rect 7725 36536 7737 36568
rect 7737 36536 7771 36568
rect 7771 36536 7777 36568
rect 7659 36495 7711 36522
rect 7659 36470 7665 36495
rect 7665 36470 7699 36495
rect 7699 36470 7711 36495
rect 7725 36495 7777 36522
rect 7725 36470 7737 36495
rect 7737 36470 7771 36495
rect 7771 36470 7777 36495
rect 7659 36422 7711 36456
rect 7725 36422 7777 36456
rect 7659 36404 7665 36422
rect 7665 36404 7711 36422
rect 7725 36404 7771 36422
rect 7771 36404 7777 36422
rect 7659 36338 7665 36390
rect 7665 36338 7711 36390
rect 7725 36338 7771 36390
rect 7771 36338 7777 36390
rect 7659 36271 7665 36323
rect 7665 36271 7711 36323
rect 7725 36271 7771 36323
rect 7771 36271 7777 36323
rect 7659 36204 7665 36256
rect 7665 36204 7711 36256
rect 7725 36204 7771 36256
rect 7771 36204 7777 36256
rect 7936 37840 7942 37892
rect 7942 37840 7988 37892
rect 8002 37840 8048 37892
rect 8048 37840 8054 37892
rect 7936 37773 7942 37825
rect 7942 37773 7988 37825
rect 8002 37773 8048 37825
rect 8048 37773 8054 37825
rect 7936 37706 7942 37758
rect 7942 37706 7988 37758
rect 8002 37706 8048 37758
rect 8048 37706 8054 37758
rect 7936 37639 7942 37691
rect 7942 37639 7988 37691
rect 8002 37639 8048 37691
rect 8048 37639 8054 37691
rect 7936 37572 7942 37624
rect 7942 37572 7988 37624
rect 8002 37572 8048 37624
rect 8048 37572 8054 37624
rect 7936 37505 7942 37557
rect 7942 37505 7988 37557
rect 8002 37505 8048 37557
rect 8048 37505 8054 37557
rect 7936 37438 7942 37490
rect 7942 37438 7988 37490
rect 8002 37438 8048 37490
rect 8048 37438 8054 37490
rect 7936 37380 7942 37423
rect 7942 37380 7988 37423
rect 8002 37380 8048 37423
rect 8048 37380 8054 37423
rect 7936 37371 7988 37380
rect 8002 37371 8054 37380
rect 7936 37304 7988 37356
rect 8002 37304 8054 37356
rect 7936 37237 7988 37289
rect 8002 37237 8054 37289
rect 7936 37170 7988 37222
rect 8002 37170 8054 37222
rect 7936 37103 7988 37155
rect 8002 37103 8054 37155
rect 7936 37036 7988 37088
rect 8002 37036 8054 37088
rect 7936 35840 7942 35892
rect 7942 35840 7988 35892
rect 8002 35840 8048 35892
rect 8048 35840 8054 35892
rect 7936 35774 7942 35826
rect 7942 35774 7988 35826
rect 8002 35774 8048 35826
rect 8048 35774 8054 35826
rect 7936 35708 7942 35760
rect 7942 35708 7988 35760
rect 8002 35708 8048 35760
rect 8048 35708 8054 35760
rect 7936 35642 7942 35694
rect 7942 35642 7988 35694
rect 8002 35642 8048 35694
rect 8048 35642 8054 35694
rect 7936 35575 7942 35627
rect 7942 35575 7988 35627
rect 8002 35575 8048 35627
rect 8048 35575 8054 35627
rect 7936 35508 7942 35560
rect 7942 35508 7988 35560
rect 8002 35508 8048 35560
rect 8048 35508 8054 35560
rect 7936 35441 7942 35493
rect 7942 35441 7988 35493
rect 8002 35441 8048 35493
rect 8048 35441 8054 35493
rect 7936 35380 7942 35426
rect 7942 35380 7988 35426
rect 8002 35380 8048 35426
rect 8048 35380 8054 35426
rect 7936 35374 7988 35380
rect 8002 35374 8054 35380
rect 8213 38714 8265 38720
rect 8213 38680 8219 38714
rect 8219 38680 8253 38714
rect 8253 38680 8265 38714
rect 8213 38668 8265 38680
rect 8279 38714 8331 38720
rect 8279 38680 8291 38714
rect 8291 38680 8325 38714
rect 8325 38680 8331 38714
rect 8279 38668 8331 38680
rect 8213 38641 8265 38654
rect 8213 38607 8219 38641
rect 8219 38607 8253 38641
rect 8253 38607 8265 38641
rect 8213 38602 8265 38607
rect 8279 38641 8331 38654
rect 8279 38607 8291 38641
rect 8291 38607 8325 38641
rect 8325 38607 8331 38641
rect 8279 38602 8331 38607
rect 8213 38568 8265 38588
rect 8213 38536 8219 38568
rect 8219 38536 8253 38568
rect 8253 38536 8265 38568
rect 8279 38568 8331 38588
rect 8279 38536 8291 38568
rect 8291 38536 8325 38568
rect 8325 38536 8331 38568
rect 8213 38495 8265 38522
rect 8213 38470 8219 38495
rect 8219 38470 8253 38495
rect 8253 38470 8265 38495
rect 8279 38495 8331 38522
rect 8279 38470 8291 38495
rect 8291 38470 8325 38495
rect 8325 38470 8331 38495
rect 8213 38422 8265 38456
rect 8279 38422 8331 38456
rect 8213 38404 8219 38422
rect 8219 38404 8265 38422
rect 8279 38404 8325 38422
rect 8325 38404 8331 38422
rect 8213 38338 8219 38390
rect 8219 38338 8265 38390
rect 8279 38338 8325 38390
rect 8325 38338 8331 38390
rect 8213 38271 8219 38323
rect 8219 38271 8265 38323
rect 8279 38271 8325 38323
rect 8325 38271 8331 38323
rect 8213 38204 8219 38256
rect 8219 38204 8265 38256
rect 8279 38204 8325 38256
rect 8325 38204 8331 38256
rect 8213 36714 8265 36720
rect 8213 36680 8219 36714
rect 8219 36680 8253 36714
rect 8253 36680 8265 36714
rect 8213 36668 8265 36680
rect 8279 36714 8331 36720
rect 8279 36680 8291 36714
rect 8291 36680 8325 36714
rect 8325 36680 8331 36714
rect 8279 36668 8331 36680
rect 8213 36641 8265 36654
rect 8213 36607 8219 36641
rect 8219 36607 8253 36641
rect 8253 36607 8265 36641
rect 8213 36602 8265 36607
rect 8279 36641 8331 36654
rect 8279 36607 8291 36641
rect 8291 36607 8325 36641
rect 8325 36607 8331 36641
rect 8279 36602 8331 36607
rect 8213 36568 8265 36588
rect 8213 36536 8219 36568
rect 8219 36536 8253 36568
rect 8253 36536 8265 36568
rect 8279 36568 8331 36588
rect 8279 36536 8291 36568
rect 8291 36536 8325 36568
rect 8325 36536 8331 36568
rect 8213 36495 8265 36522
rect 8213 36470 8219 36495
rect 8219 36470 8253 36495
rect 8253 36470 8265 36495
rect 8279 36495 8331 36522
rect 8279 36470 8291 36495
rect 8291 36470 8325 36495
rect 8325 36470 8331 36495
rect 8213 36422 8265 36456
rect 8279 36422 8331 36456
rect 8213 36404 8219 36422
rect 8219 36404 8265 36422
rect 8279 36404 8325 36422
rect 8325 36404 8331 36422
rect 8213 36338 8219 36390
rect 8219 36338 8265 36390
rect 8279 36338 8325 36390
rect 8325 36338 8331 36390
rect 8213 36271 8219 36323
rect 8219 36271 8265 36323
rect 8279 36271 8325 36323
rect 8325 36271 8331 36323
rect 8213 36204 8219 36256
rect 8219 36204 8265 36256
rect 8279 36204 8325 36256
rect 8325 36204 8331 36256
rect 8490 37840 8496 37892
rect 8496 37840 8542 37892
rect 8556 37840 8602 37892
rect 8602 37840 8608 37892
rect 8490 37773 8496 37825
rect 8496 37773 8542 37825
rect 8556 37773 8602 37825
rect 8602 37773 8608 37825
rect 8490 37706 8496 37758
rect 8496 37706 8542 37758
rect 8556 37706 8602 37758
rect 8602 37706 8608 37758
rect 8490 37639 8496 37691
rect 8496 37639 8542 37691
rect 8556 37639 8602 37691
rect 8602 37639 8608 37691
rect 8490 37572 8496 37624
rect 8496 37572 8542 37624
rect 8556 37572 8602 37624
rect 8602 37572 8608 37624
rect 8490 37505 8496 37557
rect 8496 37505 8542 37557
rect 8556 37505 8602 37557
rect 8602 37505 8608 37557
rect 8490 37438 8496 37490
rect 8496 37438 8542 37490
rect 8556 37438 8602 37490
rect 8602 37438 8608 37490
rect 8490 37380 8496 37423
rect 8496 37380 8542 37423
rect 8556 37380 8602 37423
rect 8602 37380 8608 37423
rect 8490 37371 8542 37380
rect 8556 37371 8608 37380
rect 8490 37304 8542 37356
rect 8556 37304 8608 37356
rect 8490 37237 8542 37289
rect 8556 37237 8608 37289
rect 8490 37170 8542 37222
rect 8556 37170 8608 37222
rect 8490 37103 8542 37155
rect 8556 37103 8608 37155
rect 8490 37036 8542 37088
rect 8556 37036 8608 37088
rect 8490 35840 8496 35892
rect 8496 35840 8542 35892
rect 8556 35840 8602 35892
rect 8602 35840 8608 35892
rect 8490 35774 8496 35826
rect 8496 35774 8542 35826
rect 8556 35774 8602 35826
rect 8602 35774 8608 35826
rect 8490 35708 8496 35760
rect 8496 35708 8542 35760
rect 8556 35708 8602 35760
rect 8602 35708 8608 35760
rect 8490 35642 8496 35694
rect 8496 35642 8542 35694
rect 8556 35642 8602 35694
rect 8602 35642 8608 35694
rect 8490 35575 8496 35627
rect 8496 35575 8542 35627
rect 8556 35575 8602 35627
rect 8602 35575 8608 35627
rect 8490 35508 8496 35560
rect 8496 35508 8542 35560
rect 8556 35508 8602 35560
rect 8602 35508 8608 35560
rect 8490 35441 8496 35493
rect 8496 35441 8542 35493
rect 8556 35441 8602 35493
rect 8602 35441 8608 35493
rect 8490 35380 8496 35426
rect 8496 35380 8542 35426
rect 8556 35380 8602 35426
rect 8602 35380 8608 35426
rect 8490 35374 8542 35380
rect 8556 35374 8608 35380
rect 8767 38714 8819 38720
rect 8767 38680 8773 38714
rect 8773 38680 8807 38714
rect 8807 38680 8819 38714
rect 8767 38668 8819 38680
rect 8833 38714 8885 38720
rect 8833 38680 8845 38714
rect 8845 38680 8879 38714
rect 8879 38680 8885 38714
rect 8833 38668 8885 38680
rect 8767 38641 8819 38654
rect 8767 38607 8773 38641
rect 8773 38607 8807 38641
rect 8807 38607 8819 38641
rect 8767 38602 8819 38607
rect 8833 38641 8885 38654
rect 8833 38607 8845 38641
rect 8845 38607 8879 38641
rect 8879 38607 8885 38641
rect 8833 38602 8885 38607
rect 8767 38568 8819 38588
rect 8767 38536 8773 38568
rect 8773 38536 8807 38568
rect 8807 38536 8819 38568
rect 8833 38568 8885 38588
rect 8833 38536 8845 38568
rect 8845 38536 8879 38568
rect 8879 38536 8885 38568
rect 8767 38495 8819 38522
rect 8767 38470 8773 38495
rect 8773 38470 8807 38495
rect 8807 38470 8819 38495
rect 8833 38495 8885 38522
rect 8833 38470 8845 38495
rect 8845 38470 8879 38495
rect 8879 38470 8885 38495
rect 8767 38422 8819 38456
rect 8833 38422 8885 38456
rect 8767 38404 8773 38422
rect 8773 38404 8819 38422
rect 8833 38404 8879 38422
rect 8879 38404 8885 38422
rect 8767 38338 8773 38390
rect 8773 38338 8819 38390
rect 8833 38338 8879 38390
rect 8879 38338 8885 38390
rect 8767 38271 8773 38323
rect 8773 38271 8819 38323
rect 8833 38271 8879 38323
rect 8879 38271 8885 38323
rect 8767 38204 8773 38256
rect 8773 38204 8819 38256
rect 8833 38204 8879 38256
rect 8879 38204 8885 38256
rect 8767 36714 8819 36720
rect 8767 36680 8773 36714
rect 8773 36680 8807 36714
rect 8807 36680 8819 36714
rect 8767 36668 8819 36680
rect 8833 36714 8885 36720
rect 8833 36680 8845 36714
rect 8845 36680 8879 36714
rect 8879 36680 8885 36714
rect 8833 36668 8885 36680
rect 8767 36641 8819 36654
rect 8767 36607 8773 36641
rect 8773 36607 8807 36641
rect 8807 36607 8819 36641
rect 8767 36602 8819 36607
rect 8833 36641 8885 36654
rect 8833 36607 8845 36641
rect 8845 36607 8879 36641
rect 8879 36607 8885 36641
rect 8833 36602 8885 36607
rect 8767 36568 8819 36588
rect 8767 36536 8773 36568
rect 8773 36536 8807 36568
rect 8807 36536 8819 36568
rect 8833 36568 8885 36588
rect 8833 36536 8845 36568
rect 8845 36536 8879 36568
rect 8879 36536 8885 36568
rect 8767 36495 8819 36522
rect 8767 36470 8773 36495
rect 8773 36470 8807 36495
rect 8807 36470 8819 36495
rect 8833 36495 8885 36522
rect 8833 36470 8845 36495
rect 8845 36470 8879 36495
rect 8879 36470 8885 36495
rect 8767 36422 8819 36456
rect 8833 36422 8885 36456
rect 8767 36404 8773 36422
rect 8773 36404 8819 36422
rect 8833 36404 8879 36422
rect 8879 36404 8885 36422
rect 8767 36338 8773 36390
rect 8773 36338 8819 36390
rect 8833 36338 8879 36390
rect 8879 36338 8885 36390
rect 8767 36271 8773 36323
rect 8773 36271 8819 36323
rect 8833 36271 8879 36323
rect 8879 36271 8885 36323
rect 8767 36204 8773 36256
rect 8773 36204 8819 36256
rect 8833 36204 8879 36256
rect 8879 36204 8885 36256
rect 9044 37840 9050 37892
rect 9050 37840 9096 37892
rect 9110 37840 9156 37892
rect 9156 37840 9162 37892
rect 9044 37773 9050 37825
rect 9050 37773 9096 37825
rect 9110 37773 9156 37825
rect 9156 37773 9162 37825
rect 9044 37706 9050 37758
rect 9050 37706 9096 37758
rect 9110 37706 9156 37758
rect 9156 37706 9162 37758
rect 9044 37639 9050 37691
rect 9050 37639 9096 37691
rect 9110 37639 9156 37691
rect 9156 37639 9162 37691
rect 9044 37572 9050 37624
rect 9050 37572 9096 37624
rect 9110 37572 9156 37624
rect 9156 37572 9162 37624
rect 9044 37505 9050 37557
rect 9050 37505 9096 37557
rect 9110 37505 9156 37557
rect 9156 37505 9162 37557
rect 9044 37438 9050 37490
rect 9050 37438 9096 37490
rect 9110 37438 9156 37490
rect 9156 37438 9162 37490
rect 9044 37380 9050 37423
rect 9050 37380 9096 37423
rect 9110 37380 9156 37423
rect 9156 37380 9162 37423
rect 9044 37371 9096 37380
rect 9110 37371 9162 37380
rect 9044 37304 9096 37356
rect 9110 37304 9162 37356
rect 9044 37237 9096 37289
rect 9110 37237 9162 37289
rect 9044 37170 9096 37222
rect 9110 37170 9162 37222
rect 9044 37103 9096 37155
rect 9110 37103 9162 37155
rect 9044 37036 9096 37088
rect 9110 37036 9162 37088
rect 9044 35840 9050 35892
rect 9050 35840 9096 35892
rect 9110 35840 9156 35892
rect 9156 35840 9162 35892
rect 9044 35774 9050 35826
rect 9050 35774 9096 35826
rect 9110 35774 9156 35826
rect 9156 35774 9162 35826
rect 9044 35708 9050 35760
rect 9050 35708 9096 35760
rect 9110 35708 9156 35760
rect 9156 35708 9162 35760
rect 9044 35642 9050 35694
rect 9050 35642 9096 35694
rect 9110 35642 9156 35694
rect 9156 35642 9162 35694
rect 9044 35575 9050 35627
rect 9050 35575 9096 35627
rect 9110 35575 9156 35627
rect 9156 35575 9162 35627
rect 9044 35508 9050 35560
rect 9050 35508 9096 35560
rect 9110 35508 9156 35560
rect 9156 35508 9162 35560
rect 9044 35441 9050 35493
rect 9050 35441 9096 35493
rect 9110 35441 9156 35493
rect 9156 35441 9162 35493
rect 9044 35380 9050 35426
rect 9050 35380 9096 35426
rect 9110 35380 9156 35426
rect 9156 35380 9162 35426
rect 9044 35374 9096 35380
rect 9110 35374 9162 35380
rect 9321 38714 9373 38720
rect 9321 38680 9327 38714
rect 9327 38680 9361 38714
rect 9361 38680 9373 38714
rect 9321 38668 9373 38680
rect 9387 38714 9439 38720
rect 9387 38680 9399 38714
rect 9399 38680 9433 38714
rect 9433 38680 9439 38714
rect 9387 38668 9439 38680
rect 9321 38641 9373 38654
rect 9321 38607 9327 38641
rect 9327 38607 9361 38641
rect 9361 38607 9373 38641
rect 9321 38602 9373 38607
rect 9387 38641 9439 38654
rect 9387 38607 9399 38641
rect 9399 38607 9433 38641
rect 9433 38607 9439 38641
rect 9387 38602 9439 38607
rect 9321 38568 9373 38588
rect 9321 38536 9327 38568
rect 9327 38536 9361 38568
rect 9361 38536 9373 38568
rect 9387 38568 9439 38588
rect 9387 38536 9399 38568
rect 9399 38536 9433 38568
rect 9433 38536 9439 38568
rect 9321 38495 9373 38522
rect 9321 38470 9327 38495
rect 9327 38470 9361 38495
rect 9361 38470 9373 38495
rect 9387 38495 9439 38522
rect 9387 38470 9399 38495
rect 9399 38470 9433 38495
rect 9433 38470 9439 38495
rect 9321 38422 9373 38456
rect 9387 38422 9439 38456
rect 9321 38404 9327 38422
rect 9327 38404 9373 38422
rect 9387 38404 9433 38422
rect 9433 38404 9439 38422
rect 9321 38338 9327 38390
rect 9327 38338 9373 38390
rect 9387 38338 9433 38390
rect 9433 38338 9439 38390
rect 9321 38271 9327 38323
rect 9327 38271 9373 38323
rect 9387 38271 9433 38323
rect 9433 38271 9439 38323
rect 9321 38204 9327 38256
rect 9327 38204 9373 38256
rect 9387 38204 9433 38256
rect 9433 38204 9439 38256
rect 9321 36714 9373 36720
rect 9321 36680 9327 36714
rect 9327 36680 9361 36714
rect 9361 36680 9373 36714
rect 9321 36668 9373 36680
rect 9387 36714 9439 36720
rect 9387 36680 9399 36714
rect 9399 36680 9433 36714
rect 9433 36680 9439 36714
rect 9387 36668 9439 36680
rect 9321 36641 9373 36654
rect 9321 36607 9327 36641
rect 9327 36607 9361 36641
rect 9361 36607 9373 36641
rect 9321 36602 9373 36607
rect 9387 36641 9439 36654
rect 9387 36607 9399 36641
rect 9399 36607 9433 36641
rect 9433 36607 9439 36641
rect 9387 36602 9439 36607
rect 9321 36568 9373 36588
rect 9321 36536 9327 36568
rect 9327 36536 9361 36568
rect 9361 36536 9373 36568
rect 9387 36568 9439 36588
rect 9387 36536 9399 36568
rect 9399 36536 9433 36568
rect 9433 36536 9439 36568
rect 9321 36495 9373 36522
rect 9321 36470 9327 36495
rect 9327 36470 9361 36495
rect 9361 36470 9373 36495
rect 9387 36495 9439 36522
rect 9387 36470 9399 36495
rect 9399 36470 9433 36495
rect 9433 36470 9439 36495
rect 9321 36422 9373 36456
rect 9387 36422 9439 36456
rect 9321 36404 9327 36422
rect 9327 36404 9373 36422
rect 9387 36404 9433 36422
rect 9433 36404 9439 36422
rect 9321 36338 9327 36390
rect 9327 36338 9373 36390
rect 9387 36338 9433 36390
rect 9433 36338 9439 36390
rect 9321 36271 9327 36323
rect 9327 36271 9373 36323
rect 9387 36271 9433 36323
rect 9433 36271 9439 36323
rect 9321 36204 9327 36256
rect 9327 36204 9373 36256
rect 9387 36204 9433 36256
rect 9433 36204 9439 36256
rect 9598 37840 9604 37892
rect 9604 37840 9650 37892
rect 9664 37840 9710 37892
rect 9710 37840 9716 37892
rect 9598 37773 9604 37825
rect 9604 37773 9650 37825
rect 9664 37773 9710 37825
rect 9710 37773 9716 37825
rect 9598 37706 9604 37758
rect 9604 37706 9650 37758
rect 9664 37706 9710 37758
rect 9710 37706 9716 37758
rect 9598 37639 9604 37691
rect 9604 37639 9650 37691
rect 9664 37639 9710 37691
rect 9710 37639 9716 37691
rect 9598 37572 9604 37624
rect 9604 37572 9650 37624
rect 9664 37572 9710 37624
rect 9710 37572 9716 37624
rect 9598 37505 9604 37557
rect 9604 37505 9650 37557
rect 9664 37505 9710 37557
rect 9710 37505 9716 37557
rect 9598 37438 9604 37490
rect 9604 37438 9650 37490
rect 9664 37438 9710 37490
rect 9710 37438 9716 37490
rect 9598 37380 9604 37423
rect 9604 37380 9650 37423
rect 9664 37380 9710 37423
rect 9710 37380 9716 37423
rect 9598 37371 9650 37380
rect 9664 37371 9716 37380
rect 9598 37304 9650 37356
rect 9664 37304 9716 37356
rect 9598 37237 9650 37289
rect 9664 37237 9716 37289
rect 9598 37170 9650 37222
rect 9664 37170 9716 37222
rect 9598 37103 9650 37155
rect 9664 37103 9716 37155
rect 9598 37036 9650 37088
rect 9664 37036 9716 37088
rect 9598 35840 9604 35892
rect 9604 35840 9650 35892
rect 9664 35840 9710 35892
rect 9710 35840 9716 35892
rect 9598 35774 9604 35826
rect 9604 35774 9650 35826
rect 9664 35774 9710 35826
rect 9710 35774 9716 35826
rect 9598 35708 9604 35760
rect 9604 35708 9650 35760
rect 9664 35708 9710 35760
rect 9710 35708 9716 35760
rect 9598 35642 9604 35694
rect 9604 35642 9650 35694
rect 9664 35642 9710 35694
rect 9710 35642 9716 35694
rect 9598 35575 9604 35627
rect 9604 35575 9650 35627
rect 9664 35575 9710 35627
rect 9710 35575 9716 35627
rect 9598 35508 9604 35560
rect 9604 35508 9650 35560
rect 9664 35508 9710 35560
rect 9710 35508 9716 35560
rect 9598 35441 9604 35493
rect 9604 35441 9650 35493
rect 9664 35441 9710 35493
rect 9710 35441 9716 35493
rect 9598 35380 9604 35426
rect 9604 35380 9650 35426
rect 9664 35380 9710 35426
rect 9710 35380 9716 35426
rect 9598 35374 9650 35380
rect 9664 35374 9716 35380
rect 9875 38714 9927 38720
rect 9875 38680 9881 38714
rect 9881 38680 9915 38714
rect 9915 38680 9927 38714
rect 9875 38668 9927 38680
rect 9941 38714 9993 38720
rect 9941 38680 9953 38714
rect 9953 38680 9987 38714
rect 9987 38680 9993 38714
rect 9941 38668 9993 38680
rect 9875 38641 9927 38654
rect 9875 38607 9881 38641
rect 9881 38607 9915 38641
rect 9915 38607 9927 38641
rect 9875 38602 9927 38607
rect 9941 38641 9993 38654
rect 9941 38607 9953 38641
rect 9953 38607 9987 38641
rect 9987 38607 9993 38641
rect 9941 38602 9993 38607
rect 9875 38568 9927 38588
rect 9875 38536 9881 38568
rect 9881 38536 9915 38568
rect 9915 38536 9927 38568
rect 9941 38568 9993 38588
rect 9941 38536 9953 38568
rect 9953 38536 9987 38568
rect 9987 38536 9993 38568
rect 9875 38495 9927 38522
rect 9875 38470 9881 38495
rect 9881 38470 9915 38495
rect 9915 38470 9927 38495
rect 9941 38495 9993 38522
rect 9941 38470 9953 38495
rect 9953 38470 9987 38495
rect 9987 38470 9993 38495
rect 9875 38422 9927 38456
rect 9941 38422 9993 38456
rect 9875 38404 9881 38422
rect 9881 38404 9927 38422
rect 9941 38404 9987 38422
rect 9987 38404 9993 38422
rect 9875 38338 9881 38390
rect 9881 38338 9927 38390
rect 9941 38338 9987 38390
rect 9987 38338 9993 38390
rect 9875 38271 9881 38323
rect 9881 38271 9927 38323
rect 9941 38271 9987 38323
rect 9987 38271 9993 38323
rect 9875 38204 9881 38256
rect 9881 38204 9927 38256
rect 9941 38204 9987 38256
rect 9987 38204 9993 38256
rect 9875 36714 9927 36720
rect 9875 36680 9881 36714
rect 9881 36680 9915 36714
rect 9915 36680 9927 36714
rect 9875 36668 9927 36680
rect 9941 36714 9993 36720
rect 9941 36680 9953 36714
rect 9953 36680 9987 36714
rect 9987 36680 9993 36714
rect 9941 36668 9993 36680
rect 9875 36641 9927 36654
rect 9875 36607 9881 36641
rect 9881 36607 9915 36641
rect 9915 36607 9927 36641
rect 9875 36602 9927 36607
rect 9941 36641 9993 36654
rect 9941 36607 9953 36641
rect 9953 36607 9987 36641
rect 9987 36607 9993 36641
rect 9941 36602 9993 36607
rect 9875 36568 9927 36588
rect 9875 36536 9881 36568
rect 9881 36536 9915 36568
rect 9915 36536 9927 36568
rect 9941 36568 9993 36588
rect 9941 36536 9953 36568
rect 9953 36536 9987 36568
rect 9987 36536 9993 36568
rect 9875 36495 9927 36522
rect 9875 36470 9881 36495
rect 9881 36470 9915 36495
rect 9915 36470 9927 36495
rect 9941 36495 9993 36522
rect 9941 36470 9953 36495
rect 9953 36470 9987 36495
rect 9987 36470 9993 36495
rect 9875 36422 9927 36456
rect 9941 36422 9993 36456
rect 9875 36404 9881 36422
rect 9881 36404 9927 36422
rect 9941 36404 9987 36422
rect 9987 36404 9993 36422
rect 9875 36338 9881 36390
rect 9881 36338 9927 36390
rect 9941 36338 9987 36390
rect 9987 36338 9993 36390
rect 9875 36271 9881 36323
rect 9881 36271 9927 36323
rect 9941 36271 9987 36323
rect 9987 36271 9993 36323
rect 9875 36204 9881 36256
rect 9881 36204 9927 36256
rect 9941 36204 9987 36256
rect 9987 36204 9993 36256
rect 10152 37840 10158 37892
rect 10158 37840 10204 37892
rect 10218 37840 10264 37892
rect 10264 37840 10270 37892
rect 10152 37773 10158 37825
rect 10158 37773 10204 37825
rect 10218 37773 10264 37825
rect 10264 37773 10270 37825
rect 10152 37706 10158 37758
rect 10158 37706 10204 37758
rect 10218 37706 10264 37758
rect 10264 37706 10270 37758
rect 10152 37639 10158 37691
rect 10158 37639 10204 37691
rect 10218 37639 10264 37691
rect 10264 37639 10270 37691
rect 10152 37572 10158 37624
rect 10158 37572 10204 37624
rect 10218 37572 10264 37624
rect 10264 37572 10270 37624
rect 10152 37505 10158 37557
rect 10158 37505 10204 37557
rect 10218 37505 10264 37557
rect 10264 37505 10270 37557
rect 10152 37438 10158 37490
rect 10158 37438 10204 37490
rect 10218 37438 10264 37490
rect 10264 37438 10270 37490
rect 10152 37380 10158 37423
rect 10158 37380 10204 37423
rect 10218 37380 10264 37423
rect 10264 37380 10270 37423
rect 10152 37371 10204 37380
rect 10218 37371 10270 37380
rect 10152 37304 10204 37356
rect 10218 37304 10270 37356
rect 10152 37237 10204 37289
rect 10218 37237 10270 37289
rect 10152 37170 10204 37222
rect 10218 37170 10270 37222
rect 10152 37103 10204 37155
rect 10218 37103 10270 37155
rect 10152 37036 10204 37088
rect 10218 37036 10270 37088
rect 10152 35840 10158 35892
rect 10158 35840 10204 35892
rect 10218 35840 10264 35892
rect 10264 35840 10270 35892
rect 10152 35774 10158 35826
rect 10158 35774 10204 35826
rect 10218 35774 10264 35826
rect 10264 35774 10270 35826
rect 10152 35708 10158 35760
rect 10158 35708 10204 35760
rect 10218 35708 10264 35760
rect 10264 35708 10270 35760
rect 10152 35642 10158 35694
rect 10158 35642 10204 35694
rect 10218 35642 10264 35694
rect 10264 35642 10270 35694
rect 10152 35575 10158 35627
rect 10158 35575 10204 35627
rect 10218 35575 10264 35627
rect 10264 35575 10270 35627
rect 10152 35508 10158 35560
rect 10158 35508 10204 35560
rect 10218 35508 10264 35560
rect 10264 35508 10270 35560
rect 10152 35441 10158 35493
rect 10158 35441 10204 35493
rect 10218 35441 10264 35493
rect 10264 35441 10270 35493
rect 10152 35380 10158 35426
rect 10158 35380 10204 35426
rect 10218 35380 10264 35426
rect 10264 35380 10270 35426
rect 10152 35374 10204 35380
rect 10218 35374 10270 35380
rect 10429 38714 10481 38720
rect 10429 38680 10435 38714
rect 10435 38680 10469 38714
rect 10469 38680 10481 38714
rect 10429 38668 10481 38680
rect 10495 38714 10547 38720
rect 10495 38680 10507 38714
rect 10507 38680 10541 38714
rect 10541 38680 10547 38714
rect 10495 38668 10547 38680
rect 10429 38641 10481 38654
rect 10429 38607 10435 38641
rect 10435 38607 10469 38641
rect 10469 38607 10481 38641
rect 10429 38602 10481 38607
rect 10495 38641 10547 38654
rect 10495 38607 10507 38641
rect 10507 38607 10541 38641
rect 10541 38607 10547 38641
rect 10495 38602 10547 38607
rect 10429 38568 10481 38588
rect 10429 38536 10435 38568
rect 10435 38536 10469 38568
rect 10469 38536 10481 38568
rect 10495 38568 10547 38588
rect 10495 38536 10507 38568
rect 10507 38536 10541 38568
rect 10541 38536 10547 38568
rect 10429 38495 10481 38522
rect 10429 38470 10435 38495
rect 10435 38470 10469 38495
rect 10469 38470 10481 38495
rect 10495 38495 10547 38522
rect 10495 38470 10507 38495
rect 10507 38470 10541 38495
rect 10541 38470 10547 38495
rect 10429 38422 10481 38456
rect 10495 38422 10547 38456
rect 10429 38404 10435 38422
rect 10435 38404 10481 38422
rect 10495 38404 10541 38422
rect 10541 38404 10547 38422
rect 10429 38338 10435 38390
rect 10435 38338 10481 38390
rect 10495 38338 10541 38390
rect 10541 38338 10547 38390
rect 10429 38271 10435 38323
rect 10435 38271 10481 38323
rect 10495 38271 10541 38323
rect 10541 38271 10547 38323
rect 10429 38204 10435 38256
rect 10435 38204 10481 38256
rect 10495 38204 10541 38256
rect 10541 38204 10547 38256
rect 10429 36714 10481 36720
rect 10429 36680 10435 36714
rect 10435 36680 10469 36714
rect 10469 36680 10481 36714
rect 10429 36668 10481 36680
rect 10495 36714 10547 36720
rect 10495 36680 10507 36714
rect 10507 36680 10541 36714
rect 10541 36680 10547 36714
rect 10495 36668 10547 36680
rect 10429 36641 10481 36654
rect 10429 36607 10435 36641
rect 10435 36607 10469 36641
rect 10469 36607 10481 36641
rect 10429 36602 10481 36607
rect 10495 36641 10547 36654
rect 10495 36607 10507 36641
rect 10507 36607 10541 36641
rect 10541 36607 10547 36641
rect 10495 36602 10547 36607
rect 10429 36568 10481 36588
rect 10429 36536 10435 36568
rect 10435 36536 10469 36568
rect 10469 36536 10481 36568
rect 10495 36568 10547 36588
rect 10495 36536 10507 36568
rect 10507 36536 10541 36568
rect 10541 36536 10547 36568
rect 10429 36495 10481 36522
rect 10429 36470 10435 36495
rect 10435 36470 10469 36495
rect 10469 36470 10481 36495
rect 10495 36495 10547 36522
rect 10495 36470 10507 36495
rect 10507 36470 10541 36495
rect 10541 36470 10547 36495
rect 10429 36422 10481 36456
rect 10495 36422 10547 36456
rect 10429 36404 10435 36422
rect 10435 36404 10481 36422
rect 10495 36404 10541 36422
rect 10541 36404 10547 36422
rect 10429 36338 10435 36390
rect 10435 36338 10481 36390
rect 10495 36338 10541 36390
rect 10541 36338 10547 36390
rect 10429 36271 10435 36323
rect 10435 36271 10481 36323
rect 10495 36271 10541 36323
rect 10541 36271 10547 36323
rect 10429 36204 10435 36256
rect 10435 36204 10481 36256
rect 10495 36204 10541 36256
rect 10541 36204 10547 36256
rect 10706 37840 10712 37892
rect 10712 37840 10758 37892
rect 10772 37840 10818 37892
rect 10818 37840 10824 37892
rect 10706 37773 10712 37825
rect 10712 37773 10758 37825
rect 10772 37773 10818 37825
rect 10818 37773 10824 37825
rect 10706 37706 10712 37758
rect 10712 37706 10758 37758
rect 10772 37706 10818 37758
rect 10818 37706 10824 37758
rect 10706 37639 10712 37691
rect 10712 37639 10758 37691
rect 10772 37639 10818 37691
rect 10818 37639 10824 37691
rect 10706 37572 10712 37624
rect 10712 37572 10758 37624
rect 10772 37572 10818 37624
rect 10818 37572 10824 37624
rect 10706 37505 10712 37557
rect 10712 37505 10758 37557
rect 10772 37505 10818 37557
rect 10818 37505 10824 37557
rect 10706 37438 10712 37490
rect 10712 37438 10758 37490
rect 10772 37438 10818 37490
rect 10818 37438 10824 37490
rect 10706 37380 10712 37423
rect 10712 37380 10758 37423
rect 10772 37380 10818 37423
rect 10818 37380 10824 37423
rect 10706 37371 10758 37380
rect 10772 37371 10824 37380
rect 10706 37304 10758 37356
rect 10772 37304 10824 37356
rect 10706 37237 10758 37289
rect 10772 37237 10824 37289
rect 10706 37170 10758 37222
rect 10772 37170 10824 37222
rect 10706 37103 10758 37155
rect 10772 37103 10824 37155
rect 10706 37036 10758 37088
rect 10772 37036 10824 37088
rect 10706 35840 10712 35892
rect 10712 35840 10758 35892
rect 10772 35840 10818 35892
rect 10818 35840 10824 35892
rect 10706 35774 10712 35826
rect 10712 35774 10758 35826
rect 10772 35774 10818 35826
rect 10818 35774 10824 35826
rect 10706 35708 10712 35760
rect 10712 35708 10758 35760
rect 10772 35708 10818 35760
rect 10818 35708 10824 35760
rect 10706 35642 10712 35694
rect 10712 35642 10758 35694
rect 10772 35642 10818 35694
rect 10818 35642 10824 35694
rect 10706 35575 10712 35627
rect 10712 35575 10758 35627
rect 10772 35575 10818 35627
rect 10818 35575 10824 35627
rect 10706 35508 10712 35560
rect 10712 35508 10758 35560
rect 10772 35508 10818 35560
rect 10818 35508 10824 35560
rect 10706 35441 10712 35493
rect 10712 35441 10758 35493
rect 10772 35441 10818 35493
rect 10818 35441 10824 35493
rect 10706 35380 10712 35426
rect 10712 35380 10758 35426
rect 10772 35380 10818 35426
rect 10818 35380 10824 35426
rect 10706 35374 10758 35380
rect 10772 35374 10824 35380
rect 10983 38714 11035 38720
rect 10983 38680 10989 38714
rect 10989 38680 11023 38714
rect 11023 38680 11035 38714
rect 10983 38668 11035 38680
rect 11049 38714 11101 38720
rect 11049 38680 11061 38714
rect 11061 38680 11095 38714
rect 11095 38680 11101 38714
rect 11049 38668 11101 38680
rect 10983 38641 11035 38654
rect 10983 38607 10989 38641
rect 10989 38607 11023 38641
rect 11023 38607 11035 38641
rect 10983 38602 11035 38607
rect 11049 38641 11101 38654
rect 11049 38607 11061 38641
rect 11061 38607 11095 38641
rect 11095 38607 11101 38641
rect 11049 38602 11101 38607
rect 10983 38568 11035 38588
rect 10983 38536 10989 38568
rect 10989 38536 11023 38568
rect 11023 38536 11035 38568
rect 11049 38568 11101 38588
rect 11049 38536 11061 38568
rect 11061 38536 11095 38568
rect 11095 38536 11101 38568
rect 10983 38495 11035 38522
rect 10983 38470 10989 38495
rect 10989 38470 11023 38495
rect 11023 38470 11035 38495
rect 11049 38495 11101 38522
rect 11049 38470 11061 38495
rect 11061 38470 11095 38495
rect 11095 38470 11101 38495
rect 10983 38422 11035 38456
rect 11049 38422 11101 38456
rect 10983 38404 10989 38422
rect 10989 38404 11035 38422
rect 11049 38404 11095 38422
rect 11095 38404 11101 38422
rect 10983 38338 10989 38390
rect 10989 38338 11035 38390
rect 11049 38338 11095 38390
rect 11095 38338 11101 38390
rect 10983 38271 10989 38323
rect 10989 38271 11035 38323
rect 11049 38271 11095 38323
rect 11095 38271 11101 38323
rect 10983 38204 10989 38256
rect 10989 38204 11035 38256
rect 11049 38204 11095 38256
rect 11095 38204 11101 38256
rect 10983 36714 11035 36720
rect 10983 36680 10989 36714
rect 10989 36680 11023 36714
rect 11023 36680 11035 36714
rect 10983 36668 11035 36680
rect 11049 36714 11101 36720
rect 11049 36680 11061 36714
rect 11061 36680 11095 36714
rect 11095 36680 11101 36714
rect 11049 36668 11101 36680
rect 10983 36641 11035 36654
rect 10983 36607 10989 36641
rect 10989 36607 11023 36641
rect 11023 36607 11035 36641
rect 10983 36602 11035 36607
rect 11049 36641 11101 36654
rect 11049 36607 11061 36641
rect 11061 36607 11095 36641
rect 11095 36607 11101 36641
rect 11049 36602 11101 36607
rect 10983 36568 11035 36588
rect 10983 36536 10989 36568
rect 10989 36536 11023 36568
rect 11023 36536 11035 36568
rect 11049 36568 11101 36588
rect 11049 36536 11061 36568
rect 11061 36536 11095 36568
rect 11095 36536 11101 36568
rect 10983 36495 11035 36522
rect 10983 36470 10989 36495
rect 10989 36470 11023 36495
rect 11023 36470 11035 36495
rect 11049 36495 11101 36522
rect 11049 36470 11061 36495
rect 11061 36470 11095 36495
rect 11095 36470 11101 36495
rect 10983 36422 11035 36456
rect 11049 36422 11101 36456
rect 10983 36404 10989 36422
rect 10989 36404 11035 36422
rect 11049 36404 11095 36422
rect 11095 36404 11101 36422
rect 10983 36338 10989 36390
rect 10989 36338 11035 36390
rect 11049 36338 11095 36390
rect 11095 36338 11101 36390
rect 10983 36271 10989 36323
rect 10989 36271 11035 36323
rect 11049 36271 11095 36323
rect 11095 36271 11101 36323
rect 10983 36204 10989 36256
rect 10989 36204 11035 36256
rect 11049 36204 11095 36256
rect 11095 36204 11101 36256
rect 11260 37840 11266 37892
rect 11266 37840 11312 37892
rect 11326 37840 11372 37892
rect 11372 37840 11378 37892
rect 11260 37773 11266 37825
rect 11266 37773 11312 37825
rect 11326 37773 11372 37825
rect 11372 37773 11378 37825
rect 11260 37706 11266 37758
rect 11266 37706 11312 37758
rect 11326 37706 11372 37758
rect 11372 37706 11378 37758
rect 11260 37639 11266 37691
rect 11266 37639 11312 37691
rect 11326 37639 11372 37691
rect 11372 37639 11378 37691
rect 11260 37572 11266 37624
rect 11266 37572 11312 37624
rect 11326 37572 11372 37624
rect 11372 37572 11378 37624
rect 11260 37505 11266 37557
rect 11266 37505 11312 37557
rect 11326 37505 11372 37557
rect 11372 37505 11378 37557
rect 11260 37438 11266 37490
rect 11266 37438 11312 37490
rect 11326 37438 11372 37490
rect 11372 37438 11378 37490
rect 11260 37380 11266 37423
rect 11266 37380 11312 37423
rect 11326 37380 11372 37423
rect 11372 37380 11378 37423
rect 11260 37371 11312 37380
rect 11326 37371 11378 37380
rect 11260 37304 11312 37356
rect 11326 37304 11378 37356
rect 11260 37237 11312 37289
rect 11326 37237 11378 37289
rect 11260 37170 11312 37222
rect 11326 37170 11378 37222
rect 11260 37103 11312 37155
rect 11326 37103 11378 37155
rect 11260 37036 11312 37088
rect 11326 37036 11378 37088
rect 11260 35840 11266 35892
rect 11266 35840 11312 35892
rect 11326 35840 11372 35892
rect 11372 35840 11378 35892
rect 11260 35774 11266 35826
rect 11266 35774 11312 35826
rect 11326 35774 11372 35826
rect 11372 35774 11378 35826
rect 11260 35708 11266 35760
rect 11266 35708 11312 35760
rect 11326 35708 11372 35760
rect 11372 35708 11378 35760
rect 11260 35642 11266 35694
rect 11266 35642 11312 35694
rect 11326 35642 11372 35694
rect 11372 35642 11378 35694
rect 11260 35575 11266 35627
rect 11266 35575 11312 35627
rect 11326 35575 11372 35627
rect 11372 35575 11378 35627
rect 11260 35508 11266 35560
rect 11266 35508 11312 35560
rect 11326 35508 11372 35560
rect 11372 35508 11378 35560
rect 11260 35441 11266 35493
rect 11266 35441 11312 35493
rect 11326 35441 11372 35493
rect 11372 35441 11378 35493
rect 11260 35380 11266 35426
rect 11266 35380 11312 35426
rect 11326 35380 11372 35426
rect 11372 35380 11378 35426
rect 11260 35374 11312 35380
rect 11326 35374 11378 35380
rect 11537 38714 11589 38720
rect 11537 38680 11543 38714
rect 11543 38680 11577 38714
rect 11577 38680 11589 38714
rect 11537 38668 11589 38680
rect 11603 38714 11655 38720
rect 11603 38680 11615 38714
rect 11615 38680 11649 38714
rect 11649 38680 11655 38714
rect 11603 38668 11655 38680
rect 11537 38641 11589 38654
rect 11537 38607 11543 38641
rect 11543 38607 11577 38641
rect 11577 38607 11589 38641
rect 11537 38602 11589 38607
rect 11603 38641 11655 38654
rect 11603 38607 11615 38641
rect 11615 38607 11649 38641
rect 11649 38607 11655 38641
rect 11603 38602 11655 38607
rect 11537 38568 11589 38588
rect 11537 38536 11543 38568
rect 11543 38536 11577 38568
rect 11577 38536 11589 38568
rect 11603 38568 11655 38588
rect 11603 38536 11615 38568
rect 11615 38536 11649 38568
rect 11649 38536 11655 38568
rect 11537 38495 11589 38522
rect 11537 38470 11543 38495
rect 11543 38470 11577 38495
rect 11577 38470 11589 38495
rect 11603 38495 11655 38522
rect 11603 38470 11615 38495
rect 11615 38470 11649 38495
rect 11649 38470 11655 38495
rect 11537 38422 11589 38456
rect 11603 38422 11655 38456
rect 11537 38404 11543 38422
rect 11543 38404 11589 38422
rect 11603 38404 11649 38422
rect 11649 38404 11655 38422
rect 11537 38338 11543 38390
rect 11543 38338 11589 38390
rect 11603 38338 11649 38390
rect 11649 38338 11655 38390
rect 11537 38271 11543 38323
rect 11543 38271 11589 38323
rect 11603 38271 11649 38323
rect 11649 38271 11655 38323
rect 11537 38204 11543 38256
rect 11543 38204 11589 38256
rect 11603 38204 11649 38256
rect 11649 38204 11655 38256
rect 11537 36714 11589 36720
rect 11537 36680 11543 36714
rect 11543 36680 11577 36714
rect 11577 36680 11589 36714
rect 11537 36668 11589 36680
rect 11603 36714 11655 36720
rect 11603 36680 11615 36714
rect 11615 36680 11649 36714
rect 11649 36680 11655 36714
rect 11603 36668 11655 36680
rect 11537 36641 11589 36654
rect 11537 36607 11543 36641
rect 11543 36607 11577 36641
rect 11577 36607 11589 36641
rect 11537 36602 11589 36607
rect 11603 36641 11655 36654
rect 11603 36607 11615 36641
rect 11615 36607 11649 36641
rect 11649 36607 11655 36641
rect 11603 36602 11655 36607
rect 11537 36568 11589 36588
rect 11537 36536 11543 36568
rect 11543 36536 11577 36568
rect 11577 36536 11589 36568
rect 11603 36568 11655 36588
rect 11603 36536 11615 36568
rect 11615 36536 11649 36568
rect 11649 36536 11655 36568
rect 11537 36495 11589 36522
rect 11537 36470 11543 36495
rect 11543 36470 11577 36495
rect 11577 36470 11589 36495
rect 11603 36495 11655 36522
rect 11603 36470 11615 36495
rect 11615 36470 11649 36495
rect 11649 36470 11655 36495
rect 11537 36422 11589 36456
rect 11603 36422 11655 36456
rect 11537 36404 11543 36422
rect 11543 36404 11589 36422
rect 11603 36404 11649 36422
rect 11649 36404 11655 36422
rect 11537 36338 11543 36390
rect 11543 36338 11589 36390
rect 11603 36338 11649 36390
rect 11649 36338 11655 36390
rect 11537 36271 11543 36323
rect 11543 36271 11589 36323
rect 11603 36271 11649 36323
rect 11649 36271 11655 36323
rect 11537 36204 11543 36256
rect 11543 36204 11589 36256
rect 11603 36204 11649 36256
rect 11649 36204 11655 36256
rect 11814 37840 11820 37892
rect 11820 37840 11866 37892
rect 11880 37840 11926 37892
rect 11926 37840 11932 37892
rect 11814 37773 11820 37825
rect 11820 37773 11866 37825
rect 11880 37773 11926 37825
rect 11926 37773 11932 37825
rect 11814 37706 11820 37758
rect 11820 37706 11866 37758
rect 11880 37706 11926 37758
rect 11926 37706 11932 37758
rect 11814 37639 11820 37691
rect 11820 37639 11866 37691
rect 11880 37639 11926 37691
rect 11926 37639 11932 37691
rect 11814 37572 11820 37624
rect 11820 37572 11866 37624
rect 11880 37572 11926 37624
rect 11926 37572 11932 37624
rect 11814 37505 11820 37557
rect 11820 37505 11866 37557
rect 11880 37505 11926 37557
rect 11926 37505 11932 37557
rect 11814 37438 11820 37490
rect 11820 37438 11866 37490
rect 11880 37438 11926 37490
rect 11926 37438 11932 37490
rect 11814 37380 11820 37423
rect 11820 37380 11866 37423
rect 11880 37380 11926 37423
rect 11926 37380 11932 37423
rect 11814 37371 11866 37380
rect 11880 37371 11932 37380
rect 11814 37304 11866 37356
rect 11880 37304 11932 37356
rect 11814 37237 11866 37289
rect 11880 37237 11932 37289
rect 11814 37170 11866 37222
rect 11880 37170 11932 37222
rect 11814 37103 11866 37155
rect 11880 37103 11932 37155
rect 11814 37036 11866 37088
rect 11880 37036 11932 37088
rect 11814 35840 11820 35892
rect 11820 35840 11866 35892
rect 11880 35840 11926 35892
rect 11926 35840 11932 35892
rect 11814 35774 11820 35826
rect 11820 35774 11866 35826
rect 11880 35774 11926 35826
rect 11926 35774 11932 35826
rect 11814 35708 11820 35760
rect 11820 35708 11866 35760
rect 11880 35708 11926 35760
rect 11926 35708 11932 35760
rect 11814 35642 11820 35694
rect 11820 35642 11866 35694
rect 11880 35642 11926 35694
rect 11926 35642 11932 35694
rect 11814 35575 11820 35627
rect 11820 35575 11866 35627
rect 11880 35575 11926 35627
rect 11926 35575 11932 35627
rect 11814 35508 11820 35560
rect 11820 35508 11866 35560
rect 11880 35508 11926 35560
rect 11926 35508 11932 35560
rect 11814 35441 11820 35493
rect 11820 35441 11866 35493
rect 11880 35441 11926 35493
rect 11926 35441 11932 35493
rect 11814 35380 11820 35426
rect 11820 35380 11866 35426
rect 11880 35380 11926 35426
rect 11926 35380 11932 35426
rect 11814 35374 11866 35380
rect 11880 35374 11932 35380
rect 12091 38714 12143 38720
rect 12091 38680 12097 38714
rect 12097 38680 12131 38714
rect 12131 38680 12143 38714
rect 12091 38668 12143 38680
rect 12157 38714 12209 38720
rect 12157 38680 12169 38714
rect 12169 38680 12203 38714
rect 12203 38680 12209 38714
rect 12157 38668 12209 38680
rect 12091 38641 12143 38654
rect 12091 38607 12097 38641
rect 12097 38607 12131 38641
rect 12131 38607 12143 38641
rect 12091 38602 12143 38607
rect 12157 38641 12209 38654
rect 12157 38607 12169 38641
rect 12169 38607 12203 38641
rect 12203 38607 12209 38641
rect 12157 38602 12209 38607
rect 12091 38568 12143 38588
rect 12091 38536 12097 38568
rect 12097 38536 12131 38568
rect 12131 38536 12143 38568
rect 12157 38568 12209 38588
rect 12157 38536 12169 38568
rect 12169 38536 12203 38568
rect 12203 38536 12209 38568
rect 12091 38495 12143 38522
rect 12091 38470 12097 38495
rect 12097 38470 12131 38495
rect 12131 38470 12143 38495
rect 12157 38495 12209 38522
rect 12157 38470 12169 38495
rect 12169 38470 12203 38495
rect 12203 38470 12209 38495
rect 12091 38422 12143 38456
rect 12157 38422 12209 38456
rect 12091 38404 12097 38422
rect 12097 38404 12143 38422
rect 12157 38404 12203 38422
rect 12203 38404 12209 38422
rect 12091 38338 12097 38390
rect 12097 38338 12143 38390
rect 12157 38338 12203 38390
rect 12203 38338 12209 38390
rect 12091 38271 12097 38323
rect 12097 38271 12143 38323
rect 12157 38271 12203 38323
rect 12203 38271 12209 38323
rect 12091 38204 12097 38256
rect 12097 38204 12143 38256
rect 12157 38204 12203 38256
rect 12203 38204 12209 38256
rect 12091 36714 12143 36720
rect 12091 36680 12097 36714
rect 12097 36680 12131 36714
rect 12131 36680 12143 36714
rect 12091 36668 12143 36680
rect 12157 36714 12209 36720
rect 12157 36680 12169 36714
rect 12169 36680 12203 36714
rect 12203 36680 12209 36714
rect 12157 36668 12209 36680
rect 12091 36641 12143 36654
rect 12091 36607 12097 36641
rect 12097 36607 12131 36641
rect 12131 36607 12143 36641
rect 12091 36602 12143 36607
rect 12157 36641 12209 36654
rect 12157 36607 12169 36641
rect 12169 36607 12203 36641
rect 12203 36607 12209 36641
rect 12157 36602 12209 36607
rect 12091 36568 12143 36588
rect 12091 36536 12097 36568
rect 12097 36536 12131 36568
rect 12131 36536 12143 36568
rect 12157 36568 12209 36588
rect 12157 36536 12169 36568
rect 12169 36536 12203 36568
rect 12203 36536 12209 36568
rect 12091 36495 12143 36522
rect 12091 36470 12097 36495
rect 12097 36470 12131 36495
rect 12131 36470 12143 36495
rect 12157 36495 12209 36522
rect 12157 36470 12169 36495
rect 12169 36470 12203 36495
rect 12203 36470 12209 36495
rect 12091 36422 12143 36456
rect 12157 36422 12209 36456
rect 12091 36404 12097 36422
rect 12097 36404 12143 36422
rect 12157 36404 12203 36422
rect 12203 36404 12209 36422
rect 12091 36338 12097 36390
rect 12097 36338 12143 36390
rect 12157 36338 12203 36390
rect 12203 36338 12209 36390
rect 12091 36271 12097 36323
rect 12097 36271 12143 36323
rect 12157 36271 12203 36323
rect 12203 36271 12209 36323
rect 12091 36204 12097 36256
rect 12097 36204 12143 36256
rect 12157 36204 12203 36256
rect 12203 36204 12209 36256
rect 12368 37840 12374 37892
rect 12374 37840 12420 37892
rect 12434 37840 12480 37892
rect 12480 37840 12486 37892
rect 12368 37773 12374 37825
rect 12374 37773 12420 37825
rect 12434 37773 12480 37825
rect 12480 37773 12486 37825
rect 12368 37706 12374 37758
rect 12374 37706 12420 37758
rect 12434 37706 12480 37758
rect 12480 37706 12486 37758
rect 12368 37639 12374 37691
rect 12374 37639 12420 37691
rect 12434 37639 12480 37691
rect 12480 37639 12486 37691
rect 12368 37572 12374 37624
rect 12374 37572 12420 37624
rect 12434 37572 12480 37624
rect 12480 37572 12486 37624
rect 12368 37505 12374 37557
rect 12374 37505 12420 37557
rect 12434 37505 12480 37557
rect 12480 37505 12486 37557
rect 12368 37438 12374 37490
rect 12374 37438 12420 37490
rect 12434 37438 12480 37490
rect 12480 37438 12486 37490
rect 12368 37380 12374 37423
rect 12374 37380 12420 37423
rect 12434 37380 12480 37423
rect 12480 37380 12486 37423
rect 12368 37371 12420 37380
rect 12434 37371 12486 37380
rect 12368 37304 12420 37356
rect 12434 37304 12486 37356
rect 12368 37237 12420 37289
rect 12434 37237 12486 37289
rect 12368 37170 12420 37222
rect 12434 37170 12486 37222
rect 12368 37103 12420 37155
rect 12434 37103 12486 37155
rect 12368 37036 12420 37088
rect 12434 37036 12486 37088
rect 12368 35840 12374 35892
rect 12374 35840 12420 35892
rect 12434 35840 12480 35892
rect 12480 35840 12486 35892
rect 12368 35774 12374 35826
rect 12374 35774 12420 35826
rect 12434 35774 12480 35826
rect 12480 35774 12486 35826
rect 12368 35708 12374 35760
rect 12374 35708 12420 35760
rect 12434 35708 12480 35760
rect 12480 35708 12486 35760
rect 12368 35642 12374 35694
rect 12374 35642 12420 35694
rect 12434 35642 12480 35694
rect 12480 35642 12486 35694
rect 12368 35575 12374 35627
rect 12374 35575 12420 35627
rect 12434 35575 12480 35627
rect 12480 35575 12486 35627
rect 12368 35508 12374 35560
rect 12374 35508 12420 35560
rect 12434 35508 12480 35560
rect 12480 35508 12486 35560
rect 12368 35441 12374 35493
rect 12374 35441 12420 35493
rect 12434 35441 12480 35493
rect 12480 35441 12486 35493
rect 12368 35380 12374 35426
rect 12374 35380 12420 35426
rect 12434 35380 12480 35426
rect 12480 35380 12486 35426
rect 12368 35374 12420 35380
rect 12434 35374 12486 35380
rect 12645 38714 12697 38720
rect 12645 38680 12651 38714
rect 12651 38680 12685 38714
rect 12685 38680 12697 38714
rect 12645 38668 12697 38680
rect 12711 38714 12763 38720
rect 12711 38680 12723 38714
rect 12723 38680 12757 38714
rect 12757 38680 12763 38714
rect 12711 38668 12763 38680
rect 12645 38641 12697 38654
rect 12645 38607 12651 38641
rect 12651 38607 12685 38641
rect 12685 38607 12697 38641
rect 12645 38602 12697 38607
rect 12711 38641 12763 38654
rect 12711 38607 12723 38641
rect 12723 38607 12757 38641
rect 12757 38607 12763 38641
rect 12711 38602 12763 38607
rect 12645 38568 12697 38588
rect 12645 38536 12651 38568
rect 12651 38536 12685 38568
rect 12685 38536 12697 38568
rect 12711 38568 12763 38588
rect 12711 38536 12723 38568
rect 12723 38536 12757 38568
rect 12757 38536 12763 38568
rect 12645 38495 12697 38522
rect 12645 38470 12651 38495
rect 12651 38470 12685 38495
rect 12685 38470 12697 38495
rect 12711 38495 12763 38522
rect 12711 38470 12723 38495
rect 12723 38470 12757 38495
rect 12757 38470 12763 38495
rect 12645 38422 12697 38456
rect 12711 38422 12763 38456
rect 12645 38404 12651 38422
rect 12651 38404 12697 38422
rect 12711 38404 12757 38422
rect 12757 38404 12763 38422
rect 12645 38338 12651 38390
rect 12651 38338 12697 38390
rect 12711 38338 12757 38390
rect 12757 38338 12763 38390
rect 12645 38271 12651 38323
rect 12651 38271 12697 38323
rect 12711 38271 12757 38323
rect 12757 38271 12763 38323
rect 12645 38204 12651 38256
rect 12651 38204 12697 38256
rect 12711 38204 12757 38256
rect 12757 38204 12763 38256
rect 12645 36714 12697 36720
rect 12645 36680 12651 36714
rect 12651 36680 12685 36714
rect 12685 36680 12697 36714
rect 12645 36668 12697 36680
rect 12711 36714 12763 36720
rect 12711 36680 12723 36714
rect 12723 36680 12757 36714
rect 12757 36680 12763 36714
rect 12711 36668 12763 36680
rect 12645 36641 12697 36654
rect 12645 36607 12651 36641
rect 12651 36607 12685 36641
rect 12685 36607 12697 36641
rect 12645 36602 12697 36607
rect 12711 36641 12763 36654
rect 12711 36607 12723 36641
rect 12723 36607 12757 36641
rect 12757 36607 12763 36641
rect 12711 36602 12763 36607
rect 12645 36568 12697 36588
rect 12645 36536 12651 36568
rect 12651 36536 12685 36568
rect 12685 36536 12697 36568
rect 12711 36568 12763 36588
rect 12711 36536 12723 36568
rect 12723 36536 12757 36568
rect 12757 36536 12763 36568
rect 12645 36495 12697 36522
rect 12645 36470 12651 36495
rect 12651 36470 12685 36495
rect 12685 36470 12697 36495
rect 12711 36495 12763 36522
rect 12711 36470 12723 36495
rect 12723 36470 12757 36495
rect 12757 36470 12763 36495
rect 12645 36422 12697 36456
rect 12711 36422 12763 36456
rect 12645 36404 12651 36422
rect 12651 36404 12697 36422
rect 12711 36404 12757 36422
rect 12757 36404 12763 36422
rect 12645 36338 12651 36390
rect 12651 36338 12697 36390
rect 12711 36338 12757 36390
rect 12757 36338 12763 36390
rect 12645 36271 12651 36323
rect 12651 36271 12697 36323
rect 12711 36271 12757 36323
rect 12757 36271 12763 36323
rect 12645 36204 12651 36256
rect 12651 36204 12697 36256
rect 12711 36204 12757 36256
rect 12757 36204 12763 36256
rect 12922 37840 12928 37892
rect 12928 37840 12974 37892
rect 12988 37840 13034 37892
rect 13034 37840 13040 37892
rect 12922 37773 12928 37825
rect 12928 37773 12974 37825
rect 12988 37773 13034 37825
rect 13034 37773 13040 37825
rect 12922 37706 12928 37758
rect 12928 37706 12974 37758
rect 12988 37706 13034 37758
rect 13034 37706 13040 37758
rect 12922 37639 12928 37691
rect 12928 37639 12974 37691
rect 12988 37639 13034 37691
rect 13034 37639 13040 37691
rect 12922 37572 12928 37624
rect 12928 37572 12974 37624
rect 12988 37572 13034 37624
rect 13034 37572 13040 37624
rect 12922 37505 12928 37557
rect 12928 37505 12974 37557
rect 12988 37505 13034 37557
rect 13034 37505 13040 37557
rect 12922 37438 12928 37490
rect 12928 37438 12974 37490
rect 12988 37438 13034 37490
rect 13034 37438 13040 37490
rect 12922 37380 12928 37423
rect 12928 37380 12974 37423
rect 12988 37380 13034 37423
rect 13034 37380 13040 37423
rect 12922 37371 12974 37380
rect 12988 37371 13040 37380
rect 12922 37304 12974 37356
rect 12988 37304 13040 37356
rect 12922 37237 12974 37289
rect 12988 37237 13040 37289
rect 12922 37170 12974 37222
rect 12988 37170 13040 37222
rect 12922 37103 12974 37155
rect 12988 37103 13040 37155
rect 12922 37036 12974 37088
rect 12988 37036 13040 37088
rect 12922 35840 12928 35892
rect 12928 35840 12974 35892
rect 12988 35840 13034 35892
rect 13034 35840 13040 35892
rect 12922 35774 12928 35826
rect 12928 35774 12974 35826
rect 12988 35774 13034 35826
rect 13034 35774 13040 35826
rect 12922 35708 12928 35760
rect 12928 35708 12974 35760
rect 12988 35708 13034 35760
rect 13034 35708 13040 35760
rect 12922 35642 12928 35694
rect 12928 35642 12974 35694
rect 12988 35642 13034 35694
rect 13034 35642 13040 35694
rect 12922 35575 12928 35627
rect 12928 35575 12974 35627
rect 12988 35575 13034 35627
rect 13034 35575 13040 35627
rect 12922 35508 12928 35560
rect 12928 35508 12974 35560
rect 12988 35508 13034 35560
rect 13034 35508 13040 35560
rect 12922 35441 12928 35493
rect 12928 35441 12974 35493
rect 12988 35441 13034 35493
rect 13034 35441 13040 35493
rect 12922 35380 12928 35426
rect 12928 35380 12974 35426
rect 12988 35380 13034 35426
rect 13034 35380 13040 35426
rect 12922 35374 12974 35380
rect 12988 35374 13040 35380
rect 13200 38714 13252 38720
rect 13200 38680 13205 38714
rect 13205 38680 13239 38714
rect 13239 38680 13252 38714
rect 13200 38668 13252 38680
rect 13270 38714 13322 38720
rect 13270 38680 13277 38714
rect 13277 38680 13311 38714
rect 13311 38680 13322 38714
rect 13270 38668 13322 38680
rect 13340 38668 13392 38720
rect 13410 38668 13462 38720
rect 13480 38668 13521 38720
rect 13521 38668 13532 38720
rect 13550 38668 13602 38720
rect 13200 38641 13252 38654
rect 13200 38607 13205 38641
rect 13205 38607 13239 38641
rect 13239 38607 13252 38641
rect 13200 38602 13252 38607
rect 13270 38641 13322 38654
rect 13270 38607 13277 38641
rect 13277 38607 13311 38641
rect 13311 38607 13322 38641
rect 13270 38602 13322 38607
rect 13340 38602 13392 38654
rect 13410 38602 13462 38654
rect 13480 38602 13521 38654
rect 13521 38602 13532 38654
rect 13550 38602 13602 38654
rect 13200 38568 13252 38588
rect 13200 38536 13205 38568
rect 13205 38536 13239 38568
rect 13239 38536 13252 38568
rect 13270 38568 13322 38588
rect 13270 38536 13277 38568
rect 13277 38536 13311 38568
rect 13311 38536 13322 38568
rect 13340 38536 13392 38588
rect 13410 38536 13462 38588
rect 13480 38536 13521 38588
rect 13521 38536 13532 38588
rect 13550 38536 13602 38588
rect 13200 38495 13252 38522
rect 13200 38470 13205 38495
rect 13205 38470 13239 38495
rect 13239 38470 13252 38495
rect 13270 38495 13322 38522
rect 13270 38470 13277 38495
rect 13277 38470 13311 38495
rect 13311 38470 13322 38495
rect 13340 38470 13392 38522
rect 13410 38470 13462 38522
rect 13480 38470 13521 38522
rect 13521 38470 13532 38522
rect 13550 38470 13602 38522
rect 13200 38422 13252 38456
rect 13270 38422 13322 38456
rect 13200 38404 13205 38422
rect 13205 38404 13252 38422
rect 13270 38404 13311 38422
rect 13311 38404 13322 38422
rect 13340 38404 13392 38456
rect 13410 38404 13462 38456
rect 13480 38404 13521 38456
rect 13521 38404 13532 38456
rect 13550 38404 13602 38456
rect 13200 38338 13205 38390
rect 13205 38338 13252 38390
rect 13270 38338 13311 38390
rect 13311 38338 13322 38390
rect 13340 38338 13392 38390
rect 13410 38338 13462 38390
rect 13480 38338 13521 38390
rect 13521 38338 13532 38390
rect 13550 38338 13602 38390
rect 13200 38271 13205 38323
rect 13205 38271 13252 38323
rect 13270 38271 13311 38323
rect 13311 38271 13322 38323
rect 13340 38271 13392 38323
rect 13410 38271 13462 38323
rect 13480 38271 13521 38323
rect 13521 38271 13532 38323
rect 13550 38271 13602 38323
rect 13200 38204 13205 38256
rect 13205 38204 13252 38256
rect 13270 38204 13311 38256
rect 13311 38204 13322 38256
rect 13340 38204 13392 38256
rect 13410 38204 13462 38256
rect 13480 38204 13521 38256
rect 13521 38204 13532 38256
rect 13550 38204 13602 38256
rect 13200 36714 13252 36720
rect 13200 36680 13205 36714
rect 13205 36680 13239 36714
rect 13239 36680 13252 36714
rect 13200 36668 13252 36680
rect 13270 36714 13322 36720
rect 13270 36680 13277 36714
rect 13277 36680 13311 36714
rect 13311 36680 13322 36714
rect 13270 36668 13322 36680
rect 13340 36668 13392 36720
rect 13410 36668 13462 36720
rect 13480 36668 13521 36720
rect 13521 36668 13532 36720
rect 13550 36668 13602 36720
rect 13200 36641 13252 36654
rect 13200 36607 13205 36641
rect 13205 36607 13239 36641
rect 13239 36607 13252 36641
rect 13200 36602 13252 36607
rect 13270 36641 13322 36654
rect 13270 36607 13277 36641
rect 13277 36607 13311 36641
rect 13311 36607 13322 36641
rect 13270 36602 13322 36607
rect 13340 36602 13392 36654
rect 13410 36602 13462 36654
rect 13480 36602 13521 36654
rect 13521 36602 13532 36654
rect 13550 36602 13602 36654
rect 13200 36568 13252 36588
rect 13200 36536 13205 36568
rect 13205 36536 13239 36568
rect 13239 36536 13252 36568
rect 13270 36568 13322 36588
rect 13270 36536 13277 36568
rect 13277 36536 13311 36568
rect 13311 36536 13322 36568
rect 13340 36536 13392 36588
rect 13410 36536 13462 36588
rect 13480 36536 13521 36588
rect 13521 36536 13532 36588
rect 13550 36536 13602 36588
rect 13200 36495 13252 36522
rect 13200 36470 13205 36495
rect 13205 36470 13239 36495
rect 13239 36470 13252 36495
rect 13270 36495 13322 36522
rect 13270 36470 13277 36495
rect 13277 36470 13311 36495
rect 13311 36470 13322 36495
rect 13340 36470 13392 36522
rect 13410 36470 13462 36522
rect 13480 36470 13521 36522
rect 13521 36470 13532 36522
rect 13550 36470 13602 36522
rect 13200 36422 13252 36456
rect 13270 36422 13322 36456
rect 13200 36404 13205 36422
rect 13205 36404 13252 36422
rect 13270 36404 13311 36422
rect 13311 36404 13322 36422
rect 13340 36404 13392 36456
rect 13410 36404 13462 36456
rect 13480 36404 13521 36456
rect 13521 36404 13532 36456
rect 13550 36404 13602 36456
rect 13200 36338 13205 36390
rect 13205 36338 13252 36390
rect 13270 36338 13311 36390
rect 13311 36338 13322 36390
rect 13340 36338 13392 36390
rect 13410 36338 13462 36390
rect 13480 36338 13521 36390
rect 13521 36338 13532 36390
rect 13550 36338 13602 36390
rect 13200 36271 13205 36323
rect 13205 36271 13252 36323
rect 13270 36271 13311 36323
rect 13311 36271 13322 36323
rect 13340 36271 13392 36323
rect 13410 36271 13462 36323
rect 13480 36271 13521 36323
rect 13521 36271 13532 36323
rect 13550 36271 13602 36323
rect 13200 36204 13205 36256
rect 13205 36204 13252 36256
rect 13270 36204 13311 36256
rect 13311 36204 13322 36256
rect 13340 36204 13392 36256
rect 13410 36204 13462 36256
rect 13480 36204 13521 36256
rect 13521 36204 13532 36256
rect 13550 36204 13602 36256
rect 3167 34714 3219 34720
rect 3167 34680 3173 34714
rect 3173 34680 3207 34714
rect 3207 34680 3219 34714
rect 3167 34668 3219 34680
rect 3233 34714 3285 34720
rect 3233 34680 3245 34714
rect 3245 34680 3279 34714
rect 3279 34680 3285 34714
rect 3233 34668 3285 34680
rect 3167 34641 3219 34654
rect 3167 34607 3173 34641
rect 3173 34607 3207 34641
rect 3207 34607 3219 34641
rect 3167 34602 3219 34607
rect 3233 34641 3285 34654
rect 3233 34607 3245 34641
rect 3245 34607 3279 34641
rect 3279 34607 3285 34641
rect 3233 34602 3285 34607
rect 3167 34568 3219 34588
rect 3167 34536 3173 34568
rect 3173 34536 3207 34568
rect 3207 34536 3219 34568
rect 3233 34568 3285 34588
rect 3233 34536 3245 34568
rect 3245 34536 3279 34568
rect 3279 34536 3285 34568
rect 3167 34495 3219 34522
rect 3167 34470 3173 34495
rect 3173 34470 3207 34495
rect 3207 34470 3219 34495
rect 3233 34495 3285 34522
rect 3233 34470 3245 34495
rect 3245 34470 3279 34495
rect 3279 34470 3285 34495
rect 3167 34422 3219 34456
rect 3233 34422 3285 34456
rect 3167 34404 3173 34422
rect 3173 34404 3219 34422
rect 3233 34404 3279 34422
rect 3279 34404 3285 34422
rect 3167 34338 3173 34390
rect 3173 34338 3219 34390
rect 3233 34338 3279 34390
rect 3279 34338 3285 34390
rect 3167 34271 3173 34323
rect 3173 34271 3219 34323
rect 3233 34271 3279 34323
rect 3279 34271 3285 34323
rect 3167 34204 3173 34256
rect 3173 34204 3219 34256
rect 3233 34204 3279 34256
rect 3279 34204 3285 34256
rect 3167 32714 3219 32720
rect 3167 32680 3173 32714
rect 3173 32680 3207 32714
rect 3207 32680 3219 32714
rect 3167 32668 3219 32680
rect 3233 32714 3285 32720
rect 3233 32680 3245 32714
rect 3245 32680 3279 32714
rect 3279 32680 3285 32714
rect 3233 32668 3285 32680
rect 3167 32641 3219 32654
rect 3167 32607 3173 32641
rect 3173 32607 3207 32641
rect 3207 32607 3219 32641
rect 3167 32602 3219 32607
rect 3233 32641 3285 32654
rect 3233 32607 3245 32641
rect 3245 32607 3279 32641
rect 3279 32607 3285 32641
rect 3233 32602 3285 32607
rect 3167 32568 3219 32588
rect 3167 32536 3173 32568
rect 3173 32536 3207 32568
rect 3207 32536 3219 32568
rect 3233 32568 3285 32588
rect 3233 32536 3245 32568
rect 3245 32536 3279 32568
rect 3279 32536 3285 32568
rect 3167 32495 3219 32522
rect 3167 32470 3173 32495
rect 3173 32470 3207 32495
rect 3207 32470 3219 32495
rect 3233 32495 3285 32522
rect 3233 32470 3245 32495
rect 3245 32470 3279 32495
rect 3279 32470 3285 32495
rect 3167 32422 3219 32456
rect 3233 32422 3285 32456
rect 3167 32404 3173 32422
rect 3173 32404 3219 32422
rect 3233 32404 3279 32422
rect 3279 32404 3285 32422
rect 3167 32338 3173 32390
rect 3173 32338 3219 32390
rect 3233 32338 3279 32390
rect 3279 32338 3285 32390
rect 3167 32271 3173 32323
rect 3173 32271 3219 32323
rect 3233 32271 3279 32323
rect 3279 32271 3285 32323
rect 3167 32204 3173 32256
rect 3173 32204 3219 32256
rect 3233 32204 3279 32256
rect 3279 32204 3285 32256
rect 3167 30714 3219 30720
rect 3167 30680 3173 30714
rect 3173 30680 3207 30714
rect 3207 30680 3219 30714
rect 3167 30668 3219 30680
rect 3233 30714 3285 30720
rect 3233 30680 3245 30714
rect 3245 30680 3279 30714
rect 3279 30680 3285 30714
rect 3233 30668 3285 30680
rect 3167 30641 3219 30654
rect 3167 30607 3173 30641
rect 3173 30607 3207 30641
rect 3207 30607 3219 30641
rect 3167 30602 3219 30607
rect 3233 30641 3285 30654
rect 3233 30607 3245 30641
rect 3245 30607 3279 30641
rect 3279 30607 3285 30641
rect 3233 30602 3285 30607
rect 3167 30568 3219 30588
rect 3167 30536 3173 30568
rect 3173 30536 3207 30568
rect 3207 30536 3219 30568
rect 3233 30568 3285 30588
rect 3233 30536 3245 30568
rect 3245 30536 3279 30568
rect 3279 30536 3285 30568
rect 3167 30495 3219 30522
rect 3167 30470 3173 30495
rect 3173 30470 3207 30495
rect 3207 30470 3219 30495
rect 3233 30495 3285 30522
rect 3233 30470 3245 30495
rect 3245 30470 3279 30495
rect 3279 30470 3285 30495
rect 3167 30422 3219 30456
rect 3233 30422 3285 30456
rect 3167 30404 3173 30422
rect 3173 30404 3219 30422
rect 3233 30404 3279 30422
rect 3279 30404 3285 30422
rect 3167 30338 3173 30390
rect 3173 30338 3219 30390
rect 3233 30338 3279 30390
rect 3279 30338 3285 30390
rect 3167 30271 3173 30323
rect 3173 30271 3219 30323
rect 3233 30271 3279 30323
rect 3279 30271 3285 30323
rect 3167 30204 3173 30256
rect 3173 30204 3219 30256
rect 3233 30204 3279 30256
rect 3279 30204 3285 30256
rect 3585 33840 3591 33892
rect 3591 33840 3637 33892
rect 3651 33840 3697 33892
rect 3697 33840 3703 33892
rect 3585 33774 3591 33826
rect 3591 33774 3637 33826
rect 3651 33774 3697 33826
rect 3697 33774 3703 33826
rect 3585 33708 3591 33760
rect 3591 33708 3637 33760
rect 3651 33708 3697 33760
rect 3697 33708 3703 33760
rect 3585 33642 3591 33694
rect 3591 33642 3637 33694
rect 3651 33642 3697 33694
rect 3697 33642 3703 33694
rect 3585 33575 3591 33627
rect 3591 33575 3637 33627
rect 3651 33575 3697 33627
rect 3697 33575 3703 33627
rect 3585 33508 3591 33560
rect 3591 33508 3637 33560
rect 3651 33508 3697 33560
rect 3697 33508 3703 33560
rect 3585 33441 3591 33493
rect 3591 33441 3637 33493
rect 3651 33441 3697 33493
rect 3697 33441 3703 33493
rect 3585 33380 3591 33426
rect 3591 33380 3637 33426
rect 3651 33380 3697 33426
rect 3697 33380 3703 33426
rect 3585 33374 3637 33380
rect 3651 33374 3703 33380
rect 3585 31840 3591 31892
rect 3591 31840 3637 31892
rect 3651 31840 3697 31892
rect 3697 31840 3703 31892
rect 3585 31774 3591 31826
rect 3591 31774 3637 31826
rect 3651 31774 3697 31826
rect 3697 31774 3703 31826
rect 3585 31708 3591 31760
rect 3591 31708 3637 31760
rect 3651 31708 3697 31760
rect 3697 31708 3703 31760
rect 3585 31642 3591 31694
rect 3591 31642 3637 31694
rect 3651 31642 3697 31694
rect 3697 31642 3703 31694
rect 3585 31575 3591 31627
rect 3591 31575 3637 31627
rect 3651 31575 3697 31627
rect 3697 31575 3703 31627
rect 3585 31508 3591 31560
rect 3591 31508 3637 31560
rect 3651 31508 3697 31560
rect 3697 31508 3703 31560
rect 3585 31441 3591 31493
rect 3591 31441 3637 31493
rect 3651 31441 3697 31493
rect 3697 31441 3703 31493
rect 3585 31380 3591 31426
rect 3591 31380 3637 31426
rect 3651 31380 3697 31426
rect 3697 31380 3703 31426
rect 3585 31374 3637 31380
rect 3651 31374 3703 31380
rect 3585 29840 3591 29892
rect 3591 29840 3637 29892
rect 3651 29840 3697 29892
rect 3697 29840 3703 29892
rect 3585 29774 3591 29826
rect 3591 29774 3637 29826
rect 3651 29774 3697 29826
rect 3697 29774 3703 29826
rect 3585 29708 3591 29760
rect 3591 29708 3637 29760
rect 3651 29708 3697 29760
rect 3697 29708 3703 29760
rect 3585 29642 3591 29694
rect 3591 29642 3637 29694
rect 3651 29642 3697 29694
rect 3697 29642 3703 29694
rect 3585 29575 3591 29627
rect 3591 29575 3637 29627
rect 3651 29575 3697 29627
rect 3697 29575 3703 29627
rect 3585 29508 3591 29560
rect 3591 29508 3637 29560
rect 3651 29508 3697 29560
rect 3697 29508 3703 29560
rect 3585 29441 3591 29493
rect 3591 29441 3637 29493
rect 3651 29441 3697 29493
rect 3697 29441 3703 29493
rect 3585 29380 3591 29426
rect 3591 29380 3637 29426
rect 3651 29380 3697 29426
rect 3697 29380 3703 29426
rect 3585 29374 3637 29380
rect 3651 29374 3703 29380
rect 4003 34714 4055 34720
rect 4003 34680 4009 34714
rect 4009 34680 4043 34714
rect 4043 34680 4055 34714
rect 4003 34668 4055 34680
rect 4069 34714 4121 34720
rect 4069 34680 4081 34714
rect 4081 34680 4115 34714
rect 4115 34680 4121 34714
rect 4069 34668 4121 34680
rect 4003 34641 4055 34654
rect 4003 34607 4009 34641
rect 4009 34607 4043 34641
rect 4043 34607 4055 34641
rect 4003 34602 4055 34607
rect 4069 34641 4121 34654
rect 4069 34607 4081 34641
rect 4081 34607 4115 34641
rect 4115 34607 4121 34641
rect 4069 34602 4121 34607
rect 4003 34568 4055 34588
rect 4003 34536 4009 34568
rect 4009 34536 4043 34568
rect 4043 34536 4055 34568
rect 4069 34568 4121 34588
rect 4069 34536 4081 34568
rect 4081 34536 4115 34568
rect 4115 34536 4121 34568
rect 4003 34495 4055 34522
rect 4003 34470 4009 34495
rect 4009 34470 4043 34495
rect 4043 34470 4055 34495
rect 4069 34495 4121 34522
rect 4069 34470 4081 34495
rect 4081 34470 4115 34495
rect 4115 34470 4121 34495
rect 4003 34422 4055 34456
rect 4069 34422 4121 34456
rect 4003 34404 4009 34422
rect 4009 34404 4055 34422
rect 4069 34404 4115 34422
rect 4115 34404 4121 34422
rect 4003 34338 4009 34390
rect 4009 34338 4055 34390
rect 4069 34338 4115 34390
rect 4115 34338 4121 34390
rect 4003 34271 4009 34323
rect 4009 34271 4055 34323
rect 4069 34271 4115 34323
rect 4115 34271 4121 34323
rect 4003 34204 4009 34256
rect 4009 34204 4055 34256
rect 4069 34204 4115 34256
rect 4115 34204 4121 34256
rect 4003 32714 4055 32720
rect 4003 32680 4009 32714
rect 4009 32680 4043 32714
rect 4043 32680 4055 32714
rect 4003 32668 4055 32680
rect 4069 32714 4121 32720
rect 4069 32680 4081 32714
rect 4081 32680 4115 32714
rect 4115 32680 4121 32714
rect 4069 32668 4121 32680
rect 4003 32641 4055 32654
rect 4003 32607 4009 32641
rect 4009 32607 4043 32641
rect 4043 32607 4055 32641
rect 4003 32602 4055 32607
rect 4069 32641 4121 32654
rect 4069 32607 4081 32641
rect 4081 32607 4115 32641
rect 4115 32607 4121 32641
rect 4069 32602 4121 32607
rect 4003 32568 4055 32588
rect 4003 32536 4009 32568
rect 4009 32536 4043 32568
rect 4043 32536 4055 32568
rect 4069 32568 4121 32588
rect 4069 32536 4081 32568
rect 4081 32536 4115 32568
rect 4115 32536 4121 32568
rect 4003 32495 4055 32522
rect 4003 32470 4009 32495
rect 4009 32470 4043 32495
rect 4043 32470 4055 32495
rect 4069 32495 4121 32522
rect 4069 32470 4081 32495
rect 4081 32470 4115 32495
rect 4115 32470 4121 32495
rect 4003 32422 4055 32456
rect 4069 32422 4121 32456
rect 4003 32404 4009 32422
rect 4009 32404 4055 32422
rect 4069 32404 4115 32422
rect 4115 32404 4121 32422
rect 4003 32338 4009 32390
rect 4009 32338 4055 32390
rect 4069 32338 4115 32390
rect 4115 32338 4121 32390
rect 4003 32271 4009 32323
rect 4009 32271 4055 32323
rect 4069 32271 4115 32323
rect 4115 32271 4121 32323
rect 4003 32204 4009 32256
rect 4009 32204 4055 32256
rect 4069 32204 4115 32256
rect 4115 32204 4121 32256
rect 4003 30714 4055 30720
rect 4003 30680 4009 30714
rect 4009 30680 4043 30714
rect 4043 30680 4055 30714
rect 4003 30668 4055 30680
rect 4069 30714 4121 30720
rect 4069 30680 4081 30714
rect 4081 30680 4115 30714
rect 4115 30680 4121 30714
rect 4069 30668 4121 30680
rect 4003 30641 4055 30654
rect 4003 30607 4009 30641
rect 4009 30607 4043 30641
rect 4043 30607 4055 30641
rect 4003 30602 4055 30607
rect 4069 30641 4121 30654
rect 4069 30607 4081 30641
rect 4081 30607 4115 30641
rect 4115 30607 4121 30641
rect 4069 30602 4121 30607
rect 4003 30568 4055 30588
rect 4003 30536 4009 30568
rect 4009 30536 4043 30568
rect 4043 30536 4055 30568
rect 4069 30568 4121 30588
rect 4069 30536 4081 30568
rect 4081 30536 4115 30568
rect 4115 30536 4121 30568
rect 4003 30495 4055 30522
rect 4003 30470 4009 30495
rect 4009 30470 4043 30495
rect 4043 30470 4055 30495
rect 4069 30495 4121 30522
rect 4069 30470 4081 30495
rect 4081 30470 4115 30495
rect 4115 30470 4121 30495
rect 4003 30422 4055 30456
rect 4069 30422 4121 30456
rect 4003 30404 4009 30422
rect 4009 30404 4055 30422
rect 4069 30404 4115 30422
rect 4115 30404 4121 30422
rect 4003 30338 4009 30390
rect 4009 30338 4055 30390
rect 4069 30338 4115 30390
rect 4115 30338 4121 30390
rect 4003 30271 4009 30323
rect 4009 30271 4055 30323
rect 4069 30271 4115 30323
rect 4115 30271 4121 30323
rect 4003 30204 4009 30256
rect 4009 30204 4055 30256
rect 4069 30204 4115 30256
rect 4115 30204 4121 30256
rect 4421 33840 4427 33892
rect 4427 33840 4473 33892
rect 4487 33840 4533 33892
rect 4533 33840 4539 33892
rect 4421 33774 4427 33826
rect 4427 33774 4473 33826
rect 4487 33774 4533 33826
rect 4533 33774 4539 33826
rect 4421 33708 4427 33760
rect 4427 33708 4473 33760
rect 4487 33708 4533 33760
rect 4533 33708 4539 33760
rect 4421 33642 4427 33694
rect 4427 33642 4473 33694
rect 4487 33642 4533 33694
rect 4533 33642 4539 33694
rect 4421 33575 4427 33627
rect 4427 33575 4473 33627
rect 4487 33575 4533 33627
rect 4533 33575 4539 33627
rect 4421 33508 4427 33560
rect 4427 33508 4473 33560
rect 4487 33508 4533 33560
rect 4533 33508 4539 33560
rect 4421 33441 4427 33493
rect 4427 33441 4473 33493
rect 4487 33441 4533 33493
rect 4533 33441 4539 33493
rect 4421 33380 4427 33426
rect 4427 33380 4473 33426
rect 4487 33380 4533 33426
rect 4533 33380 4539 33426
rect 4421 33374 4473 33380
rect 4487 33374 4539 33380
rect 4421 31840 4427 31892
rect 4427 31840 4473 31892
rect 4487 31840 4533 31892
rect 4533 31840 4539 31892
rect 4421 31774 4427 31826
rect 4427 31774 4473 31826
rect 4487 31774 4533 31826
rect 4533 31774 4539 31826
rect 4421 31708 4427 31760
rect 4427 31708 4473 31760
rect 4487 31708 4533 31760
rect 4533 31708 4539 31760
rect 4421 31642 4427 31694
rect 4427 31642 4473 31694
rect 4487 31642 4533 31694
rect 4533 31642 4539 31694
rect 4421 31575 4427 31627
rect 4427 31575 4473 31627
rect 4487 31575 4533 31627
rect 4533 31575 4539 31627
rect 4421 31508 4427 31560
rect 4427 31508 4473 31560
rect 4487 31508 4533 31560
rect 4533 31508 4539 31560
rect 4421 31441 4427 31493
rect 4427 31441 4473 31493
rect 4487 31441 4533 31493
rect 4533 31441 4539 31493
rect 4421 31380 4427 31426
rect 4427 31380 4473 31426
rect 4487 31380 4533 31426
rect 4533 31380 4539 31426
rect 4421 31374 4473 31380
rect 4487 31374 4539 31380
rect 4421 29840 4427 29892
rect 4427 29840 4473 29892
rect 4487 29840 4533 29892
rect 4533 29840 4539 29892
rect 4421 29774 4427 29826
rect 4427 29774 4473 29826
rect 4487 29774 4533 29826
rect 4533 29774 4539 29826
rect 4421 29708 4427 29760
rect 4427 29708 4473 29760
rect 4487 29708 4533 29760
rect 4533 29708 4539 29760
rect 4421 29642 4427 29694
rect 4427 29642 4473 29694
rect 4487 29642 4533 29694
rect 4533 29642 4539 29694
rect 4421 29575 4427 29627
rect 4427 29575 4473 29627
rect 4487 29575 4533 29627
rect 4533 29575 4539 29627
rect 4421 29508 4427 29560
rect 4427 29508 4473 29560
rect 4487 29508 4533 29560
rect 4533 29508 4539 29560
rect 4421 29441 4427 29493
rect 4427 29441 4473 29493
rect 4487 29441 4533 29493
rect 4533 29441 4539 29493
rect 4421 29380 4427 29426
rect 4427 29380 4473 29426
rect 4487 29380 4533 29426
rect 4533 29380 4539 29426
rect 4421 29374 4473 29380
rect 4487 29374 4539 29380
rect 4839 34714 4891 34720
rect 4839 34680 4845 34714
rect 4845 34680 4879 34714
rect 4879 34680 4891 34714
rect 4839 34668 4891 34680
rect 4905 34714 4957 34720
rect 4905 34680 4917 34714
rect 4917 34680 4951 34714
rect 4951 34680 4957 34714
rect 4905 34668 4957 34680
rect 4839 34641 4891 34654
rect 4839 34607 4845 34641
rect 4845 34607 4879 34641
rect 4879 34607 4891 34641
rect 4839 34602 4891 34607
rect 4905 34641 4957 34654
rect 4905 34607 4917 34641
rect 4917 34607 4951 34641
rect 4951 34607 4957 34641
rect 4905 34602 4957 34607
rect 4839 34568 4891 34588
rect 4839 34536 4845 34568
rect 4845 34536 4879 34568
rect 4879 34536 4891 34568
rect 4905 34568 4957 34588
rect 4905 34536 4917 34568
rect 4917 34536 4951 34568
rect 4951 34536 4957 34568
rect 4839 34495 4891 34522
rect 4839 34470 4845 34495
rect 4845 34470 4879 34495
rect 4879 34470 4891 34495
rect 4905 34495 4957 34522
rect 4905 34470 4917 34495
rect 4917 34470 4951 34495
rect 4951 34470 4957 34495
rect 4839 34422 4891 34456
rect 4905 34422 4957 34456
rect 4839 34404 4845 34422
rect 4845 34404 4891 34422
rect 4905 34404 4951 34422
rect 4951 34404 4957 34422
rect 4839 34338 4845 34390
rect 4845 34338 4891 34390
rect 4905 34338 4951 34390
rect 4951 34338 4957 34390
rect 4839 34271 4845 34323
rect 4845 34271 4891 34323
rect 4905 34271 4951 34323
rect 4951 34271 4957 34323
rect 4839 34204 4845 34256
rect 4845 34204 4891 34256
rect 4905 34204 4951 34256
rect 4951 34204 4957 34256
rect 4839 32714 4891 32720
rect 4839 32680 4845 32714
rect 4845 32680 4879 32714
rect 4879 32680 4891 32714
rect 4839 32668 4891 32680
rect 4905 32714 4957 32720
rect 4905 32680 4917 32714
rect 4917 32680 4951 32714
rect 4951 32680 4957 32714
rect 4905 32668 4957 32680
rect 4839 32641 4891 32654
rect 4839 32607 4845 32641
rect 4845 32607 4879 32641
rect 4879 32607 4891 32641
rect 4839 32602 4891 32607
rect 4905 32641 4957 32654
rect 4905 32607 4917 32641
rect 4917 32607 4951 32641
rect 4951 32607 4957 32641
rect 4905 32602 4957 32607
rect 4839 32568 4891 32588
rect 4839 32536 4845 32568
rect 4845 32536 4879 32568
rect 4879 32536 4891 32568
rect 4905 32568 4957 32588
rect 4905 32536 4917 32568
rect 4917 32536 4951 32568
rect 4951 32536 4957 32568
rect 4839 32495 4891 32522
rect 4839 32470 4845 32495
rect 4845 32470 4879 32495
rect 4879 32470 4891 32495
rect 4905 32495 4957 32522
rect 4905 32470 4917 32495
rect 4917 32470 4951 32495
rect 4951 32470 4957 32495
rect 4839 32422 4891 32456
rect 4905 32422 4957 32456
rect 4839 32404 4845 32422
rect 4845 32404 4891 32422
rect 4905 32404 4951 32422
rect 4951 32404 4957 32422
rect 4839 32338 4845 32390
rect 4845 32338 4891 32390
rect 4905 32338 4951 32390
rect 4951 32338 4957 32390
rect 4839 32271 4845 32323
rect 4845 32271 4891 32323
rect 4905 32271 4951 32323
rect 4951 32271 4957 32323
rect 4839 32204 4845 32256
rect 4845 32204 4891 32256
rect 4905 32204 4951 32256
rect 4951 32204 4957 32256
rect 4839 30714 4891 30720
rect 4839 30680 4845 30714
rect 4845 30680 4879 30714
rect 4879 30680 4891 30714
rect 4839 30668 4891 30680
rect 4905 30714 4957 30720
rect 4905 30680 4917 30714
rect 4917 30680 4951 30714
rect 4951 30680 4957 30714
rect 4905 30668 4957 30680
rect 4839 30641 4891 30654
rect 4839 30607 4845 30641
rect 4845 30607 4879 30641
rect 4879 30607 4891 30641
rect 4839 30602 4891 30607
rect 4905 30641 4957 30654
rect 4905 30607 4917 30641
rect 4917 30607 4951 30641
rect 4951 30607 4957 30641
rect 4905 30602 4957 30607
rect 4839 30568 4891 30588
rect 4839 30536 4845 30568
rect 4845 30536 4879 30568
rect 4879 30536 4891 30568
rect 4905 30568 4957 30588
rect 4905 30536 4917 30568
rect 4917 30536 4951 30568
rect 4951 30536 4957 30568
rect 4839 30495 4891 30522
rect 4839 30470 4845 30495
rect 4845 30470 4879 30495
rect 4879 30470 4891 30495
rect 4905 30495 4957 30522
rect 4905 30470 4917 30495
rect 4917 30470 4951 30495
rect 4951 30470 4957 30495
rect 4839 30422 4891 30456
rect 4905 30422 4957 30456
rect 4839 30404 4845 30422
rect 4845 30404 4891 30422
rect 4905 30404 4951 30422
rect 4951 30404 4957 30422
rect 4839 30338 4845 30390
rect 4845 30338 4891 30390
rect 4905 30338 4951 30390
rect 4951 30338 4957 30390
rect 4839 30271 4845 30323
rect 4845 30271 4891 30323
rect 4905 30271 4951 30323
rect 4951 30271 4957 30323
rect 4839 30204 4845 30256
rect 4845 30204 4891 30256
rect 4905 30204 4951 30256
rect 4951 30204 4957 30256
rect 3757 23645 3809 23697
rect 3831 23645 3883 23697
rect 3757 23573 3809 23625
rect 3831 23573 3883 23625
rect 3757 23501 3809 23553
rect 3831 23501 3883 23553
rect 3757 23428 3809 23480
rect 3831 23428 3883 23480
rect 3762 21723 3814 21775
rect 3826 21723 3878 21775
rect 4839 28714 4891 28720
rect 4839 28680 4845 28714
rect 4845 28680 4879 28714
rect 4879 28680 4891 28714
rect 4839 28668 4891 28680
rect 4905 28714 4957 28720
rect 4905 28680 4917 28714
rect 4917 28680 4951 28714
rect 4951 28680 4957 28714
rect 4905 28668 4957 28680
rect 4839 28641 4891 28654
rect 4839 28607 4845 28641
rect 4845 28607 4879 28641
rect 4879 28607 4891 28641
rect 4839 28602 4891 28607
rect 4905 28641 4957 28654
rect 4905 28607 4917 28641
rect 4917 28607 4951 28641
rect 4951 28607 4957 28641
rect 4905 28602 4957 28607
rect 4839 28568 4891 28588
rect 4839 28536 4845 28568
rect 4845 28536 4879 28568
rect 4879 28536 4891 28568
rect 4905 28568 4957 28588
rect 4905 28536 4917 28568
rect 4917 28536 4951 28568
rect 4951 28536 4957 28568
rect 4839 28495 4891 28522
rect 4839 28470 4845 28495
rect 4845 28470 4879 28495
rect 4879 28470 4891 28495
rect 4905 28495 4957 28522
rect 4905 28470 4917 28495
rect 4917 28470 4951 28495
rect 4951 28470 4957 28495
rect 4839 28422 4891 28456
rect 4905 28422 4957 28456
rect 4839 28404 4845 28422
rect 4845 28404 4891 28422
rect 4905 28404 4951 28422
rect 4951 28404 4957 28422
rect 4839 28338 4845 28390
rect 4845 28338 4891 28390
rect 4905 28338 4951 28390
rect 4951 28338 4957 28390
rect 4839 28271 4845 28323
rect 4845 28271 4891 28323
rect 4905 28271 4951 28323
rect 4951 28271 4957 28323
rect 4839 28204 4845 28256
rect 4845 28204 4891 28256
rect 4905 28204 4951 28256
rect 4951 28204 4957 28256
rect 4839 26718 4845 26720
rect 4845 26718 4879 26720
rect 4879 26718 4891 26720
rect 4839 26677 4891 26718
rect 4839 26668 4845 26677
rect 4845 26668 4879 26677
rect 4879 26668 4891 26677
rect 4905 26718 4917 26720
rect 4917 26718 4951 26720
rect 4951 26718 4957 26720
rect 4905 26677 4957 26718
rect 4905 26668 4917 26677
rect 4917 26668 4951 26677
rect 4951 26668 4957 26677
rect 4839 26643 4845 26654
rect 4845 26643 4879 26654
rect 4879 26643 4891 26654
rect 4839 26602 4891 26643
rect 4905 26643 4917 26654
rect 4917 26643 4951 26654
rect 4951 26643 4957 26654
rect 4905 26602 4957 26643
rect 4839 26568 4845 26588
rect 4845 26568 4879 26588
rect 4879 26568 4891 26588
rect 4839 26536 4891 26568
rect 4905 26568 4917 26588
rect 4917 26568 4951 26588
rect 4951 26568 4957 26588
rect 4905 26536 4957 26568
rect 4839 26493 4845 26522
rect 4845 26493 4879 26522
rect 4879 26493 4891 26522
rect 4839 26470 4891 26493
rect 4905 26493 4917 26522
rect 4917 26493 4951 26522
rect 4951 26493 4957 26522
rect 4905 26470 4957 26493
rect 4839 26452 4891 26456
rect 4839 26418 4845 26452
rect 4845 26418 4879 26452
rect 4879 26418 4891 26452
rect 4839 26404 4891 26418
rect 4905 26452 4957 26456
rect 4905 26418 4917 26452
rect 4917 26418 4951 26452
rect 4951 26418 4957 26452
rect 4905 26404 4957 26418
rect 4839 26377 4891 26389
rect 4839 26343 4845 26377
rect 4845 26343 4879 26377
rect 4879 26343 4891 26377
rect 4839 26337 4891 26343
rect 4905 26377 4957 26389
rect 4905 26343 4917 26377
rect 4917 26343 4951 26377
rect 4951 26343 4957 26377
rect 4905 26337 4957 26343
rect 4839 26302 4891 26322
rect 4839 26270 4845 26302
rect 4845 26270 4879 26302
rect 4879 26270 4891 26302
rect 4905 26302 4957 26322
rect 4905 26270 4917 26302
rect 4917 26270 4951 26302
rect 4951 26270 4957 26302
rect 4839 26227 4891 26255
rect 4839 26203 4845 26227
rect 4845 26203 4879 26227
rect 4879 26203 4891 26227
rect 4905 26227 4957 26255
rect 4905 26203 4917 26227
rect 4917 26203 4951 26227
rect 4951 26203 4957 26227
rect 5257 33840 5263 33892
rect 5263 33840 5309 33892
rect 5323 33840 5369 33892
rect 5369 33840 5375 33892
rect 5257 33774 5263 33826
rect 5263 33774 5309 33826
rect 5323 33774 5369 33826
rect 5369 33774 5375 33826
rect 5257 33708 5263 33760
rect 5263 33708 5309 33760
rect 5323 33708 5369 33760
rect 5369 33708 5375 33760
rect 5257 33642 5263 33694
rect 5263 33642 5309 33694
rect 5323 33642 5369 33694
rect 5369 33642 5375 33694
rect 5257 33575 5263 33627
rect 5263 33575 5309 33627
rect 5323 33575 5369 33627
rect 5369 33575 5375 33627
rect 5257 33508 5263 33560
rect 5263 33508 5309 33560
rect 5323 33508 5369 33560
rect 5369 33508 5375 33560
rect 5257 33441 5263 33493
rect 5263 33441 5309 33493
rect 5323 33441 5369 33493
rect 5369 33441 5375 33493
rect 5257 33380 5263 33426
rect 5263 33380 5309 33426
rect 5323 33380 5369 33426
rect 5369 33380 5375 33426
rect 5257 33374 5309 33380
rect 5323 33374 5375 33380
rect 5257 31840 5263 31892
rect 5263 31840 5309 31892
rect 5323 31840 5369 31892
rect 5369 31840 5375 31892
rect 5257 31774 5263 31826
rect 5263 31774 5309 31826
rect 5323 31774 5369 31826
rect 5369 31774 5375 31826
rect 5257 31708 5263 31760
rect 5263 31708 5309 31760
rect 5323 31708 5369 31760
rect 5369 31708 5375 31760
rect 5257 31642 5263 31694
rect 5263 31642 5309 31694
rect 5323 31642 5369 31694
rect 5369 31642 5375 31694
rect 5257 31575 5263 31627
rect 5263 31575 5309 31627
rect 5323 31575 5369 31627
rect 5369 31575 5375 31627
rect 5257 31508 5263 31560
rect 5263 31508 5309 31560
rect 5323 31508 5369 31560
rect 5369 31508 5375 31560
rect 5257 31441 5263 31493
rect 5263 31441 5309 31493
rect 5323 31441 5369 31493
rect 5369 31441 5375 31493
rect 5257 31380 5263 31426
rect 5263 31380 5309 31426
rect 5323 31380 5369 31426
rect 5369 31380 5375 31426
rect 5257 31374 5309 31380
rect 5323 31374 5375 31380
rect 5257 29840 5263 29892
rect 5263 29840 5309 29892
rect 5323 29840 5369 29892
rect 5369 29840 5375 29892
rect 5257 29774 5263 29826
rect 5263 29774 5309 29826
rect 5323 29774 5369 29826
rect 5369 29774 5375 29826
rect 5257 29708 5263 29760
rect 5263 29708 5309 29760
rect 5323 29708 5369 29760
rect 5369 29708 5375 29760
rect 5257 29642 5263 29694
rect 5263 29642 5309 29694
rect 5323 29642 5369 29694
rect 5369 29642 5375 29694
rect 5257 29575 5263 29627
rect 5263 29575 5309 29627
rect 5323 29575 5369 29627
rect 5369 29575 5375 29627
rect 5257 29508 5263 29560
rect 5263 29508 5309 29560
rect 5323 29508 5369 29560
rect 5369 29508 5375 29560
rect 5257 29441 5263 29493
rect 5263 29441 5309 29493
rect 5323 29441 5369 29493
rect 5369 29441 5375 29493
rect 5257 29380 5263 29426
rect 5263 29380 5309 29426
rect 5323 29380 5369 29426
rect 5369 29380 5375 29426
rect 5257 29374 5309 29380
rect 5323 29374 5375 29380
rect 5257 27840 5263 27892
rect 5263 27840 5309 27892
rect 5323 27840 5369 27892
rect 5369 27840 5375 27892
rect 5257 27774 5263 27826
rect 5263 27774 5309 27826
rect 5323 27774 5369 27826
rect 5369 27774 5375 27826
rect 5257 27708 5263 27760
rect 5263 27708 5309 27760
rect 5323 27708 5369 27760
rect 5369 27708 5375 27760
rect 5257 27642 5263 27694
rect 5263 27642 5309 27694
rect 5323 27642 5369 27694
rect 5369 27642 5375 27694
rect 5257 27575 5263 27627
rect 5263 27575 5309 27627
rect 5323 27575 5369 27627
rect 5369 27575 5375 27627
rect 5257 27508 5263 27560
rect 5263 27508 5309 27560
rect 5323 27508 5369 27560
rect 5369 27508 5375 27560
rect 5257 27441 5263 27493
rect 5263 27441 5309 27493
rect 5323 27441 5369 27493
rect 5369 27441 5375 27493
rect 5257 27380 5263 27426
rect 5263 27380 5309 27426
rect 5323 27380 5369 27426
rect 5369 27380 5375 27426
rect 5257 27374 5309 27380
rect 5323 27374 5375 27380
rect 5257 25854 5309 25891
rect 5257 25839 5263 25854
rect 5263 25839 5297 25854
rect 5297 25839 5309 25854
rect 5323 25854 5375 25891
rect 5323 25839 5335 25854
rect 5335 25839 5369 25854
rect 5369 25839 5375 25854
rect 5257 25820 5263 25825
rect 5263 25820 5297 25825
rect 5297 25820 5309 25825
rect 5257 25780 5309 25820
rect 5257 25773 5263 25780
rect 5263 25773 5297 25780
rect 5297 25773 5309 25780
rect 5323 25820 5335 25825
rect 5335 25820 5369 25825
rect 5369 25820 5375 25825
rect 5323 25780 5375 25820
rect 5323 25773 5335 25780
rect 5335 25773 5369 25780
rect 5369 25773 5375 25780
rect 5257 25746 5263 25759
rect 5263 25746 5297 25759
rect 5297 25746 5309 25759
rect 5257 25707 5309 25746
rect 5323 25746 5335 25759
rect 5335 25746 5369 25759
rect 5369 25746 5375 25759
rect 5323 25707 5375 25746
rect 5675 34714 5727 34720
rect 5675 34680 5681 34714
rect 5681 34680 5715 34714
rect 5715 34680 5727 34714
rect 5675 34668 5727 34680
rect 5741 34714 5793 34720
rect 5741 34680 5753 34714
rect 5753 34680 5787 34714
rect 5787 34680 5793 34714
rect 5741 34668 5793 34680
rect 5675 34641 5727 34654
rect 5675 34607 5681 34641
rect 5681 34607 5715 34641
rect 5715 34607 5727 34641
rect 5675 34602 5727 34607
rect 5741 34641 5793 34654
rect 5741 34607 5753 34641
rect 5753 34607 5787 34641
rect 5787 34607 5793 34641
rect 5741 34602 5793 34607
rect 5675 34568 5727 34588
rect 5675 34536 5681 34568
rect 5681 34536 5715 34568
rect 5715 34536 5727 34568
rect 5741 34568 5793 34588
rect 5741 34536 5753 34568
rect 5753 34536 5787 34568
rect 5787 34536 5793 34568
rect 5675 34495 5727 34522
rect 5675 34470 5681 34495
rect 5681 34470 5715 34495
rect 5715 34470 5727 34495
rect 5741 34495 5793 34522
rect 5741 34470 5753 34495
rect 5753 34470 5787 34495
rect 5787 34470 5793 34495
rect 5675 34422 5727 34456
rect 5741 34422 5793 34456
rect 5675 34404 5681 34422
rect 5681 34404 5727 34422
rect 5741 34404 5787 34422
rect 5787 34404 5793 34422
rect 5675 34338 5681 34390
rect 5681 34338 5727 34390
rect 5741 34338 5787 34390
rect 5787 34338 5793 34390
rect 5675 34271 5681 34323
rect 5681 34271 5727 34323
rect 5741 34271 5787 34323
rect 5787 34271 5793 34323
rect 5675 34204 5681 34256
rect 5681 34204 5727 34256
rect 5741 34204 5787 34256
rect 5787 34204 5793 34256
rect 5675 32714 5727 32720
rect 5675 32680 5681 32714
rect 5681 32680 5715 32714
rect 5715 32680 5727 32714
rect 5675 32668 5727 32680
rect 5741 32714 5793 32720
rect 5741 32680 5753 32714
rect 5753 32680 5787 32714
rect 5787 32680 5793 32714
rect 5741 32668 5793 32680
rect 5675 32641 5727 32654
rect 5675 32607 5681 32641
rect 5681 32607 5715 32641
rect 5715 32607 5727 32641
rect 5675 32602 5727 32607
rect 5741 32641 5793 32654
rect 5741 32607 5753 32641
rect 5753 32607 5787 32641
rect 5787 32607 5793 32641
rect 5741 32602 5793 32607
rect 5675 32568 5727 32588
rect 5675 32536 5681 32568
rect 5681 32536 5715 32568
rect 5715 32536 5727 32568
rect 5741 32568 5793 32588
rect 5741 32536 5753 32568
rect 5753 32536 5787 32568
rect 5787 32536 5793 32568
rect 5675 32495 5727 32522
rect 5675 32470 5681 32495
rect 5681 32470 5715 32495
rect 5715 32470 5727 32495
rect 5741 32495 5793 32522
rect 5741 32470 5753 32495
rect 5753 32470 5787 32495
rect 5787 32470 5793 32495
rect 5675 32422 5727 32456
rect 5741 32422 5793 32456
rect 5675 32404 5681 32422
rect 5681 32404 5727 32422
rect 5741 32404 5787 32422
rect 5787 32404 5793 32422
rect 5675 32338 5681 32390
rect 5681 32338 5727 32390
rect 5741 32338 5787 32390
rect 5787 32338 5793 32390
rect 5675 32271 5681 32323
rect 5681 32271 5727 32323
rect 5741 32271 5787 32323
rect 5787 32271 5793 32323
rect 5675 32204 5681 32256
rect 5681 32204 5727 32256
rect 5741 32204 5787 32256
rect 5787 32204 5793 32256
rect 5675 30714 5727 30720
rect 5675 30680 5681 30714
rect 5681 30680 5715 30714
rect 5715 30680 5727 30714
rect 5675 30668 5727 30680
rect 5741 30714 5793 30720
rect 5741 30680 5753 30714
rect 5753 30680 5787 30714
rect 5787 30680 5793 30714
rect 5741 30668 5793 30680
rect 5675 30641 5727 30654
rect 5675 30607 5681 30641
rect 5681 30607 5715 30641
rect 5715 30607 5727 30641
rect 5675 30602 5727 30607
rect 5741 30641 5793 30654
rect 5741 30607 5753 30641
rect 5753 30607 5787 30641
rect 5787 30607 5793 30641
rect 5741 30602 5793 30607
rect 5675 30568 5727 30588
rect 5675 30536 5681 30568
rect 5681 30536 5715 30568
rect 5715 30536 5727 30568
rect 5741 30568 5793 30588
rect 5741 30536 5753 30568
rect 5753 30536 5787 30568
rect 5787 30536 5793 30568
rect 5675 30495 5727 30522
rect 5675 30470 5681 30495
rect 5681 30470 5715 30495
rect 5715 30470 5727 30495
rect 5741 30495 5793 30522
rect 5741 30470 5753 30495
rect 5753 30470 5787 30495
rect 5787 30470 5793 30495
rect 5675 30422 5727 30456
rect 5741 30422 5793 30456
rect 5675 30404 5681 30422
rect 5681 30404 5727 30422
rect 5741 30404 5787 30422
rect 5787 30404 5793 30422
rect 5675 30338 5681 30390
rect 5681 30338 5727 30390
rect 5741 30338 5787 30390
rect 5787 30338 5793 30390
rect 5675 30271 5681 30323
rect 5681 30271 5727 30323
rect 5741 30271 5787 30323
rect 5787 30271 5793 30323
rect 5675 30204 5681 30256
rect 5681 30204 5727 30256
rect 5741 30204 5787 30256
rect 5787 30204 5793 30256
rect 5675 28714 5727 28720
rect 5675 28680 5681 28714
rect 5681 28680 5715 28714
rect 5715 28680 5727 28714
rect 5675 28668 5727 28680
rect 5741 28714 5793 28720
rect 5741 28680 5753 28714
rect 5753 28680 5787 28714
rect 5787 28680 5793 28714
rect 5741 28668 5793 28680
rect 5675 28641 5727 28654
rect 5675 28607 5681 28641
rect 5681 28607 5715 28641
rect 5715 28607 5727 28641
rect 5675 28602 5727 28607
rect 5741 28641 5793 28654
rect 5741 28607 5753 28641
rect 5753 28607 5787 28641
rect 5787 28607 5793 28641
rect 5741 28602 5793 28607
rect 5675 28568 5727 28588
rect 5675 28536 5681 28568
rect 5681 28536 5715 28568
rect 5715 28536 5727 28568
rect 5741 28568 5793 28588
rect 5741 28536 5753 28568
rect 5753 28536 5787 28568
rect 5787 28536 5793 28568
rect 5675 28495 5727 28522
rect 5675 28470 5681 28495
rect 5681 28470 5715 28495
rect 5715 28470 5727 28495
rect 5741 28495 5793 28522
rect 5741 28470 5753 28495
rect 5753 28470 5787 28495
rect 5787 28470 5793 28495
rect 5675 28422 5727 28456
rect 5741 28422 5793 28456
rect 5675 28404 5681 28422
rect 5681 28404 5727 28422
rect 5741 28404 5787 28422
rect 5787 28404 5793 28422
rect 5675 28338 5681 28390
rect 5681 28338 5727 28390
rect 5741 28338 5787 28390
rect 5787 28338 5793 28390
rect 5675 28271 5681 28323
rect 5681 28271 5727 28323
rect 5741 28271 5787 28323
rect 5787 28271 5793 28323
rect 5675 28204 5681 28256
rect 5681 28204 5727 28256
rect 5741 28204 5787 28256
rect 5787 28204 5793 28256
rect 5675 26718 5681 26720
rect 5681 26718 5715 26720
rect 5715 26718 5727 26720
rect 5675 26679 5727 26718
rect 5675 26668 5681 26679
rect 5681 26668 5715 26679
rect 5715 26668 5727 26679
rect 5741 26718 5753 26720
rect 5753 26718 5787 26720
rect 5787 26718 5793 26720
rect 5741 26679 5793 26718
rect 5741 26668 5753 26679
rect 5753 26668 5787 26679
rect 5787 26668 5793 26679
rect 5675 26645 5681 26654
rect 5681 26645 5715 26654
rect 5715 26645 5727 26654
rect 5675 26606 5727 26645
rect 5675 26602 5681 26606
rect 5681 26602 5715 26606
rect 5715 26602 5727 26606
rect 5741 26645 5753 26654
rect 5753 26645 5787 26654
rect 5787 26645 5793 26654
rect 5741 26606 5793 26645
rect 5741 26602 5753 26606
rect 5753 26602 5787 26606
rect 5787 26602 5793 26606
rect 5675 26572 5681 26588
rect 5681 26572 5715 26588
rect 5715 26572 5727 26588
rect 5675 26536 5727 26572
rect 5741 26572 5753 26588
rect 5753 26572 5787 26588
rect 5787 26572 5793 26588
rect 5741 26536 5793 26572
rect 5675 26499 5681 26522
rect 5681 26499 5715 26522
rect 5715 26499 5727 26522
rect 5675 26470 5727 26499
rect 5741 26499 5753 26522
rect 5753 26499 5787 26522
rect 5787 26499 5793 26522
rect 5741 26470 5793 26499
rect 5675 26426 5681 26456
rect 5681 26426 5715 26456
rect 5715 26426 5727 26456
rect 5675 26404 5727 26426
rect 5741 26426 5753 26456
rect 5753 26426 5787 26456
rect 5787 26426 5793 26456
rect 5741 26404 5793 26426
rect 5675 26387 5727 26389
rect 5675 26353 5681 26387
rect 5681 26353 5715 26387
rect 5715 26353 5727 26387
rect 5675 26337 5727 26353
rect 5741 26387 5793 26389
rect 5741 26353 5753 26387
rect 5753 26353 5787 26387
rect 5787 26353 5793 26387
rect 5741 26337 5793 26353
rect 5675 26314 5727 26322
rect 5675 26280 5681 26314
rect 5681 26280 5715 26314
rect 5715 26280 5727 26314
rect 5675 26270 5727 26280
rect 5741 26314 5793 26322
rect 5741 26280 5753 26314
rect 5753 26280 5787 26314
rect 5787 26280 5793 26314
rect 5741 26270 5793 26280
rect 5675 26241 5727 26255
rect 5675 26207 5681 26241
rect 5681 26207 5715 26241
rect 5715 26207 5727 26241
rect 5675 26203 5727 26207
rect 5741 26241 5793 26255
rect 5741 26207 5753 26241
rect 5753 26207 5787 26241
rect 5787 26207 5793 26241
rect 5741 26203 5793 26207
rect 6093 33840 6099 33892
rect 6099 33840 6145 33892
rect 6159 33840 6205 33892
rect 6205 33840 6211 33892
rect 6093 33774 6099 33826
rect 6099 33774 6145 33826
rect 6159 33774 6205 33826
rect 6205 33774 6211 33826
rect 6093 33708 6099 33760
rect 6099 33708 6145 33760
rect 6159 33708 6205 33760
rect 6205 33708 6211 33760
rect 6093 33642 6099 33694
rect 6099 33642 6145 33694
rect 6159 33642 6205 33694
rect 6205 33642 6211 33694
rect 6093 33575 6099 33627
rect 6099 33575 6145 33627
rect 6159 33575 6205 33627
rect 6205 33575 6211 33627
rect 6093 33508 6099 33560
rect 6099 33508 6145 33560
rect 6159 33508 6205 33560
rect 6205 33508 6211 33560
rect 6093 33441 6099 33493
rect 6099 33441 6145 33493
rect 6159 33441 6205 33493
rect 6205 33441 6211 33493
rect 6093 33380 6099 33426
rect 6099 33380 6145 33426
rect 6159 33380 6205 33426
rect 6205 33380 6211 33426
rect 6093 33374 6145 33380
rect 6159 33374 6211 33380
rect 6093 31840 6099 31892
rect 6099 31840 6145 31892
rect 6159 31840 6205 31892
rect 6205 31840 6211 31892
rect 6093 31774 6099 31826
rect 6099 31774 6145 31826
rect 6159 31774 6205 31826
rect 6205 31774 6211 31826
rect 6093 31708 6099 31760
rect 6099 31708 6145 31760
rect 6159 31708 6205 31760
rect 6205 31708 6211 31760
rect 6093 31642 6099 31694
rect 6099 31642 6145 31694
rect 6159 31642 6205 31694
rect 6205 31642 6211 31694
rect 6093 31575 6099 31627
rect 6099 31575 6145 31627
rect 6159 31575 6205 31627
rect 6205 31575 6211 31627
rect 6093 31508 6099 31560
rect 6099 31508 6145 31560
rect 6159 31508 6205 31560
rect 6205 31508 6211 31560
rect 6093 31441 6099 31493
rect 6099 31441 6145 31493
rect 6159 31441 6205 31493
rect 6205 31441 6211 31493
rect 6093 31380 6099 31426
rect 6099 31380 6145 31426
rect 6159 31380 6205 31426
rect 6205 31380 6211 31426
rect 6093 31374 6145 31380
rect 6159 31374 6211 31380
rect 6093 29840 6099 29892
rect 6099 29840 6145 29892
rect 6159 29840 6205 29892
rect 6205 29840 6211 29892
rect 6093 29774 6099 29826
rect 6099 29774 6145 29826
rect 6159 29774 6205 29826
rect 6205 29774 6211 29826
rect 6093 29708 6099 29760
rect 6099 29708 6145 29760
rect 6159 29708 6205 29760
rect 6205 29708 6211 29760
rect 6093 29642 6099 29694
rect 6099 29642 6145 29694
rect 6159 29642 6205 29694
rect 6205 29642 6211 29694
rect 6093 29575 6099 29627
rect 6099 29575 6145 29627
rect 6159 29575 6205 29627
rect 6205 29575 6211 29627
rect 6093 29508 6099 29560
rect 6099 29508 6145 29560
rect 6159 29508 6205 29560
rect 6205 29508 6211 29560
rect 6093 29441 6099 29493
rect 6099 29441 6145 29493
rect 6159 29441 6205 29493
rect 6205 29441 6211 29493
rect 6093 29380 6099 29426
rect 6099 29380 6145 29426
rect 6159 29380 6205 29426
rect 6205 29380 6211 29426
rect 6093 29374 6145 29380
rect 6159 29374 6211 29380
rect 6093 27840 6099 27892
rect 6099 27840 6145 27892
rect 6159 27840 6205 27892
rect 6205 27840 6211 27892
rect 6093 27774 6099 27826
rect 6099 27774 6145 27826
rect 6159 27774 6205 27826
rect 6205 27774 6211 27826
rect 6093 27708 6099 27760
rect 6099 27708 6145 27760
rect 6159 27708 6205 27760
rect 6205 27708 6211 27760
rect 6093 27642 6099 27694
rect 6099 27642 6145 27694
rect 6159 27642 6205 27694
rect 6205 27642 6211 27694
rect 6093 27575 6099 27627
rect 6099 27575 6145 27627
rect 6159 27575 6205 27627
rect 6205 27575 6211 27627
rect 6093 27508 6099 27560
rect 6099 27508 6145 27560
rect 6159 27508 6205 27560
rect 6205 27508 6211 27560
rect 6093 27441 6099 27493
rect 6099 27441 6145 27493
rect 6159 27441 6205 27493
rect 6205 27441 6211 27493
rect 6093 27380 6099 27426
rect 6099 27380 6145 27426
rect 6159 27380 6205 27426
rect 6205 27380 6211 27426
rect 6093 27374 6145 27380
rect 6159 27374 6211 27380
rect 6093 25854 6145 25891
rect 6093 25839 6099 25854
rect 6099 25839 6133 25854
rect 6133 25839 6145 25854
rect 6159 25854 6211 25891
rect 6159 25839 6171 25854
rect 6171 25839 6205 25854
rect 6205 25839 6211 25854
rect 6093 25820 6099 25825
rect 6099 25820 6133 25825
rect 6133 25820 6145 25825
rect 6093 25780 6145 25820
rect 6093 25773 6099 25780
rect 6099 25773 6133 25780
rect 6133 25773 6145 25780
rect 6159 25820 6171 25825
rect 6171 25820 6205 25825
rect 6205 25820 6211 25825
rect 6159 25780 6211 25820
rect 6159 25773 6171 25780
rect 6171 25773 6205 25780
rect 6205 25773 6211 25780
rect 6093 25746 6099 25759
rect 6099 25746 6133 25759
rect 6133 25746 6145 25759
rect 5257 25641 5309 25693
rect 5323 25641 5375 25693
rect 5257 25574 5309 25626
rect 5323 25574 5375 25626
rect 5257 25507 5309 25559
rect 5323 25507 5375 25559
rect 5257 25440 5309 25492
rect 5323 25440 5375 25492
rect 5257 25373 5309 25425
rect 5323 25373 5375 25425
rect 6093 25707 6145 25746
rect 6159 25746 6171 25759
rect 6171 25746 6205 25759
rect 6205 25746 6211 25759
rect 6159 25707 6211 25746
rect 6511 34714 6563 34720
rect 6511 34680 6517 34714
rect 6517 34680 6551 34714
rect 6551 34680 6563 34714
rect 6511 34668 6563 34680
rect 6577 34714 6629 34720
rect 6577 34680 6589 34714
rect 6589 34680 6623 34714
rect 6623 34680 6629 34714
rect 6577 34668 6629 34680
rect 6511 34641 6563 34654
rect 6511 34607 6517 34641
rect 6517 34607 6551 34641
rect 6551 34607 6563 34641
rect 6511 34602 6563 34607
rect 6577 34641 6629 34654
rect 6577 34607 6589 34641
rect 6589 34607 6623 34641
rect 6623 34607 6629 34641
rect 6577 34602 6629 34607
rect 6511 34568 6563 34588
rect 6511 34536 6517 34568
rect 6517 34536 6551 34568
rect 6551 34536 6563 34568
rect 6577 34568 6629 34588
rect 6577 34536 6589 34568
rect 6589 34536 6623 34568
rect 6623 34536 6629 34568
rect 6511 34495 6563 34522
rect 6511 34470 6517 34495
rect 6517 34470 6551 34495
rect 6551 34470 6563 34495
rect 6577 34495 6629 34522
rect 6577 34470 6589 34495
rect 6589 34470 6623 34495
rect 6623 34470 6629 34495
rect 6511 34422 6563 34456
rect 6577 34422 6629 34456
rect 6511 34404 6517 34422
rect 6517 34404 6563 34422
rect 6577 34404 6623 34422
rect 6623 34404 6629 34422
rect 6511 34338 6517 34390
rect 6517 34338 6563 34390
rect 6577 34338 6623 34390
rect 6623 34338 6629 34390
rect 6511 34271 6517 34323
rect 6517 34271 6563 34323
rect 6577 34271 6623 34323
rect 6623 34271 6629 34323
rect 6511 34204 6517 34256
rect 6517 34204 6563 34256
rect 6577 34204 6623 34256
rect 6623 34204 6629 34256
rect 6511 32714 6563 32720
rect 6511 32680 6517 32714
rect 6517 32680 6551 32714
rect 6551 32680 6563 32714
rect 6511 32668 6563 32680
rect 6577 32714 6629 32720
rect 6577 32680 6589 32714
rect 6589 32680 6623 32714
rect 6623 32680 6629 32714
rect 6577 32668 6629 32680
rect 6511 32641 6563 32654
rect 6511 32607 6517 32641
rect 6517 32607 6551 32641
rect 6551 32607 6563 32641
rect 6511 32602 6563 32607
rect 6577 32641 6629 32654
rect 6577 32607 6589 32641
rect 6589 32607 6623 32641
rect 6623 32607 6629 32641
rect 6577 32602 6629 32607
rect 6511 32568 6563 32588
rect 6511 32536 6517 32568
rect 6517 32536 6551 32568
rect 6551 32536 6563 32568
rect 6577 32568 6629 32588
rect 6577 32536 6589 32568
rect 6589 32536 6623 32568
rect 6623 32536 6629 32568
rect 6511 32495 6563 32522
rect 6511 32470 6517 32495
rect 6517 32470 6551 32495
rect 6551 32470 6563 32495
rect 6577 32495 6629 32522
rect 6577 32470 6589 32495
rect 6589 32470 6623 32495
rect 6623 32470 6629 32495
rect 6511 32422 6563 32456
rect 6577 32422 6629 32456
rect 6511 32404 6517 32422
rect 6517 32404 6563 32422
rect 6577 32404 6623 32422
rect 6623 32404 6629 32422
rect 6511 32338 6517 32390
rect 6517 32338 6563 32390
rect 6577 32338 6623 32390
rect 6623 32338 6629 32390
rect 6511 32271 6517 32323
rect 6517 32271 6563 32323
rect 6577 32271 6623 32323
rect 6623 32271 6629 32323
rect 6511 32204 6517 32256
rect 6517 32204 6563 32256
rect 6577 32204 6623 32256
rect 6623 32204 6629 32256
rect 6511 30714 6563 30720
rect 6511 30680 6517 30714
rect 6517 30680 6551 30714
rect 6551 30680 6563 30714
rect 6511 30668 6563 30680
rect 6577 30714 6629 30720
rect 6577 30680 6589 30714
rect 6589 30680 6623 30714
rect 6623 30680 6629 30714
rect 6577 30668 6629 30680
rect 6511 30641 6563 30654
rect 6511 30607 6517 30641
rect 6517 30607 6551 30641
rect 6551 30607 6563 30641
rect 6511 30602 6563 30607
rect 6577 30641 6629 30654
rect 6577 30607 6589 30641
rect 6589 30607 6623 30641
rect 6623 30607 6629 30641
rect 6577 30602 6629 30607
rect 6511 30568 6563 30588
rect 6511 30536 6517 30568
rect 6517 30536 6551 30568
rect 6551 30536 6563 30568
rect 6577 30568 6629 30588
rect 6577 30536 6589 30568
rect 6589 30536 6623 30568
rect 6623 30536 6629 30568
rect 6511 30495 6563 30522
rect 6511 30470 6517 30495
rect 6517 30470 6551 30495
rect 6551 30470 6563 30495
rect 6577 30495 6629 30522
rect 6577 30470 6589 30495
rect 6589 30470 6623 30495
rect 6623 30470 6629 30495
rect 6511 30422 6563 30456
rect 6577 30422 6629 30456
rect 6511 30404 6517 30422
rect 6517 30404 6563 30422
rect 6577 30404 6623 30422
rect 6623 30404 6629 30422
rect 6511 30338 6517 30390
rect 6517 30338 6563 30390
rect 6577 30338 6623 30390
rect 6623 30338 6629 30390
rect 6511 30271 6517 30323
rect 6517 30271 6563 30323
rect 6577 30271 6623 30323
rect 6623 30271 6629 30323
rect 6511 30204 6517 30256
rect 6517 30204 6563 30256
rect 6577 30204 6623 30256
rect 6623 30204 6629 30256
rect 6511 28714 6563 28720
rect 6511 28680 6517 28714
rect 6517 28680 6551 28714
rect 6551 28680 6563 28714
rect 6511 28668 6563 28680
rect 6577 28714 6629 28720
rect 6577 28680 6589 28714
rect 6589 28680 6623 28714
rect 6623 28680 6629 28714
rect 6577 28668 6629 28680
rect 6511 28641 6563 28654
rect 6511 28607 6517 28641
rect 6517 28607 6551 28641
rect 6551 28607 6563 28641
rect 6511 28602 6563 28607
rect 6577 28641 6629 28654
rect 6577 28607 6589 28641
rect 6589 28607 6623 28641
rect 6623 28607 6629 28641
rect 6577 28602 6629 28607
rect 6511 28568 6563 28588
rect 6511 28536 6517 28568
rect 6517 28536 6551 28568
rect 6551 28536 6563 28568
rect 6577 28568 6629 28588
rect 6577 28536 6589 28568
rect 6589 28536 6623 28568
rect 6623 28536 6629 28568
rect 6511 28495 6563 28522
rect 6511 28470 6517 28495
rect 6517 28470 6551 28495
rect 6551 28470 6563 28495
rect 6577 28495 6629 28522
rect 6577 28470 6589 28495
rect 6589 28470 6623 28495
rect 6623 28470 6629 28495
rect 6511 28422 6563 28456
rect 6577 28422 6629 28456
rect 6511 28404 6517 28422
rect 6517 28404 6563 28422
rect 6577 28404 6623 28422
rect 6623 28404 6629 28422
rect 6511 28338 6517 28390
rect 6517 28338 6563 28390
rect 6577 28338 6623 28390
rect 6623 28338 6629 28390
rect 6511 28271 6517 28323
rect 6517 28271 6563 28323
rect 6577 28271 6623 28323
rect 6623 28271 6629 28323
rect 6511 28204 6517 28256
rect 6517 28204 6563 28256
rect 6577 28204 6623 28256
rect 6623 28204 6629 28256
rect 6511 26717 6517 26720
rect 6517 26717 6551 26720
rect 6551 26717 6563 26720
rect 6511 26676 6563 26717
rect 6511 26668 6517 26676
rect 6517 26668 6551 26676
rect 6551 26668 6563 26676
rect 6577 26717 6589 26720
rect 6589 26717 6623 26720
rect 6623 26717 6629 26720
rect 6577 26676 6629 26717
rect 6577 26668 6589 26676
rect 6589 26668 6623 26676
rect 6623 26668 6629 26676
rect 6511 26642 6517 26654
rect 6517 26642 6551 26654
rect 6551 26642 6563 26654
rect 6511 26602 6563 26642
rect 6577 26642 6589 26654
rect 6589 26642 6623 26654
rect 6623 26642 6629 26654
rect 6577 26602 6629 26642
rect 6511 26567 6517 26588
rect 6517 26567 6551 26588
rect 6551 26567 6563 26588
rect 6511 26536 6563 26567
rect 6577 26567 6589 26588
rect 6589 26567 6623 26588
rect 6623 26567 6629 26588
rect 6577 26536 6629 26567
rect 6511 26492 6517 26522
rect 6517 26492 6551 26522
rect 6551 26492 6563 26522
rect 6511 26470 6563 26492
rect 6577 26492 6589 26522
rect 6589 26492 6623 26522
rect 6623 26492 6629 26522
rect 6577 26470 6629 26492
rect 6511 26451 6563 26456
rect 6511 26417 6517 26451
rect 6517 26417 6551 26451
rect 6551 26417 6563 26451
rect 6511 26404 6563 26417
rect 6577 26451 6629 26456
rect 6577 26417 6589 26451
rect 6589 26417 6623 26451
rect 6623 26417 6629 26451
rect 6577 26404 6629 26417
rect 6511 26376 6563 26389
rect 6511 26342 6517 26376
rect 6517 26342 6551 26376
rect 6551 26342 6563 26376
rect 6511 26337 6563 26342
rect 6577 26376 6629 26389
rect 6577 26342 6589 26376
rect 6589 26342 6623 26376
rect 6623 26342 6629 26376
rect 6577 26337 6629 26342
rect 6511 26301 6563 26322
rect 6511 26270 6517 26301
rect 6517 26270 6551 26301
rect 6551 26270 6563 26301
rect 6577 26301 6629 26322
rect 6577 26270 6589 26301
rect 6589 26270 6623 26301
rect 6623 26270 6629 26301
rect 6511 26226 6563 26255
rect 6511 26203 6517 26226
rect 6517 26203 6551 26226
rect 6551 26203 6563 26226
rect 6577 26226 6629 26255
rect 6577 26203 6589 26226
rect 6589 26203 6623 26226
rect 6623 26203 6629 26226
rect 6929 33840 6935 33892
rect 6935 33840 6981 33892
rect 6995 33840 7041 33892
rect 7041 33840 7047 33892
rect 6929 33774 6935 33826
rect 6935 33774 6981 33826
rect 6995 33774 7041 33826
rect 7041 33774 7047 33826
rect 6929 33708 6935 33760
rect 6935 33708 6981 33760
rect 6995 33708 7041 33760
rect 7041 33708 7047 33760
rect 6929 33642 6935 33694
rect 6935 33642 6981 33694
rect 6995 33642 7041 33694
rect 7041 33642 7047 33694
rect 6929 33575 6935 33627
rect 6935 33575 6981 33627
rect 6995 33575 7041 33627
rect 7041 33575 7047 33627
rect 6929 33508 6935 33560
rect 6935 33508 6981 33560
rect 6995 33508 7041 33560
rect 7041 33508 7047 33560
rect 6929 33441 6935 33493
rect 6935 33441 6981 33493
rect 6995 33441 7041 33493
rect 7041 33441 7047 33493
rect 6929 33380 6935 33426
rect 6935 33380 6981 33426
rect 6995 33380 7041 33426
rect 7041 33380 7047 33426
rect 6929 33374 6981 33380
rect 6995 33374 7047 33380
rect 6929 31840 6935 31892
rect 6935 31840 6981 31892
rect 6995 31840 7041 31892
rect 7041 31840 7047 31892
rect 6929 31774 6935 31826
rect 6935 31774 6981 31826
rect 6995 31774 7041 31826
rect 7041 31774 7047 31826
rect 6929 31708 6935 31760
rect 6935 31708 6981 31760
rect 6995 31708 7041 31760
rect 7041 31708 7047 31760
rect 6929 31642 6935 31694
rect 6935 31642 6981 31694
rect 6995 31642 7041 31694
rect 7041 31642 7047 31694
rect 6929 31575 6935 31627
rect 6935 31575 6981 31627
rect 6995 31575 7041 31627
rect 7041 31575 7047 31627
rect 6929 31508 6935 31560
rect 6935 31508 6981 31560
rect 6995 31508 7041 31560
rect 7041 31508 7047 31560
rect 6929 31441 6935 31493
rect 6935 31441 6981 31493
rect 6995 31441 7041 31493
rect 7041 31441 7047 31493
rect 6929 31380 6935 31426
rect 6935 31380 6981 31426
rect 6995 31380 7041 31426
rect 7041 31380 7047 31426
rect 6929 31374 6981 31380
rect 6995 31374 7047 31380
rect 6929 29840 6935 29892
rect 6935 29840 6981 29892
rect 6995 29840 7041 29892
rect 7041 29840 7047 29892
rect 6929 29774 6935 29826
rect 6935 29774 6981 29826
rect 6995 29774 7041 29826
rect 7041 29774 7047 29826
rect 6929 29708 6935 29760
rect 6935 29708 6981 29760
rect 6995 29708 7041 29760
rect 7041 29708 7047 29760
rect 6929 29642 6935 29694
rect 6935 29642 6981 29694
rect 6995 29642 7041 29694
rect 7041 29642 7047 29694
rect 6929 29575 6935 29627
rect 6935 29575 6981 29627
rect 6995 29575 7041 29627
rect 7041 29575 7047 29627
rect 6929 29508 6935 29560
rect 6935 29508 6981 29560
rect 6995 29508 7041 29560
rect 7041 29508 7047 29560
rect 6929 29441 6935 29493
rect 6935 29441 6981 29493
rect 6995 29441 7041 29493
rect 7041 29441 7047 29493
rect 6929 29380 6935 29426
rect 6935 29380 6981 29426
rect 6995 29380 7041 29426
rect 7041 29380 7047 29426
rect 6929 29374 6981 29380
rect 6995 29374 7047 29380
rect 6929 27840 6935 27892
rect 6935 27840 6981 27892
rect 6995 27840 7041 27892
rect 7041 27840 7047 27892
rect 6929 27774 6935 27826
rect 6935 27774 6981 27826
rect 6995 27774 7041 27826
rect 7041 27774 7047 27826
rect 6929 27708 6935 27760
rect 6935 27708 6981 27760
rect 6995 27708 7041 27760
rect 7041 27708 7047 27760
rect 6929 27642 6935 27694
rect 6935 27642 6981 27694
rect 6995 27642 7041 27694
rect 7041 27642 7047 27694
rect 6929 27575 6935 27627
rect 6935 27575 6981 27627
rect 6995 27575 7041 27627
rect 7041 27575 7047 27627
rect 6929 27508 6935 27560
rect 6935 27508 6981 27560
rect 6995 27508 7041 27560
rect 7041 27508 7047 27560
rect 6929 27441 6935 27493
rect 6935 27441 6981 27493
rect 6995 27441 7041 27493
rect 7041 27441 7047 27493
rect 6929 27380 6935 27426
rect 6935 27380 6981 27426
rect 6995 27380 7041 27426
rect 7041 27380 7047 27426
rect 6929 27374 6981 27380
rect 6995 27374 7047 27380
rect 6929 25856 6981 25891
rect 6929 25839 6935 25856
rect 6935 25839 6969 25856
rect 6969 25839 6981 25856
rect 6995 25856 7047 25891
rect 6995 25839 7007 25856
rect 7007 25839 7041 25856
rect 7041 25839 7047 25856
rect 6929 25822 6935 25825
rect 6935 25822 6969 25825
rect 6969 25822 6981 25825
rect 6929 25780 6981 25822
rect 6929 25773 6935 25780
rect 6935 25773 6969 25780
rect 6969 25773 6981 25780
rect 6995 25822 7007 25825
rect 7007 25822 7041 25825
rect 7041 25822 7047 25825
rect 6995 25780 7047 25822
rect 6995 25773 7007 25780
rect 7007 25773 7041 25780
rect 7041 25773 7047 25780
rect 6929 25746 6935 25759
rect 6935 25746 6969 25759
rect 6969 25746 6981 25759
rect 6093 25641 6145 25693
rect 6159 25641 6211 25693
rect 6093 25574 6145 25626
rect 6159 25574 6211 25626
rect 6093 25507 6145 25559
rect 6159 25507 6211 25559
rect 6093 25440 6145 25492
rect 6159 25440 6211 25492
rect 6093 25373 6145 25425
rect 6159 25373 6211 25425
rect 6929 25707 6981 25746
rect 6995 25746 7007 25759
rect 7007 25746 7041 25759
rect 7041 25746 7047 25759
rect 6995 25707 7047 25746
rect 7347 34714 7399 34720
rect 7347 34680 7353 34714
rect 7353 34680 7387 34714
rect 7387 34680 7399 34714
rect 7347 34668 7399 34680
rect 7413 34714 7465 34720
rect 7413 34680 7425 34714
rect 7425 34680 7459 34714
rect 7459 34680 7465 34714
rect 7413 34668 7465 34680
rect 7347 34641 7399 34654
rect 7347 34607 7353 34641
rect 7353 34607 7387 34641
rect 7387 34607 7399 34641
rect 7347 34602 7399 34607
rect 7413 34641 7465 34654
rect 7413 34607 7425 34641
rect 7425 34607 7459 34641
rect 7459 34607 7465 34641
rect 7413 34602 7465 34607
rect 7347 34568 7399 34588
rect 7347 34536 7353 34568
rect 7353 34536 7387 34568
rect 7387 34536 7399 34568
rect 7413 34568 7465 34588
rect 7413 34536 7425 34568
rect 7425 34536 7459 34568
rect 7459 34536 7465 34568
rect 7347 34495 7399 34522
rect 7347 34470 7353 34495
rect 7353 34470 7387 34495
rect 7387 34470 7399 34495
rect 7413 34495 7465 34522
rect 7413 34470 7425 34495
rect 7425 34470 7459 34495
rect 7459 34470 7465 34495
rect 7347 34422 7399 34456
rect 7413 34422 7465 34456
rect 7347 34404 7353 34422
rect 7353 34404 7399 34422
rect 7413 34404 7459 34422
rect 7459 34404 7465 34422
rect 7347 34338 7353 34390
rect 7353 34338 7399 34390
rect 7413 34338 7459 34390
rect 7459 34338 7465 34390
rect 7347 34271 7353 34323
rect 7353 34271 7399 34323
rect 7413 34271 7459 34323
rect 7459 34271 7465 34323
rect 7347 34204 7353 34256
rect 7353 34204 7399 34256
rect 7413 34204 7459 34256
rect 7459 34204 7465 34256
rect 7347 32714 7399 32720
rect 7347 32680 7353 32714
rect 7353 32680 7387 32714
rect 7387 32680 7399 32714
rect 7347 32668 7399 32680
rect 7413 32714 7465 32720
rect 7413 32680 7425 32714
rect 7425 32680 7459 32714
rect 7459 32680 7465 32714
rect 7413 32668 7465 32680
rect 7347 32641 7399 32654
rect 7347 32607 7353 32641
rect 7353 32607 7387 32641
rect 7387 32607 7399 32641
rect 7347 32602 7399 32607
rect 7413 32641 7465 32654
rect 7413 32607 7425 32641
rect 7425 32607 7459 32641
rect 7459 32607 7465 32641
rect 7413 32602 7465 32607
rect 7347 32568 7399 32588
rect 7347 32536 7353 32568
rect 7353 32536 7387 32568
rect 7387 32536 7399 32568
rect 7413 32568 7465 32588
rect 7413 32536 7425 32568
rect 7425 32536 7459 32568
rect 7459 32536 7465 32568
rect 7347 32495 7399 32522
rect 7347 32470 7353 32495
rect 7353 32470 7387 32495
rect 7387 32470 7399 32495
rect 7413 32495 7465 32522
rect 7413 32470 7425 32495
rect 7425 32470 7459 32495
rect 7459 32470 7465 32495
rect 7347 32422 7399 32456
rect 7413 32422 7465 32456
rect 7347 32404 7353 32422
rect 7353 32404 7399 32422
rect 7413 32404 7459 32422
rect 7459 32404 7465 32422
rect 7347 32338 7353 32390
rect 7353 32338 7399 32390
rect 7413 32338 7459 32390
rect 7459 32338 7465 32390
rect 7347 32271 7353 32323
rect 7353 32271 7399 32323
rect 7413 32271 7459 32323
rect 7459 32271 7465 32323
rect 7347 32204 7353 32256
rect 7353 32204 7399 32256
rect 7413 32204 7459 32256
rect 7459 32204 7465 32256
rect 7347 30714 7399 30720
rect 7347 30680 7353 30714
rect 7353 30680 7387 30714
rect 7387 30680 7399 30714
rect 7347 30668 7399 30680
rect 7413 30714 7465 30720
rect 7413 30680 7425 30714
rect 7425 30680 7459 30714
rect 7459 30680 7465 30714
rect 7413 30668 7465 30680
rect 7347 30641 7399 30654
rect 7347 30607 7353 30641
rect 7353 30607 7387 30641
rect 7387 30607 7399 30641
rect 7347 30602 7399 30607
rect 7413 30641 7465 30654
rect 7413 30607 7425 30641
rect 7425 30607 7459 30641
rect 7459 30607 7465 30641
rect 7413 30602 7465 30607
rect 7347 30568 7399 30588
rect 7347 30536 7353 30568
rect 7353 30536 7387 30568
rect 7387 30536 7399 30568
rect 7413 30568 7465 30588
rect 7413 30536 7425 30568
rect 7425 30536 7459 30568
rect 7459 30536 7465 30568
rect 7347 30495 7399 30522
rect 7347 30470 7353 30495
rect 7353 30470 7387 30495
rect 7387 30470 7399 30495
rect 7413 30495 7465 30522
rect 7413 30470 7425 30495
rect 7425 30470 7459 30495
rect 7459 30470 7465 30495
rect 7347 30422 7399 30456
rect 7413 30422 7465 30456
rect 7347 30404 7353 30422
rect 7353 30404 7399 30422
rect 7413 30404 7459 30422
rect 7459 30404 7465 30422
rect 7347 30338 7353 30390
rect 7353 30338 7399 30390
rect 7413 30338 7459 30390
rect 7459 30338 7465 30390
rect 7347 30271 7353 30323
rect 7353 30271 7399 30323
rect 7413 30271 7459 30323
rect 7459 30271 7465 30323
rect 7347 30204 7353 30256
rect 7353 30204 7399 30256
rect 7413 30204 7459 30256
rect 7459 30204 7465 30256
rect 7347 28714 7399 28720
rect 7347 28680 7353 28714
rect 7353 28680 7387 28714
rect 7387 28680 7399 28714
rect 7347 28668 7399 28680
rect 7413 28714 7465 28720
rect 7413 28680 7425 28714
rect 7425 28680 7459 28714
rect 7459 28680 7465 28714
rect 7413 28668 7465 28680
rect 7347 28641 7399 28654
rect 7347 28607 7353 28641
rect 7353 28607 7387 28641
rect 7387 28607 7399 28641
rect 7347 28602 7399 28607
rect 7413 28641 7465 28654
rect 7413 28607 7425 28641
rect 7425 28607 7459 28641
rect 7459 28607 7465 28641
rect 7413 28602 7465 28607
rect 7347 28568 7399 28588
rect 7347 28536 7353 28568
rect 7353 28536 7387 28568
rect 7387 28536 7399 28568
rect 7413 28568 7465 28588
rect 7413 28536 7425 28568
rect 7425 28536 7459 28568
rect 7459 28536 7465 28568
rect 7347 28495 7399 28522
rect 7347 28470 7353 28495
rect 7353 28470 7387 28495
rect 7387 28470 7399 28495
rect 7413 28495 7465 28522
rect 7413 28470 7425 28495
rect 7425 28470 7459 28495
rect 7459 28470 7465 28495
rect 7347 28422 7399 28456
rect 7413 28422 7465 28456
rect 7347 28404 7353 28422
rect 7353 28404 7399 28422
rect 7413 28404 7459 28422
rect 7459 28404 7465 28422
rect 7347 28338 7353 28390
rect 7353 28338 7399 28390
rect 7413 28338 7459 28390
rect 7459 28338 7465 28390
rect 7347 28271 7353 28323
rect 7353 28271 7399 28323
rect 7413 28271 7459 28323
rect 7459 28271 7465 28323
rect 7347 28204 7353 28256
rect 7353 28204 7399 28256
rect 7413 28204 7459 28256
rect 7459 28204 7465 28256
rect 7347 26717 7353 26720
rect 7353 26717 7387 26720
rect 7387 26717 7399 26720
rect 7347 26676 7399 26717
rect 7347 26668 7353 26676
rect 7353 26668 7387 26676
rect 7387 26668 7399 26676
rect 7413 26717 7425 26720
rect 7425 26717 7459 26720
rect 7459 26717 7465 26720
rect 7413 26676 7465 26717
rect 7413 26668 7425 26676
rect 7425 26668 7459 26676
rect 7459 26668 7465 26676
rect 7347 26642 7353 26654
rect 7353 26642 7387 26654
rect 7387 26642 7399 26654
rect 7347 26602 7399 26642
rect 7413 26642 7425 26654
rect 7425 26642 7459 26654
rect 7459 26642 7465 26654
rect 7413 26602 7465 26642
rect 7347 26567 7353 26588
rect 7353 26567 7387 26588
rect 7387 26567 7399 26588
rect 7347 26536 7399 26567
rect 7413 26567 7425 26588
rect 7425 26567 7459 26588
rect 7459 26567 7465 26588
rect 7413 26536 7465 26567
rect 7347 26492 7353 26522
rect 7353 26492 7387 26522
rect 7387 26492 7399 26522
rect 7347 26470 7399 26492
rect 7413 26492 7425 26522
rect 7425 26492 7459 26522
rect 7459 26492 7465 26522
rect 7413 26470 7465 26492
rect 7347 26451 7399 26456
rect 7347 26417 7353 26451
rect 7353 26417 7387 26451
rect 7387 26417 7399 26451
rect 7347 26404 7399 26417
rect 7413 26451 7465 26456
rect 7413 26417 7425 26451
rect 7425 26417 7459 26451
rect 7459 26417 7465 26451
rect 7413 26404 7465 26417
rect 7347 26376 7399 26389
rect 7347 26342 7353 26376
rect 7353 26342 7387 26376
rect 7387 26342 7399 26376
rect 7347 26337 7399 26342
rect 7413 26376 7465 26389
rect 7413 26342 7425 26376
rect 7425 26342 7459 26376
rect 7459 26342 7465 26376
rect 7413 26337 7465 26342
rect 7347 26301 7399 26322
rect 7347 26270 7353 26301
rect 7353 26270 7387 26301
rect 7387 26270 7399 26301
rect 7413 26301 7465 26322
rect 7413 26270 7425 26301
rect 7425 26270 7459 26301
rect 7459 26270 7465 26301
rect 7347 26226 7399 26255
rect 7347 26203 7353 26226
rect 7353 26203 7387 26226
rect 7387 26203 7399 26226
rect 7413 26226 7465 26255
rect 7413 26203 7425 26226
rect 7425 26203 7459 26226
rect 7459 26203 7465 26226
rect 7765 33840 7771 33892
rect 7771 33840 7817 33892
rect 7831 33840 7877 33892
rect 7877 33840 7883 33892
rect 7765 33774 7771 33826
rect 7771 33774 7817 33826
rect 7831 33774 7877 33826
rect 7877 33774 7883 33826
rect 7765 33708 7771 33760
rect 7771 33708 7817 33760
rect 7831 33708 7877 33760
rect 7877 33708 7883 33760
rect 7765 33642 7771 33694
rect 7771 33642 7817 33694
rect 7831 33642 7877 33694
rect 7877 33642 7883 33694
rect 7765 33575 7771 33627
rect 7771 33575 7817 33627
rect 7831 33575 7877 33627
rect 7877 33575 7883 33627
rect 7765 33508 7771 33560
rect 7771 33508 7817 33560
rect 7831 33508 7877 33560
rect 7877 33508 7883 33560
rect 7765 33441 7771 33493
rect 7771 33441 7817 33493
rect 7831 33441 7877 33493
rect 7877 33441 7883 33493
rect 7765 33380 7771 33426
rect 7771 33380 7817 33426
rect 7831 33380 7877 33426
rect 7877 33380 7883 33426
rect 7765 33374 7817 33380
rect 7831 33374 7883 33380
rect 7765 31840 7771 31892
rect 7771 31840 7817 31892
rect 7831 31840 7877 31892
rect 7877 31840 7883 31892
rect 7765 31774 7771 31826
rect 7771 31774 7817 31826
rect 7831 31774 7877 31826
rect 7877 31774 7883 31826
rect 7765 31708 7771 31760
rect 7771 31708 7817 31760
rect 7831 31708 7877 31760
rect 7877 31708 7883 31760
rect 7765 31642 7771 31694
rect 7771 31642 7817 31694
rect 7831 31642 7877 31694
rect 7877 31642 7883 31694
rect 7765 31575 7771 31627
rect 7771 31575 7817 31627
rect 7831 31575 7877 31627
rect 7877 31575 7883 31627
rect 7765 31508 7771 31560
rect 7771 31508 7817 31560
rect 7831 31508 7877 31560
rect 7877 31508 7883 31560
rect 7765 31441 7771 31493
rect 7771 31441 7817 31493
rect 7831 31441 7877 31493
rect 7877 31441 7883 31493
rect 7765 31380 7771 31426
rect 7771 31380 7817 31426
rect 7831 31380 7877 31426
rect 7877 31380 7883 31426
rect 7765 31374 7817 31380
rect 7831 31374 7883 31380
rect 7765 29840 7771 29892
rect 7771 29840 7817 29892
rect 7831 29840 7877 29892
rect 7877 29840 7883 29892
rect 7765 29774 7771 29826
rect 7771 29774 7817 29826
rect 7831 29774 7877 29826
rect 7877 29774 7883 29826
rect 7765 29708 7771 29760
rect 7771 29708 7817 29760
rect 7831 29708 7877 29760
rect 7877 29708 7883 29760
rect 7765 29642 7771 29694
rect 7771 29642 7817 29694
rect 7831 29642 7877 29694
rect 7877 29642 7883 29694
rect 7765 29575 7771 29627
rect 7771 29575 7817 29627
rect 7831 29575 7877 29627
rect 7877 29575 7883 29627
rect 7765 29508 7771 29560
rect 7771 29508 7817 29560
rect 7831 29508 7877 29560
rect 7877 29508 7883 29560
rect 7765 29441 7771 29493
rect 7771 29441 7817 29493
rect 7831 29441 7877 29493
rect 7877 29441 7883 29493
rect 7765 29380 7771 29426
rect 7771 29380 7817 29426
rect 7831 29380 7877 29426
rect 7877 29380 7883 29426
rect 7765 29374 7817 29380
rect 7831 29374 7883 29380
rect 7765 27840 7771 27892
rect 7771 27840 7817 27892
rect 7831 27840 7877 27892
rect 7877 27840 7883 27892
rect 7765 27774 7771 27826
rect 7771 27774 7817 27826
rect 7831 27774 7877 27826
rect 7877 27774 7883 27826
rect 7765 27708 7771 27760
rect 7771 27708 7817 27760
rect 7831 27708 7877 27760
rect 7877 27708 7883 27760
rect 7765 27642 7771 27694
rect 7771 27642 7817 27694
rect 7831 27642 7877 27694
rect 7877 27642 7883 27694
rect 7765 27575 7771 27627
rect 7771 27575 7817 27627
rect 7831 27575 7877 27627
rect 7877 27575 7883 27627
rect 7765 27508 7771 27560
rect 7771 27508 7817 27560
rect 7831 27508 7877 27560
rect 7877 27508 7883 27560
rect 7765 27441 7771 27493
rect 7771 27441 7817 27493
rect 7831 27441 7877 27493
rect 7877 27441 7883 27493
rect 7765 27380 7771 27426
rect 7771 27380 7817 27426
rect 7831 27380 7877 27426
rect 7877 27380 7883 27426
rect 7765 27374 7817 27380
rect 7831 27374 7883 27380
rect 7765 25857 7817 25891
rect 7765 25839 7771 25857
rect 7771 25839 7805 25857
rect 7805 25839 7817 25857
rect 7831 25857 7883 25891
rect 7831 25839 7843 25857
rect 7843 25839 7877 25857
rect 7877 25839 7883 25857
rect 7765 25823 7771 25825
rect 7771 25823 7805 25825
rect 7805 25823 7817 25825
rect 7765 25780 7817 25823
rect 7765 25773 7771 25780
rect 7771 25773 7805 25780
rect 7805 25773 7817 25780
rect 7831 25823 7843 25825
rect 7843 25823 7877 25825
rect 7877 25823 7883 25825
rect 7831 25780 7883 25823
rect 7831 25773 7843 25780
rect 7843 25773 7877 25780
rect 7877 25773 7883 25780
rect 7765 25746 7771 25759
rect 7771 25746 7805 25759
rect 7805 25746 7817 25759
rect 6929 25641 6981 25693
rect 6995 25641 7047 25693
rect 6929 25574 6981 25626
rect 6995 25574 7047 25626
rect 6929 25507 6981 25559
rect 6995 25507 7047 25559
rect 6929 25440 6981 25492
rect 6995 25440 7047 25492
rect 6929 25373 6981 25425
rect 6995 25373 7047 25425
rect 7765 25707 7817 25746
rect 7831 25746 7843 25759
rect 7843 25746 7877 25759
rect 7877 25746 7883 25759
rect 7831 25707 7883 25746
rect 8183 34714 8235 34720
rect 8183 34680 8189 34714
rect 8189 34680 8223 34714
rect 8223 34680 8235 34714
rect 8183 34668 8235 34680
rect 8249 34714 8301 34720
rect 8249 34680 8261 34714
rect 8261 34680 8295 34714
rect 8295 34680 8301 34714
rect 8249 34668 8301 34680
rect 8183 34641 8235 34654
rect 8183 34607 8189 34641
rect 8189 34607 8223 34641
rect 8223 34607 8235 34641
rect 8183 34602 8235 34607
rect 8249 34641 8301 34654
rect 8249 34607 8261 34641
rect 8261 34607 8295 34641
rect 8295 34607 8301 34641
rect 8249 34602 8301 34607
rect 8183 34568 8235 34588
rect 8183 34536 8189 34568
rect 8189 34536 8223 34568
rect 8223 34536 8235 34568
rect 8249 34568 8301 34588
rect 8249 34536 8261 34568
rect 8261 34536 8295 34568
rect 8295 34536 8301 34568
rect 8183 34495 8235 34522
rect 8183 34470 8189 34495
rect 8189 34470 8223 34495
rect 8223 34470 8235 34495
rect 8249 34495 8301 34522
rect 8249 34470 8261 34495
rect 8261 34470 8295 34495
rect 8295 34470 8301 34495
rect 8183 34422 8235 34456
rect 8249 34422 8301 34456
rect 8183 34404 8189 34422
rect 8189 34404 8235 34422
rect 8249 34404 8295 34422
rect 8295 34404 8301 34422
rect 8183 34338 8189 34390
rect 8189 34338 8235 34390
rect 8249 34338 8295 34390
rect 8295 34338 8301 34390
rect 8183 34271 8189 34323
rect 8189 34271 8235 34323
rect 8249 34271 8295 34323
rect 8295 34271 8301 34323
rect 8183 34204 8189 34256
rect 8189 34204 8235 34256
rect 8249 34204 8295 34256
rect 8295 34204 8301 34256
rect 8183 32714 8235 32720
rect 8183 32680 8189 32714
rect 8189 32680 8223 32714
rect 8223 32680 8235 32714
rect 8183 32668 8235 32680
rect 8249 32714 8301 32720
rect 8249 32680 8261 32714
rect 8261 32680 8295 32714
rect 8295 32680 8301 32714
rect 8249 32668 8301 32680
rect 8183 32641 8235 32654
rect 8183 32607 8189 32641
rect 8189 32607 8223 32641
rect 8223 32607 8235 32641
rect 8183 32602 8235 32607
rect 8249 32641 8301 32654
rect 8249 32607 8261 32641
rect 8261 32607 8295 32641
rect 8295 32607 8301 32641
rect 8249 32602 8301 32607
rect 8183 32568 8235 32588
rect 8183 32536 8189 32568
rect 8189 32536 8223 32568
rect 8223 32536 8235 32568
rect 8249 32568 8301 32588
rect 8249 32536 8261 32568
rect 8261 32536 8295 32568
rect 8295 32536 8301 32568
rect 8183 32495 8235 32522
rect 8183 32470 8189 32495
rect 8189 32470 8223 32495
rect 8223 32470 8235 32495
rect 8249 32495 8301 32522
rect 8249 32470 8261 32495
rect 8261 32470 8295 32495
rect 8295 32470 8301 32495
rect 8183 32422 8235 32456
rect 8249 32422 8301 32456
rect 8183 32404 8189 32422
rect 8189 32404 8235 32422
rect 8249 32404 8295 32422
rect 8295 32404 8301 32422
rect 8183 32338 8189 32390
rect 8189 32338 8235 32390
rect 8249 32338 8295 32390
rect 8295 32338 8301 32390
rect 8183 32271 8189 32323
rect 8189 32271 8235 32323
rect 8249 32271 8295 32323
rect 8295 32271 8301 32323
rect 8183 32204 8189 32256
rect 8189 32204 8235 32256
rect 8249 32204 8295 32256
rect 8295 32204 8301 32256
rect 8183 30714 8235 30720
rect 8183 30680 8189 30714
rect 8189 30680 8223 30714
rect 8223 30680 8235 30714
rect 8183 30668 8235 30680
rect 8249 30714 8301 30720
rect 8249 30680 8261 30714
rect 8261 30680 8295 30714
rect 8295 30680 8301 30714
rect 8249 30668 8301 30680
rect 8183 30641 8235 30654
rect 8183 30607 8189 30641
rect 8189 30607 8223 30641
rect 8223 30607 8235 30641
rect 8183 30602 8235 30607
rect 8249 30641 8301 30654
rect 8249 30607 8261 30641
rect 8261 30607 8295 30641
rect 8295 30607 8301 30641
rect 8249 30602 8301 30607
rect 8183 30568 8235 30588
rect 8183 30536 8189 30568
rect 8189 30536 8223 30568
rect 8223 30536 8235 30568
rect 8249 30568 8301 30588
rect 8249 30536 8261 30568
rect 8261 30536 8295 30568
rect 8295 30536 8301 30568
rect 8183 30495 8235 30522
rect 8183 30470 8189 30495
rect 8189 30470 8223 30495
rect 8223 30470 8235 30495
rect 8249 30495 8301 30522
rect 8249 30470 8261 30495
rect 8261 30470 8295 30495
rect 8295 30470 8301 30495
rect 8183 30422 8235 30456
rect 8249 30422 8301 30456
rect 8183 30404 8189 30422
rect 8189 30404 8235 30422
rect 8249 30404 8295 30422
rect 8295 30404 8301 30422
rect 8183 30338 8189 30390
rect 8189 30338 8235 30390
rect 8249 30338 8295 30390
rect 8295 30338 8301 30390
rect 8183 30271 8189 30323
rect 8189 30271 8235 30323
rect 8249 30271 8295 30323
rect 8295 30271 8301 30323
rect 8183 30204 8189 30256
rect 8189 30204 8235 30256
rect 8249 30204 8295 30256
rect 8295 30204 8301 30256
rect 8183 28714 8235 28720
rect 8183 28680 8189 28714
rect 8189 28680 8223 28714
rect 8223 28680 8235 28714
rect 8183 28668 8235 28680
rect 8249 28714 8301 28720
rect 8249 28680 8261 28714
rect 8261 28680 8295 28714
rect 8295 28680 8301 28714
rect 8249 28668 8301 28680
rect 8183 28641 8235 28654
rect 8183 28607 8189 28641
rect 8189 28607 8223 28641
rect 8223 28607 8235 28641
rect 8183 28602 8235 28607
rect 8249 28641 8301 28654
rect 8249 28607 8261 28641
rect 8261 28607 8295 28641
rect 8295 28607 8301 28641
rect 8249 28602 8301 28607
rect 8183 28568 8235 28588
rect 8183 28536 8189 28568
rect 8189 28536 8223 28568
rect 8223 28536 8235 28568
rect 8249 28568 8301 28588
rect 8249 28536 8261 28568
rect 8261 28536 8295 28568
rect 8295 28536 8301 28568
rect 8183 28495 8235 28522
rect 8183 28470 8189 28495
rect 8189 28470 8223 28495
rect 8223 28470 8235 28495
rect 8249 28495 8301 28522
rect 8249 28470 8261 28495
rect 8261 28470 8295 28495
rect 8295 28470 8301 28495
rect 8183 28422 8235 28456
rect 8249 28422 8301 28456
rect 8183 28404 8189 28422
rect 8189 28404 8235 28422
rect 8249 28404 8295 28422
rect 8295 28404 8301 28422
rect 8183 28338 8189 28390
rect 8189 28338 8235 28390
rect 8249 28338 8295 28390
rect 8295 28338 8301 28390
rect 8183 28271 8189 28323
rect 8189 28271 8235 28323
rect 8249 28271 8295 28323
rect 8295 28271 8301 28323
rect 8183 28204 8189 28256
rect 8189 28204 8235 28256
rect 8249 28204 8295 28256
rect 8295 28204 8301 28256
rect 8183 26717 8189 26720
rect 8189 26717 8223 26720
rect 8223 26717 8235 26720
rect 8183 26676 8235 26717
rect 8183 26668 8189 26676
rect 8189 26668 8223 26676
rect 8223 26668 8235 26676
rect 8249 26717 8261 26720
rect 8261 26717 8295 26720
rect 8295 26717 8301 26720
rect 8249 26676 8301 26717
rect 8249 26668 8261 26676
rect 8261 26668 8295 26676
rect 8295 26668 8301 26676
rect 8183 26642 8189 26654
rect 8189 26642 8223 26654
rect 8223 26642 8235 26654
rect 8183 26602 8235 26642
rect 8249 26642 8261 26654
rect 8261 26642 8295 26654
rect 8295 26642 8301 26654
rect 8249 26602 8301 26642
rect 8183 26567 8189 26588
rect 8189 26567 8223 26588
rect 8223 26567 8235 26588
rect 8183 26536 8235 26567
rect 8249 26567 8261 26588
rect 8261 26567 8295 26588
rect 8295 26567 8301 26588
rect 8249 26536 8301 26567
rect 8183 26492 8189 26522
rect 8189 26492 8223 26522
rect 8223 26492 8235 26522
rect 8183 26470 8235 26492
rect 8249 26492 8261 26522
rect 8261 26492 8295 26522
rect 8295 26492 8301 26522
rect 8249 26470 8301 26492
rect 8183 26451 8235 26456
rect 8183 26417 8189 26451
rect 8189 26417 8223 26451
rect 8223 26417 8235 26451
rect 8183 26404 8235 26417
rect 8249 26451 8301 26456
rect 8249 26417 8261 26451
rect 8261 26417 8295 26451
rect 8295 26417 8301 26451
rect 8249 26404 8301 26417
rect 8183 26376 8235 26389
rect 8183 26342 8189 26376
rect 8189 26342 8223 26376
rect 8223 26342 8235 26376
rect 8183 26337 8235 26342
rect 8249 26376 8301 26389
rect 8249 26342 8261 26376
rect 8261 26342 8295 26376
rect 8295 26342 8301 26376
rect 8249 26337 8301 26342
rect 8183 26301 8235 26322
rect 8183 26270 8189 26301
rect 8189 26270 8223 26301
rect 8223 26270 8235 26301
rect 8249 26301 8301 26322
rect 8249 26270 8261 26301
rect 8261 26270 8295 26301
rect 8295 26270 8301 26301
rect 8183 26226 8235 26255
rect 8183 26203 8189 26226
rect 8189 26203 8223 26226
rect 8223 26203 8235 26226
rect 8249 26226 8301 26255
rect 8249 26203 8261 26226
rect 8261 26203 8295 26226
rect 8295 26203 8301 26226
rect 8601 33840 8607 33892
rect 8607 33840 8653 33892
rect 8667 33840 8713 33892
rect 8713 33840 8719 33892
rect 8601 33774 8607 33826
rect 8607 33774 8653 33826
rect 8667 33774 8713 33826
rect 8713 33774 8719 33826
rect 8601 33708 8607 33760
rect 8607 33708 8653 33760
rect 8667 33708 8713 33760
rect 8713 33708 8719 33760
rect 8601 33642 8607 33694
rect 8607 33642 8653 33694
rect 8667 33642 8713 33694
rect 8713 33642 8719 33694
rect 8601 33575 8607 33627
rect 8607 33575 8653 33627
rect 8667 33575 8713 33627
rect 8713 33575 8719 33627
rect 8601 33508 8607 33560
rect 8607 33508 8653 33560
rect 8667 33508 8713 33560
rect 8713 33508 8719 33560
rect 8601 33441 8607 33493
rect 8607 33441 8653 33493
rect 8667 33441 8713 33493
rect 8713 33441 8719 33493
rect 8601 33380 8607 33426
rect 8607 33380 8653 33426
rect 8667 33380 8713 33426
rect 8713 33380 8719 33426
rect 8601 33374 8653 33380
rect 8667 33374 8719 33380
rect 8601 31840 8607 31892
rect 8607 31840 8653 31892
rect 8667 31840 8713 31892
rect 8713 31840 8719 31892
rect 8601 31774 8607 31826
rect 8607 31774 8653 31826
rect 8667 31774 8713 31826
rect 8713 31774 8719 31826
rect 8601 31708 8607 31760
rect 8607 31708 8653 31760
rect 8667 31708 8713 31760
rect 8713 31708 8719 31760
rect 8601 31642 8607 31694
rect 8607 31642 8653 31694
rect 8667 31642 8713 31694
rect 8713 31642 8719 31694
rect 8601 31575 8607 31627
rect 8607 31575 8653 31627
rect 8667 31575 8713 31627
rect 8713 31575 8719 31627
rect 8601 31508 8607 31560
rect 8607 31508 8653 31560
rect 8667 31508 8713 31560
rect 8713 31508 8719 31560
rect 8601 31441 8607 31493
rect 8607 31441 8653 31493
rect 8667 31441 8713 31493
rect 8713 31441 8719 31493
rect 8601 31380 8607 31426
rect 8607 31380 8653 31426
rect 8667 31380 8713 31426
rect 8713 31380 8719 31426
rect 8601 31374 8653 31380
rect 8667 31374 8719 31380
rect 8601 29840 8607 29892
rect 8607 29840 8653 29892
rect 8667 29840 8713 29892
rect 8713 29840 8719 29892
rect 8601 29774 8607 29826
rect 8607 29774 8653 29826
rect 8667 29774 8713 29826
rect 8713 29774 8719 29826
rect 8601 29708 8607 29760
rect 8607 29708 8653 29760
rect 8667 29708 8713 29760
rect 8713 29708 8719 29760
rect 8601 29642 8607 29694
rect 8607 29642 8653 29694
rect 8667 29642 8713 29694
rect 8713 29642 8719 29694
rect 8601 29575 8607 29627
rect 8607 29575 8653 29627
rect 8667 29575 8713 29627
rect 8713 29575 8719 29627
rect 8601 29508 8607 29560
rect 8607 29508 8653 29560
rect 8667 29508 8713 29560
rect 8713 29508 8719 29560
rect 8601 29441 8607 29493
rect 8607 29441 8653 29493
rect 8667 29441 8713 29493
rect 8713 29441 8719 29493
rect 8601 29380 8607 29426
rect 8607 29380 8653 29426
rect 8667 29380 8713 29426
rect 8713 29380 8719 29426
rect 8601 29374 8653 29380
rect 8667 29374 8719 29380
rect 8601 27840 8607 27892
rect 8607 27840 8653 27892
rect 8667 27840 8713 27892
rect 8713 27840 8719 27892
rect 8601 27774 8607 27826
rect 8607 27774 8653 27826
rect 8667 27774 8713 27826
rect 8713 27774 8719 27826
rect 8601 27708 8607 27760
rect 8607 27708 8653 27760
rect 8667 27708 8713 27760
rect 8713 27708 8719 27760
rect 8601 27642 8607 27694
rect 8607 27642 8653 27694
rect 8667 27642 8713 27694
rect 8713 27642 8719 27694
rect 8601 27575 8607 27627
rect 8607 27575 8653 27627
rect 8667 27575 8713 27627
rect 8713 27575 8719 27627
rect 8601 27508 8607 27560
rect 8607 27508 8653 27560
rect 8667 27508 8713 27560
rect 8713 27508 8719 27560
rect 8601 27441 8607 27493
rect 8607 27441 8653 27493
rect 8667 27441 8713 27493
rect 8713 27441 8719 27493
rect 8601 27380 8607 27426
rect 8607 27380 8653 27426
rect 8667 27380 8713 27426
rect 8713 27380 8719 27426
rect 8601 27374 8653 27380
rect 8667 27374 8719 27380
rect 8601 25857 8653 25891
rect 8601 25839 8607 25857
rect 8607 25839 8641 25857
rect 8641 25839 8653 25857
rect 8667 25857 8719 25891
rect 8667 25839 8679 25857
rect 8679 25839 8713 25857
rect 8713 25839 8719 25857
rect 8601 25823 8607 25825
rect 8607 25823 8641 25825
rect 8641 25823 8653 25825
rect 8601 25780 8653 25823
rect 8601 25773 8607 25780
rect 8607 25773 8641 25780
rect 8641 25773 8653 25780
rect 8667 25823 8679 25825
rect 8679 25823 8713 25825
rect 8713 25823 8719 25825
rect 8667 25780 8719 25823
rect 8667 25773 8679 25780
rect 8679 25773 8713 25780
rect 8713 25773 8719 25780
rect 8601 25746 8607 25759
rect 8607 25746 8641 25759
rect 8641 25746 8653 25759
rect 7765 25641 7817 25693
rect 7831 25641 7883 25693
rect 7765 25574 7817 25626
rect 7831 25574 7883 25626
rect 7765 25507 7817 25559
rect 7831 25507 7883 25559
rect 7765 25440 7817 25492
rect 7831 25440 7883 25492
rect 7765 25373 7817 25425
rect 7831 25373 7883 25425
rect 8601 25707 8653 25746
rect 8667 25746 8679 25759
rect 8679 25746 8713 25759
rect 8713 25746 8719 25759
rect 8667 25707 8719 25746
rect 9019 34714 9071 34720
rect 9019 34680 9025 34714
rect 9025 34680 9059 34714
rect 9059 34680 9071 34714
rect 9019 34668 9071 34680
rect 9085 34714 9137 34720
rect 9085 34680 9097 34714
rect 9097 34680 9131 34714
rect 9131 34680 9137 34714
rect 9085 34668 9137 34680
rect 9019 34641 9071 34654
rect 9019 34607 9025 34641
rect 9025 34607 9059 34641
rect 9059 34607 9071 34641
rect 9019 34602 9071 34607
rect 9085 34641 9137 34654
rect 9085 34607 9097 34641
rect 9097 34607 9131 34641
rect 9131 34607 9137 34641
rect 9085 34602 9137 34607
rect 9019 34568 9071 34588
rect 9019 34536 9025 34568
rect 9025 34536 9059 34568
rect 9059 34536 9071 34568
rect 9085 34568 9137 34588
rect 9085 34536 9097 34568
rect 9097 34536 9131 34568
rect 9131 34536 9137 34568
rect 9019 34495 9071 34522
rect 9019 34470 9025 34495
rect 9025 34470 9059 34495
rect 9059 34470 9071 34495
rect 9085 34495 9137 34522
rect 9085 34470 9097 34495
rect 9097 34470 9131 34495
rect 9131 34470 9137 34495
rect 9019 34422 9071 34456
rect 9085 34422 9137 34456
rect 9019 34404 9025 34422
rect 9025 34404 9071 34422
rect 9085 34404 9131 34422
rect 9131 34404 9137 34422
rect 9019 34338 9025 34390
rect 9025 34338 9071 34390
rect 9085 34338 9131 34390
rect 9131 34338 9137 34390
rect 9019 34271 9025 34323
rect 9025 34271 9071 34323
rect 9085 34271 9131 34323
rect 9131 34271 9137 34323
rect 9019 34204 9025 34256
rect 9025 34204 9071 34256
rect 9085 34204 9131 34256
rect 9131 34204 9137 34256
rect 9019 32714 9071 32720
rect 9019 32680 9025 32714
rect 9025 32680 9059 32714
rect 9059 32680 9071 32714
rect 9019 32668 9071 32680
rect 9085 32714 9137 32720
rect 9085 32680 9097 32714
rect 9097 32680 9131 32714
rect 9131 32680 9137 32714
rect 9085 32668 9137 32680
rect 9019 32641 9071 32654
rect 9019 32607 9025 32641
rect 9025 32607 9059 32641
rect 9059 32607 9071 32641
rect 9019 32602 9071 32607
rect 9085 32641 9137 32654
rect 9085 32607 9097 32641
rect 9097 32607 9131 32641
rect 9131 32607 9137 32641
rect 9085 32602 9137 32607
rect 9019 32568 9071 32588
rect 9019 32536 9025 32568
rect 9025 32536 9059 32568
rect 9059 32536 9071 32568
rect 9085 32568 9137 32588
rect 9085 32536 9097 32568
rect 9097 32536 9131 32568
rect 9131 32536 9137 32568
rect 9019 32495 9071 32522
rect 9019 32470 9025 32495
rect 9025 32470 9059 32495
rect 9059 32470 9071 32495
rect 9085 32495 9137 32522
rect 9085 32470 9097 32495
rect 9097 32470 9131 32495
rect 9131 32470 9137 32495
rect 9019 32422 9071 32456
rect 9085 32422 9137 32456
rect 9019 32404 9025 32422
rect 9025 32404 9071 32422
rect 9085 32404 9131 32422
rect 9131 32404 9137 32422
rect 9019 32338 9025 32390
rect 9025 32338 9071 32390
rect 9085 32338 9131 32390
rect 9131 32338 9137 32390
rect 9019 32271 9025 32323
rect 9025 32271 9071 32323
rect 9085 32271 9131 32323
rect 9131 32271 9137 32323
rect 9019 32204 9025 32256
rect 9025 32204 9071 32256
rect 9085 32204 9131 32256
rect 9131 32204 9137 32256
rect 9019 30714 9071 30720
rect 9019 30680 9025 30714
rect 9025 30680 9059 30714
rect 9059 30680 9071 30714
rect 9019 30668 9071 30680
rect 9085 30714 9137 30720
rect 9085 30680 9097 30714
rect 9097 30680 9131 30714
rect 9131 30680 9137 30714
rect 9085 30668 9137 30680
rect 9019 30641 9071 30654
rect 9019 30607 9025 30641
rect 9025 30607 9059 30641
rect 9059 30607 9071 30641
rect 9019 30602 9071 30607
rect 9085 30641 9137 30654
rect 9085 30607 9097 30641
rect 9097 30607 9131 30641
rect 9131 30607 9137 30641
rect 9085 30602 9137 30607
rect 9019 30568 9071 30588
rect 9019 30536 9025 30568
rect 9025 30536 9059 30568
rect 9059 30536 9071 30568
rect 9085 30568 9137 30588
rect 9085 30536 9097 30568
rect 9097 30536 9131 30568
rect 9131 30536 9137 30568
rect 9019 30495 9071 30522
rect 9019 30470 9025 30495
rect 9025 30470 9059 30495
rect 9059 30470 9071 30495
rect 9085 30495 9137 30522
rect 9085 30470 9097 30495
rect 9097 30470 9131 30495
rect 9131 30470 9137 30495
rect 9019 30422 9071 30456
rect 9085 30422 9137 30456
rect 9019 30404 9025 30422
rect 9025 30404 9071 30422
rect 9085 30404 9131 30422
rect 9131 30404 9137 30422
rect 9019 30338 9025 30390
rect 9025 30338 9071 30390
rect 9085 30338 9131 30390
rect 9131 30338 9137 30390
rect 9019 30271 9025 30323
rect 9025 30271 9071 30323
rect 9085 30271 9131 30323
rect 9131 30271 9137 30323
rect 9019 30204 9025 30256
rect 9025 30204 9071 30256
rect 9085 30204 9131 30256
rect 9131 30204 9137 30256
rect 9019 28714 9071 28720
rect 9019 28680 9025 28714
rect 9025 28680 9059 28714
rect 9059 28680 9071 28714
rect 9019 28668 9071 28680
rect 9085 28714 9137 28720
rect 9085 28680 9097 28714
rect 9097 28680 9131 28714
rect 9131 28680 9137 28714
rect 9085 28668 9137 28680
rect 9019 28641 9071 28654
rect 9019 28607 9025 28641
rect 9025 28607 9059 28641
rect 9059 28607 9071 28641
rect 9019 28602 9071 28607
rect 9085 28641 9137 28654
rect 9085 28607 9097 28641
rect 9097 28607 9131 28641
rect 9131 28607 9137 28641
rect 9085 28602 9137 28607
rect 9019 28568 9071 28588
rect 9019 28536 9025 28568
rect 9025 28536 9059 28568
rect 9059 28536 9071 28568
rect 9085 28568 9137 28588
rect 9085 28536 9097 28568
rect 9097 28536 9131 28568
rect 9131 28536 9137 28568
rect 9019 28495 9071 28522
rect 9019 28470 9025 28495
rect 9025 28470 9059 28495
rect 9059 28470 9071 28495
rect 9085 28495 9137 28522
rect 9085 28470 9097 28495
rect 9097 28470 9131 28495
rect 9131 28470 9137 28495
rect 9019 28422 9071 28456
rect 9085 28422 9137 28456
rect 9019 28404 9025 28422
rect 9025 28404 9071 28422
rect 9085 28404 9131 28422
rect 9131 28404 9137 28422
rect 9019 28338 9025 28390
rect 9025 28338 9071 28390
rect 9085 28338 9131 28390
rect 9131 28338 9137 28390
rect 9019 28271 9025 28323
rect 9025 28271 9071 28323
rect 9085 28271 9131 28323
rect 9131 28271 9137 28323
rect 9019 28204 9025 28256
rect 9025 28204 9071 28256
rect 9085 28204 9131 28256
rect 9131 28204 9137 28256
rect 9019 26717 9025 26720
rect 9025 26717 9059 26720
rect 9059 26717 9071 26720
rect 9019 26676 9071 26717
rect 9019 26668 9025 26676
rect 9025 26668 9059 26676
rect 9059 26668 9071 26676
rect 9085 26717 9097 26720
rect 9097 26717 9131 26720
rect 9131 26717 9137 26720
rect 9085 26676 9137 26717
rect 9085 26668 9097 26676
rect 9097 26668 9131 26676
rect 9131 26668 9137 26676
rect 9019 26642 9025 26654
rect 9025 26642 9059 26654
rect 9059 26642 9071 26654
rect 9019 26602 9071 26642
rect 9085 26642 9097 26654
rect 9097 26642 9131 26654
rect 9131 26642 9137 26654
rect 9085 26602 9137 26642
rect 9019 26567 9025 26588
rect 9025 26567 9059 26588
rect 9059 26567 9071 26588
rect 9019 26536 9071 26567
rect 9085 26567 9097 26588
rect 9097 26567 9131 26588
rect 9131 26567 9137 26588
rect 9085 26536 9137 26567
rect 9019 26492 9025 26522
rect 9025 26492 9059 26522
rect 9059 26492 9071 26522
rect 9019 26470 9071 26492
rect 9085 26492 9097 26522
rect 9097 26492 9131 26522
rect 9131 26492 9137 26522
rect 9085 26470 9137 26492
rect 9019 26451 9071 26456
rect 9019 26417 9025 26451
rect 9025 26417 9059 26451
rect 9059 26417 9071 26451
rect 9019 26404 9071 26417
rect 9085 26451 9137 26456
rect 9085 26417 9097 26451
rect 9097 26417 9131 26451
rect 9131 26417 9137 26451
rect 9085 26404 9137 26417
rect 9019 26376 9071 26389
rect 9019 26342 9025 26376
rect 9025 26342 9059 26376
rect 9059 26342 9071 26376
rect 9019 26337 9071 26342
rect 9085 26376 9137 26389
rect 9085 26342 9097 26376
rect 9097 26342 9131 26376
rect 9131 26342 9137 26376
rect 9085 26337 9137 26342
rect 9019 26301 9071 26322
rect 9019 26270 9025 26301
rect 9025 26270 9059 26301
rect 9059 26270 9071 26301
rect 9085 26301 9137 26322
rect 9085 26270 9097 26301
rect 9097 26270 9131 26301
rect 9131 26270 9137 26301
rect 9019 26226 9071 26255
rect 9019 26203 9025 26226
rect 9025 26203 9059 26226
rect 9059 26203 9071 26226
rect 9085 26226 9137 26255
rect 9085 26203 9097 26226
rect 9097 26203 9131 26226
rect 9131 26203 9137 26226
rect 9437 33840 9443 33892
rect 9443 33840 9489 33892
rect 9503 33840 9549 33892
rect 9549 33840 9555 33892
rect 9437 33774 9443 33826
rect 9443 33774 9489 33826
rect 9503 33774 9549 33826
rect 9549 33774 9555 33826
rect 9437 33708 9443 33760
rect 9443 33708 9489 33760
rect 9503 33708 9549 33760
rect 9549 33708 9555 33760
rect 9437 33642 9443 33694
rect 9443 33642 9489 33694
rect 9503 33642 9549 33694
rect 9549 33642 9555 33694
rect 9437 33575 9443 33627
rect 9443 33575 9489 33627
rect 9503 33575 9549 33627
rect 9549 33575 9555 33627
rect 9437 33508 9443 33560
rect 9443 33508 9489 33560
rect 9503 33508 9549 33560
rect 9549 33508 9555 33560
rect 9437 33441 9443 33493
rect 9443 33441 9489 33493
rect 9503 33441 9549 33493
rect 9549 33441 9555 33493
rect 9437 33380 9443 33426
rect 9443 33380 9489 33426
rect 9503 33380 9549 33426
rect 9549 33380 9555 33426
rect 9437 33374 9489 33380
rect 9503 33374 9555 33380
rect 9437 31840 9443 31892
rect 9443 31840 9489 31892
rect 9503 31840 9549 31892
rect 9549 31840 9555 31892
rect 9437 31774 9443 31826
rect 9443 31774 9489 31826
rect 9503 31774 9549 31826
rect 9549 31774 9555 31826
rect 9437 31708 9443 31760
rect 9443 31708 9489 31760
rect 9503 31708 9549 31760
rect 9549 31708 9555 31760
rect 9437 31642 9443 31694
rect 9443 31642 9489 31694
rect 9503 31642 9549 31694
rect 9549 31642 9555 31694
rect 9437 31575 9443 31627
rect 9443 31575 9489 31627
rect 9503 31575 9549 31627
rect 9549 31575 9555 31627
rect 9437 31508 9443 31560
rect 9443 31508 9489 31560
rect 9503 31508 9549 31560
rect 9549 31508 9555 31560
rect 9437 31441 9443 31493
rect 9443 31441 9489 31493
rect 9503 31441 9549 31493
rect 9549 31441 9555 31493
rect 9437 31380 9443 31426
rect 9443 31380 9489 31426
rect 9503 31380 9549 31426
rect 9549 31380 9555 31426
rect 9437 31374 9489 31380
rect 9503 31374 9555 31380
rect 9437 29840 9443 29892
rect 9443 29840 9489 29892
rect 9503 29840 9549 29892
rect 9549 29840 9555 29892
rect 9437 29774 9443 29826
rect 9443 29774 9489 29826
rect 9503 29774 9549 29826
rect 9549 29774 9555 29826
rect 9437 29708 9443 29760
rect 9443 29708 9489 29760
rect 9503 29708 9549 29760
rect 9549 29708 9555 29760
rect 9437 29642 9443 29694
rect 9443 29642 9489 29694
rect 9503 29642 9549 29694
rect 9549 29642 9555 29694
rect 9437 29575 9443 29627
rect 9443 29575 9489 29627
rect 9503 29575 9549 29627
rect 9549 29575 9555 29627
rect 9437 29508 9443 29560
rect 9443 29508 9489 29560
rect 9503 29508 9549 29560
rect 9549 29508 9555 29560
rect 9437 29441 9443 29493
rect 9443 29441 9489 29493
rect 9503 29441 9549 29493
rect 9549 29441 9555 29493
rect 9437 29380 9443 29426
rect 9443 29380 9489 29426
rect 9503 29380 9549 29426
rect 9549 29380 9555 29426
rect 9437 29374 9489 29380
rect 9503 29374 9555 29380
rect 9437 27840 9443 27892
rect 9443 27840 9489 27892
rect 9503 27840 9549 27892
rect 9549 27840 9555 27892
rect 9437 27774 9443 27826
rect 9443 27774 9489 27826
rect 9503 27774 9549 27826
rect 9549 27774 9555 27826
rect 9437 27708 9443 27760
rect 9443 27708 9489 27760
rect 9503 27708 9549 27760
rect 9549 27708 9555 27760
rect 9437 27642 9443 27694
rect 9443 27642 9489 27694
rect 9503 27642 9549 27694
rect 9549 27642 9555 27694
rect 9437 27575 9443 27627
rect 9443 27575 9489 27627
rect 9503 27575 9549 27627
rect 9549 27575 9555 27627
rect 9437 27508 9443 27560
rect 9443 27508 9489 27560
rect 9503 27508 9549 27560
rect 9549 27508 9555 27560
rect 9437 27441 9443 27493
rect 9443 27441 9489 27493
rect 9503 27441 9549 27493
rect 9549 27441 9555 27493
rect 9437 27380 9443 27426
rect 9443 27380 9489 27426
rect 9503 27380 9549 27426
rect 9549 27380 9555 27426
rect 9437 27374 9489 27380
rect 9503 27374 9555 27380
rect 9437 25857 9489 25891
rect 9437 25839 9443 25857
rect 9443 25839 9477 25857
rect 9477 25839 9489 25857
rect 9503 25857 9555 25891
rect 9503 25839 9515 25857
rect 9515 25839 9549 25857
rect 9549 25839 9555 25857
rect 9437 25823 9443 25825
rect 9443 25823 9477 25825
rect 9477 25823 9489 25825
rect 9437 25780 9489 25823
rect 9437 25773 9443 25780
rect 9443 25773 9477 25780
rect 9477 25773 9489 25780
rect 9503 25823 9515 25825
rect 9515 25823 9549 25825
rect 9549 25823 9555 25825
rect 9503 25780 9555 25823
rect 9503 25773 9515 25780
rect 9515 25773 9549 25780
rect 9549 25773 9555 25780
rect 9437 25746 9443 25759
rect 9443 25746 9477 25759
rect 9477 25746 9489 25759
rect 8601 25641 8653 25693
rect 8667 25641 8719 25693
rect 8601 25574 8653 25626
rect 8667 25574 8719 25626
rect 8601 25507 8653 25559
rect 8667 25507 8719 25559
rect 8601 25440 8653 25492
rect 8667 25440 8719 25492
rect 8601 25373 8653 25425
rect 8667 25373 8719 25425
rect 9437 25707 9489 25746
rect 9503 25746 9515 25759
rect 9515 25746 9549 25759
rect 9549 25746 9555 25759
rect 9503 25707 9555 25746
rect 9855 34714 9907 34720
rect 9855 34680 9861 34714
rect 9861 34680 9895 34714
rect 9895 34680 9907 34714
rect 9855 34668 9907 34680
rect 9921 34714 9973 34720
rect 9921 34680 9933 34714
rect 9933 34680 9967 34714
rect 9967 34680 9973 34714
rect 9921 34668 9973 34680
rect 9855 34641 9907 34654
rect 9855 34607 9861 34641
rect 9861 34607 9895 34641
rect 9895 34607 9907 34641
rect 9855 34602 9907 34607
rect 9921 34641 9973 34654
rect 9921 34607 9933 34641
rect 9933 34607 9967 34641
rect 9967 34607 9973 34641
rect 9921 34602 9973 34607
rect 9855 34568 9907 34588
rect 9855 34536 9861 34568
rect 9861 34536 9895 34568
rect 9895 34536 9907 34568
rect 9921 34568 9973 34588
rect 9921 34536 9933 34568
rect 9933 34536 9967 34568
rect 9967 34536 9973 34568
rect 9855 34495 9907 34522
rect 9855 34470 9861 34495
rect 9861 34470 9895 34495
rect 9895 34470 9907 34495
rect 9921 34495 9973 34522
rect 9921 34470 9933 34495
rect 9933 34470 9967 34495
rect 9967 34470 9973 34495
rect 9855 34422 9907 34456
rect 9921 34422 9973 34456
rect 9855 34404 9861 34422
rect 9861 34404 9907 34422
rect 9921 34404 9967 34422
rect 9967 34404 9973 34422
rect 9855 34338 9861 34390
rect 9861 34338 9907 34390
rect 9921 34338 9967 34390
rect 9967 34338 9973 34390
rect 9855 34271 9861 34323
rect 9861 34271 9907 34323
rect 9921 34271 9967 34323
rect 9967 34271 9973 34323
rect 9855 34204 9861 34256
rect 9861 34204 9907 34256
rect 9921 34204 9967 34256
rect 9967 34204 9973 34256
rect 9855 32714 9907 32720
rect 9855 32680 9861 32714
rect 9861 32680 9895 32714
rect 9895 32680 9907 32714
rect 9855 32668 9907 32680
rect 9921 32714 9973 32720
rect 9921 32680 9933 32714
rect 9933 32680 9967 32714
rect 9967 32680 9973 32714
rect 9921 32668 9973 32680
rect 9855 32641 9907 32654
rect 9855 32607 9861 32641
rect 9861 32607 9895 32641
rect 9895 32607 9907 32641
rect 9855 32602 9907 32607
rect 9921 32641 9973 32654
rect 9921 32607 9933 32641
rect 9933 32607 9967 32641
rect 9967 32607 9973 32641
rect 9921 32602 9973 32607
rect 9855 32568 9907 32588
rect 9855 32536 9861 32568
rect 9861 32536 9895 32568
rect 9895 32536 9907 32568
rect 9921 32568 9973 32588
rect 9921 32536 9933 32568
rect 9933 32536 9967 32568
rect 9967 32536 9973 32568
rect 9855 32495 9907 32522
rect 9855 32470 9861 32495
rect 9861 32470 9895 32495
rect 9895 32470 9907 32495
rect 9921 32495 9973 32522
rect 9921 32470 9933 32495
rect 9933 32470 9967 32495
rect 9967 32470 9973 32495
rect 9855 32422 9907 32456
rect 9921 32422 9973 32456
rect 9855 32404 9861 32422
rect 9861 32404 9907 32422
rect 9921 32404 9967 32422
rect 9967 32404 9973 32422
rect 9855 32338 9861 32390
rect 9861 32338 9907 32390
rect 9921 32338 9967 32390
rect 9967 32338 9973 32390
rect 9855 32271 9861 32323
rect 9861 32271 9907 32323
rect 9921 32271 9967 32323
rect 9967 32271 9973 32323
rect 9855 32204 9861 32256
rect 9861 32204 9907 32256
rect 9921 32204 9967 32256
rect 9967 32204 9973 32256
rect 9855 30714 9907 30720
rect 9855 30680 9861 30714
rect 9861 30680 9895 30714
rect 9895 30680 9907 30714
rect 9855 30668 9907 30680
rect 9921 30714 9973 30720
rect 9921 30680 9933 30714
rect 9933 30680 9967 30714
rect 9967 30680 9973 30714
rect 9921 30668 9973 30680
rect 9855 30641 9907 30654
rect 9855 30607 9861 30641
rect 9861 30607 9895 30641
rect 9895 30607 9907 30641
rect 9855 30602 9907 30607
rect 9921 30641 9973 30654
rect 9921 30607 9933 30641
rect 9933 30607 9967 30641
rect 9967 30607 9973 30641
rect 9921 30602 9973 30607
rect 9855 30568 9907 30588
rect 9855 30536 9861 30568
rect 9861 30536 9895 30568
rect 9895 30536 9907 30568
rect 9921 30568 9973 30588
rect 9921 30536 9933 30568
rect 9933 30536 9967 30568
rect 9967 30536 9973 30568
rect 9855 30495 9907 30522
rect 9855 30470 9861 30495
rect 9861 30470 9895 30495
rect 9895 30470 9907 30495
rect 9921 30495 9973 30522
rect 9921 30470 9933 30495
rect 9933 30470 9967 30495
rect 9967 30470 9973 30495
rect 9855 30422 9907 30456
rect 9921 30422 9973 30456
rect 9855 30404 9861 30422
rect 9861 30404 9907 30422
rect 9921 30404 9967 30422
rect 9967 30404 9973 30422
rect 9855 30338 9861 30390
rect 9861 30338 9907 30390
rect 9921 30338 9967 30390
rect 9967 30338 9973 30390
rect 9855 30271 9861 30323
rect 9861 30271 9907 30323
rect 9921 30271 9967 30323
rect 9967 30271 9973 30323
rect 9855 30204 9861 30256
rect 9861 30204 9907 30256
rect 9921 30204 9967 30256
rect 9967 30204 9973 30256
rect 9855 28714 9907 28720
rect 9855 28680 9861 28714
rect 9861 28680 9895 28714
rect 9895 28680 9907 28714
rect 9855 28668 9907 28680
rect 9921 28714 9973 28720
rect 9921 28680 9933 28714
rect 9933 28680 9967 28714
rect 9967 28680 9973 28714
rect 9921 28668 9973 28680
rect 9855 28641 9907 28654
rect 9855 28607 9861 28641
rect 9861 28607 9895 28641
rect 9895 28607 9907 28641
rect 9855 28602 9907 28607
rect 9921 28641 9973 28654
rect 9921 28607 9933 28641
rect 9933 28607 9967 28641
rect 9967 28607 9973 28641
rect 9921 28602 9973 28607
rect 9855 28568 9907 28588
rect 9855 28536 9861 28568
rect 9861 28536 9895 28568
rect 9895 28536 9907 28568
rect 9921 28568 9973 28588
rect 9921 28536 9933 28568
rect 9933 28536 9967 28568
rect 9967 28536 9973 28568
rect 9855 28495 9907 28522
rect 9855 28470 9861 28495
rect 9861 28470 9895 28495
rect 9895 28470 9907 28495
rect 9921 28495 9973 28522
rect 9921 28470 9933 28495
rect 9933 28470 9967 28495
rect 9967 28470 9973 28495
rect 9855 28422 9907 28456
rect 9921 28422 9973 28456
rect 9855 28404 9861 28422
rect 9861 28404 9907 28422
rect 9921 28404 9967 28422
rect 9967 28404 9973 28422
rect 9855 28338 9861 28390
rect 9861 28338 9907 28390
rect 9921 28338 9967 28390
rect 9967 28338 9973 28390
rect 9855 28271 9861 28323
rect 9861 28271 9907 28323
rect 9921 28271 9967 28323
rect 9967 28271 9973 28323
rect 9855 28204 9861 28256
rect 9861 28204 9907 28256
rect 9921 28204 9967 28256
rect 9967 28204 9973 28256
rect 9855 26717 9861 26720
rect 9861 26717 9895 26720
rect 9895 26717 9907 26720
rect 9855 26676 9907 26717
rect 9855 26668 9861 26676
rect 9861 26668 9895 26676
rect 9895 26668 9907 26676
rect 9921 26717 9933 26720
rect 9933 26717 9967 26720
rect 9967 26717 9973 26720
rect 9921 26676 9973 26717
rect 9921 26668 9933 26676
rect 9933 26668 9967 26676
rect 9967 26668 9973 26676
rect 9855 26642 9861 26654
rect 9861 26642 9895 26654
rect 9895 26642 9907 26654
rect 9855 26602 9907 26642
rect 9921 26642 9933 26654
rect 9933 26642 9967 26654
rect 9967 26642 9973 26654
rect 9921 26602 9973 26642
rect 9855 26567 9861 26588
rect 9861 26567 9895 26588
rect 9895 26567 9907 26588
rect 9855 26536 9907 26567
rect 9921 26567 9933 26588
rect 9933 26567 9967 26588
rect 9967 26567 9973 26588
rect 9921 26536 9973 26567
rect 9855 26492 9861 26522
rect 9861 26492 9895 26522
rect 9895 26492 9907 26522
rect 9855 26470 9907 26492
rect 9921 26492 9933 26522
rect 9933 26492 9967 26522
rect 9967 26492 9973 26522
rect 9921 26470 9973 26492
rect 9855 26451 9907 26456
rect 9855 26417 9861 26451
rect 9861 26417 9895 26451
rect 9895 26417 9907 26451
rect 9855 26404 9907 26417
rect 9921 26451 9973 26456
rect 9921 26417 9933 26451
rect 9933 26417 9967 26451
rect 9967 26417 9973 26451
rect 9921 26404 9973 26417
rect 9855 26376 9907 26389
rect 9855 26342 9861 26376
rect 9861 26342 9895 26376
rect 9895 26342 9907 26376
rect 9855 26337 9907 26342
rect 9921 26376 9973 26389
rect 9921 26342 9933 26376
rect 9933 26342 9967 26376
rect 9967 26342 9973 26376
rect 9921 26337 9973 26342
rect 9855 26301 9907 26322
rect 9855 26270 9861 26301
rect 9861 26270 9895 26301
rect 9895 26270 9907 26301
rect 9921 26301 9973 26322
rect 9921 26270 9933 26301
rect 9933 26270 9967 26301
rect 9967 26270 9973 26301
rect 9855 26226 9907 26255
rect 9855 26203 9861 26226
rect 9861 26203 9895 26226
rect 9895 26203 9907 26226
rect 9921 26226 9973 26255
rect 9921 26203 9933 26226
rect 9933 26203 9967 26226
rect 9967 26203 9973 26226
rect 10273 33840 10279 33892
rect 10279 33840 10325 33892
rect 10339 33840 10385 33892
rect 10385 33840 10391 33892
rect 10273 33774 10279 33826
rect 10279 33774 10325 33826
rect 10339 33774 10385 33826
rect 10385 33774 10391 33826
rect 10273 33708 10279 33760
rect 10279 33708 10325 33760
rect 10339 33708 10385 33760
rect 10385 33708 10391 33760
rect 10273 33642 10279 33694
rect 10279 33642 10325 33694
rect 10339 33642 10385 33694
rect 10385 33642 10391 33694
rect 10273 33575 10279 33627
rect 10279 33575 10325 33627
rect 10339 33575 10385 33627
rect 10385 33575 10391 33627
rect 10273 33508 10279 33560
rect 10279 33508 10325 33560
rect 10339 33508 10385 33560
rect 10385 33508 10391 33560
rect 10273 33441 10279 33493
rect 10279 33441 10325 33493
rect 10339 33441 10385 33493
rect 10385 33441 10391 33493
rect 10273 33380 10279 33426
rect 10279 33380 10325 33426
rect 10339 33380 10385 33426
rect 10385 33380 10391 33426
rect 10273 33374 10325 33380
rect 10339 33374 10391 33380
rect 10273 31840 10279 31892
rect 10279 31840 10325 31892
rect 10339 31840 10385 31892
rect 10385 31840 10391 31892
rect 10273 31774 10279 31826
rect 10279 31774 10325 31826
rect 10339 31774 10385 31826
rect 10385 31774 10391 31826
rect 10273 31708 10279 31760
rect 10279 31708 10325 31760
rect 10339 31708 10385 31760
rect 10385 31708 10391 31760
rect 10273 31642 10279 31694
rect 10279 31642 10325 31694
rect 10339 31642 10385 31694
rect 10385 31642 10391 31694
rect 10273 31575 10279 31627
rect 10279 31575 10325 31627
rect 10339 31575 10385 31627
rect 10385 31575 10391 31627
rect 10273 31508 10279 31560
rect 10279 31508 10325 31560
rect 10339 31508 10385 31560
rect 10385 31508 10391 31560
rect 10273 31441 10279 31493
rect 10279 31441 10325 31493
rect 10339 31441 10385 31493
rect 10385 31441 10391 31493
rect 10273 31380 10279 31426
rect 10279 31380 10325 31426
rect 10339 31380 10385 31426
rect 10385 31380 10391 31426
rect 10273 31374 10325 31380
rect 10339 31374 10391 31380
rect 10273 29840 10279 29892
rect 10279 29840 10325 29892
rect 10339 29840 10385 29892
rect 10385 29840 10391 29892
rect 10273 29774 10279 29826
rect 10279 29774 10325 29826
rect 10339 29774 10385 29826
rect 10385 29774 10391 29826
rect 10273 29708 10279 29760
rect 10279 29708 10325 29760
rect 10339 29708 10385 29760
rect 10385 29708 10391 29760
rect 10273 29642 10279 29694
rect 10279 29642 10325 29694
rect 10339 29642 10385 29694
rect 10385 29642 10391 29694
rect 10273 29575 10279 29627
rect 10279 29575 10325 29627
rect 10339 29575 10385 29627
rect 10385 29575 10391 29627
rect 10273 29508 10279 29560
rect 10279 29508 10325 29560
rect 10339 29508 10385 29560
rect 10385 29508 10391 29560
rect 10273 29441 10279 29493
rect 10279 29441 10325 29493
rect 10339 29441 10385 29493
rect 10385 29441 10391 29493
rect 10273 29380 10279 29426
rect 10279 29380 10325 29426
rect 10339 29380 10385 29426
rect 10385 29380 10391 29426
rect 10273 29374 10325 29380
rect 10339 29374 10391 29380
rect 10273 27840 10279 27892
rect 10279 27840 10325 27892
rect 10339 27840 10385 27892
rect 10385 27840 10391 27892
rect 10273 27774 10279 27826
rect 10279 27774 10325 27826
rect 10339 27774 10385 27826
rect 10385 27774 10391 27826
rect 10273 27708 10279 27760
rect 10279 27708 10325 27760
rect 10339 27708 10385 27760
rect 10385 27708 10391 27760
rect 10273 27642 10279 27694
rect 10279 27642 10325 27694
rect 10339 27642 10385 27694
rect 10385 27642 10391 27694
rect 10273 27575 10279 27627
rect 10279 27575 10325 27627
rect 10339 27575 10385 27627
rect 10385 27575 10391 27627
rect 10273 27508 10279 27560
rect 10279 27508 10325 27560
rect 10339 27508 10385 27560
rect 10385 27508 10391 27560
rect 10273 27441 10279 27493
rect 10279 27441 10325 27493
rect 10339 27441 10385 27493
rect 10385 27441 10391 27493
rect 10273 27380 10279 27426
rect 10279 27380 10325 27426
rect 10339 27380 10385 27426
rect 10385 27380 10391 27426
rect 10273 27374 10325 27380
rect 10339 27374 10391 27380
rect 10273 25857 10325 25891
rect 10273 25839 10279 25857
rect 10279 25839 10313 25857
rect 10313 25839 10325 25857
rect 10339 25857 10391 25891
rect 10339 25839 10351 25857
rect 10351 25839 10385 25857
rect 10385 25839 10391 25857
rect 10273 25823 10279 25825
rect 10279 25823 10313 25825
rect 10313 25823 10325 25825
rect 10273 25780 10325 25823
rect 10273 25773 10279 25780
rect 10279 25773 10313 25780
rect 10313 25773 10325 25780
rect 10339 25823 10351 25825
rect 10351 25823 10385 25825
rect 10385 25823 10391 25825
rect 10339 25780 10391 25823
rect 10339 25773 10351 25780
rect 10351 25773 10385 25780
rect 10385 25773 10391 25780
rect 10273 25746 10279 25759
rect 10279 25746 10313 25759
rect 10313 25746 10325 25759
rect 9437 25641 9489 25693
rect 9503 25641 9555 25693
rect 9437 25574 9489 25626
rect 9503 25574 9555 25626
rect 9437 25507 9489 25559
rect 9503 25507 9555 25559
rect 9437 25440 9489 25492
rect 9503 25440 9555 25492
rect 9437 25373 9489 25425
rect 9503 25373 9555 25425
rect 10273 25707 10325 25746
rect 10339 25746 10351 25759
rect 10351 25746 10385 25759
rect 10385 25746 10391 25759
rect 10339 25707 10391 25746
rect 10691 34714 10743 34720
rect 10691 34680 10697 34714
rect 10697 34680 10731 34714
rect 10731 34680 10743 34714
rect 10691 34668 10743 34680
rect 10757 34714 10809 34720
rect 10757 34680 10769 34714
rect 10769 34680 10803 34714
rect 10803 34680 10809 34714
rect 10757 34668 10809 34680
rect 10691 34641 10743 34654
rect 10691 34607 10697 34641
rect 10697 34607 10731 34641
rect 10731 34607 10743 34641
rect 10691 34602 10743 34607
rect 10757 34641 10809 34654
rect 10757 34607 10769 34641
rect 10769 34607 10803 34641
rect 10803 34607 10809 34641
rect 10757 34602 10809 34607
rect 10691 34568 10743 34588
rect 10691 34536 10697 34568
rect 10697 34536 10731 34568
rect 10731 34536 10743 34568
rect 10757 34568 10809 34588
rect 10757 34536 10769 34568
rect 10769 34536 10803 34568
rect 10803 34536 10809 34568
rect 10691 34495 10743 34522
rect 10691 34470 10697 34495
rect 10697 34470 10731 34495
rect 10731 34470 10743 34495
rect 10757 34495 10809 34522
rect 10757 34470 10769 34495
rect 10769 34470 10803 34495
rect 10803 34470 10809 34495
rect 10691 34422 10743 34456
rect 10757 34422 10809 34456
rect 10691 34404 10697 34422
rect 10697 34404 10743 34422
rect 10757 34404 10803 34422
rect 10803 34404 10809 34422
rect 10691 34338 10697 34390
rect 10697 34338 10743 34390
rect 10757 34338 10803 34390
rect 10803 34338 10809 34390
rect 10691 34271 10697 34323
rect 10697 34271 10743 34323
rect 10757 34271 10803 34323
rect 10803 34271 10809 34323
rect 10691 34204 10697 34256
rect 10697 34204 10743 34256
rect 10757 34204 10803 34256
rect 10803 34204 10809 34256
rect 10691 32714 10743 32720
rect 10691 32680 10697 32714
rect 10697 32680 10731 32714
rect 10731 32680 10743 32714
rect 10691 32668 10743 32680
rect 10757 32714 10809 32720
rect 10757 32680 10769 32714
rect 10769 32680 10803 32714
rect 10803 32680 10809 32714
rect 10757 32668 10809 32680
rect 10691 32641 10743 32654
rect 10691 32607 10697 32641
rect 10697 32607 10731 32641
rect 10731 32607 10743 32641
rect 10691 32602 10743 32607
rect 10757 32641 10809 32654
rect 10757 32607 10769 32641
rect 10769 32607 10803 32641
rect 10803 32607 10809 32641
rect 10757 32602 10809 32607
rect 10691 32568 10743 32588
rect 10691 32536 10697 32568
rect 10697 32536 10731 32568
rect 10731 32536 10743 32568
rect 10757 32568 10809 32588
rect 10757 32536 10769 32568
rect 10769 32536 10803 32568
rect 10803 32536 10809 32568
rect 10691 32495 10743 32522
rect 10691 32470 10697 32495
rect 10697 32470 10731 32495
rect 10731 32470 10743 32495
rect 10757 32495 10809 32522
rect 10757 32470 10769 32495
rect 10769 32470 10803 32495
rect 10803 32470 10809 32495
rect 10691 32422 10743 32456
rect 10757 32422 10809 32456
rect 10691 32404 10697 32422
rect 10697 32404 10743 32422
rect 10757 32404 10803 32422
rect 10803 32404 10809 32422
rect 10691 32338 10697 32390
rect 10697 32338 10743 32390
rect 10757 32338 10803 32390
rect 10803 32338 10809 32390
rect 10691 32271 10697 32323
rect 10697 32271 10743 32323
rect 10757 32271 10803 32323
rect 10803 32271 10809 32323
rect 10691 32204 10697 32256
rect 10697 32204 10743 32256
rect 10757 32204 10803 32256
rect 10803 32204 10809 32256
rect 10691 30714 10743 30720
rect 10691 30680 10697 30714
rect 10697 30680 10731 30714
rect 10731 30680 10743 30714
rect 10691 30668 10743 30680
rect 10757 30714 10809 30720
rect 10757 30680 10769 30714
rect 10769 30680 10803 30714
rect 10803 30680 10809 30714
rect 10757 30668 10809 30680
rect 10691 30641 10743 30654
rect 10691 30607 10697 30641
rect 10697 30607 10731 30641
rect 10731 30607 10743 30641
rect 10691 30602 10743 30607
rect 10757 30641 10809 30654
rect 10757 30607 10769 30641
rect 10769 30607 10803 30641
rect 10803 30607 10809 30641
rect 10757 30602 10809 30607
rect 10691 30568 10743 30588
rect 10691 30536 10697 30568
rect 10697 30536 10731 30568
rect 10731 30536 10743 30568
rect 10757 30568 10809 30588
rect 10757 30536 10769 30568
rect 10769 30536 10803 30568
rect 10803 30536 10809 30568
rect 10691 30495 10743 30522
rect 10691 30470 10697 30495
rect 10697 30470 10731 30495
rect 10731 30470 10743 30495
rect 10757 30495 10809 30522
rect 10757 30470 10769 30495
rect 10769 30470 10803 30495
rect 10803 30470 10809 30495
rect 10691 30422 10743 30456
rect 10757 30422 10809 30456
rect 10691 30404 10697 30422
rect 10697 30404 10743 30422
rect 10757 30404 10803 30422
rect 10803 30404 10809 30422
rect 10691 30338 10697 30390
rect 10697 30338 10743 30390
rect 10757 30338 10803 30390
rect 10803 30338 10809 30390
rect 10691 30271 10697 30323
rect 10697 30271 10743 30323
rect 10757 30271 10803 30323
rect 10803 30271 10809 30323
rect 10691 30204 10697 30256
rect 10697 30204 10743 30256
rect 10757 30204 10803 30256
rect 10803 30204 10809 30256
rect 10691 28714 10743 28720
rect 10691 28680 10697 28714
rect 10697 28680 10731 28714
rect 10731 28680 10743 28714
rect 10691 28668 10743 28680
rect 10757 28714 10809 28720
rect 10757 28680 10769 28714
rect 10769 28680 10803 28714
rect 10803 28680 10809 28714
rect 10757 28668 10809 28680
rect 10691 28641 10743 28654
rect 10691 28607 10697 28641
rect 10697 28607 10731 28641
rect 10731 28607 10743 28641
rect 10691 28602 10743 28607
rect 10757 28641 10809 28654
rect 10757 28607 10769 28641
rect 10769 28607 10803 28641
rect 10803 28607 10809 28641
rect 10757 28602 10809 28607
rect 10691 28568 10743 28588
rect 10691 28536 10697 28568
rect 10697 28536 10731 28568
rect 10731 28536 10743 28568
rect 10757 28568 10809 28588
rect 10757 28536 10769 28568
rect 10769 28536 10803 28568
rect 10803 28536 10809 28568
rect 10691 28495 10743 28522
rect 10691 28470 10697 28495
rect 10697 28470 10731 28495
rect 10731 28470 10743 28495
rect 10757 28495 10809 28522
rect 10757 28470 10769 28495
rect 10769 28470 10803 28495
rect 10803 28470 10809 28495
rect 10691 28422 10743 28456
rect 10757 28422 10809 28456
rect 10691 28404 10697 28422
rect 10697 28404 10743 28422
rect 10757 28404 10803 28422
rect 10803 28404 10809 28422
rect 10691 28338 10697 28390
rect 10697 28338 10743 28390
rect 10757 28338 10803 28390
rect 10803 28338 10809 28390
rect 10691 28271 10697 28323
rect 10697 28271 10743 28323
rect 10757 28271 10803 28323
rect 10803 28271 10809 28323
rect 10691 28204 10697 28256
rect 10697 28204 10743 28256
rect 10757 28204 10803 28256
rect 10803 28204 10809 28256
rect 10691 26717 10697 26720
rect 10697 26717 10731 26720
rect 10731 26717 10743 26720
rect 10691 26676 10743 26717
rect 10691 26668 10697 26676
rect 10697 26668 10731 26676
rect 10731 26668 10743 26676
rect 10757 26717 10769 26720
rect 10769 26717 10803 26720
rect 10803 26717 10809 26720
rect 10757 26676 10809 26717
rect 10757 26668 10769 26676
rect 10769 26668 10803 26676
rect 10803 26668 10809 26676
rect 10691 26642 10697 26654
rect 10697 26642 10731 26654
rect 10731 26642 10743 26654
rect 10691 26602 10743 26642
rect 10757 26642 10769 26654
rect 10769 26642 10803 26654
rect 10803 26642 10809 26654
rect 10757 26602 10809 26642
rect 10691 26567 10697 26588
rect 10697 26567 10731 26588
rect 10731 26567 10743 26588
rect 10691 26536 10743 26567
rect 10757 26567 10769 26588
rect 10769 26567 10803 26588
rect 10803 26567 10809 26588
rect 10757 26536 10809 26567
rect 10691 26492 10697 26522
rect 10697 26492 10731 26522
rect 10731 26492 10743 26522
rect 10691 26470 10743 26492
rect 10757 26492 10769 26522
rect 10769 26492 10803 26522
rect 10803 26492 10809 26522
rect 10757 26470 10809 26492
rect 10691 26451 10743 26456
rect 10691 26417 10697 26451
rect 10697 26417 10731 26451
rect 10731 26417 10743 26451
rect 10691 26404 10743 26417
rect 10757 26451 10809 26456
rect 10757 26417 10769 26451
rect 10769 26417 10803 26451
rect 10803 26417 10809 26451
rect 10757 26404 10809 26417
rect 10691 26376 10743 26389
rect 10691 26342 10697 26376
rect 10697 26342 10731 26376
rect 10731 26342 10743 26376
rect 10691 26337 10743 26342
rect 10757 26376 10809 26389
rect 10757 26342 10769 26376
rect 10769 26342 10803 26376
rect 10803 26342 10809 26376
rect 10757 26337 10809 26342
rect 10691 26301 10743 26322
rect 10691 26270 10697 26301
rect 10697 26270 10731 26301
rect 10731 26270 10743 26301
rect 10757 26301 10809 26322
rect 10757 26270 10769 26301
rect 10769 26270 10803 26301
rect 10803 26270 10809 26301
rect 10691 26226 10743 26255
rect 10691 26203 10697 26226
rect 10697 26203 10731 26226
rect 10731 26203 10743 26226
rect 10757 26226 10809 26255
rect 10757 26203 10769 26226
rect 10769 26203 10803 26226
rect 10803 26203 10809 26226
rect 11109 33840 11115 33892
rect 11115 33840 11161 33892
rect 11175 33840 11221 33892
rect 11221 33840 11227 33892
rect 11109 33774 11115 33826
rect 11115 33774 11161 33826
rect 11175 33774 11221 33826
rect 11221 33774 11227 33826
rect 11109 33708 11115 33760
rect 11115 33708 11161 33760
rect 11175 33708 11221 33760
rect 11221 33708 11227 33760
rect 11109 33642 11115 33694
rect 11115 33642 11161 33694
rect 11175 33642 11221 33694
rect 11221 33642 11227 33694
rect 11109 33575 11115 33627
rect 11115 33575 11161 33627
rect 11175 33575 11221 33627
rect 11221 33575 11227 33627
rect 11109 33508 11115 33560
rect 11115 33508 11161 33560
rect 11175 33508 11221 33560
rect 11221 33508 11227 33560
rect 11109 33441 11115 33493
rect 11115 33441 11161 33493
rect 11175 33441 11221 33493
rect 11221 33441 11227 33493
rect 11109 33380 11115 33426
rect 11115 33380 11161 33426
rect 11175 33380 11221 33426
rect 11221 33380 11227 33426
rect 11109 33374 11161 33380
rect 11175 33374 11227 33380
rect 11109 31840 11115 31892
rect 11115 31840 11161 31892
rect 11175 31840 11221 31892
rect 11221 31840 11227 31892
rect 11109 31774 11115 31826
rect 11115 31774 11161 31826
rect 11175 31774 11221 31826
rect 11221 31774 11227 31826
rect 11109 31708 11115 31760
rect 11115 31708 11161 31760
rect 11175 31708 11221 31760
rect 11221 31708 11227 31760
rect 11109 31642 11115 31694
rect 11115 31642 11161 31694
rect 11175 31642 11221 31694
rect 11221 31642 11227 31694
rect 11109 31575 11115 31627
rect 11115 31575 11161 31627
rect 11175 31575 11221 31627
rect 11221 31575 11227 31627
rect 11109 31508 11115 31560
rect 11115 31508 11161 31560
rect 11175 31508 11221 31560
rect 11221 31508 11227 31560
rect 11109 31441 11115 31493
rect 11115 31441 11161 31493
rect 11175 31441 11221 31493
rect 11221 31441 11227 31493
rect 11109 31380 11115 31426
rect 11115 31380 11161 31426
rect 11175 31380 11221 31426
rect 11221 31380 11227 31426
rect 11109 31374 11161 31380
rect 11175 31374 11227 31380
rect 11109 29840 11115 29892
rect 11115 29840 11161 29892
rect 11175 29840 11221 29892
rect 11221 29840 11227 29892
rect 11109 29774 11115 29826
rect 11115 29774 11161 29826
rect 11175 29774 11221 29826
rect 11221 29774 11227 29826
rect 11109 29708 11115 29760
rect 11115 29708 11161 29760
rect 11175 29708 11221 29760
rect 11221 29708 11227 29760
rect 11109 29642 11115 29694
rect 11115 29642 11161 29694
rect 11175 29642 11221 29694
rect 11221 29642 11227 29694
rect 11109 29575 11115 29627
rect 11115 29575 11161 29627
rect 11175 29575 11221 29627
rect 11221 29575 11227 29627
rect 11109 29508 11115 29560
rect 11115 29508 11161 29560
rect 11175 29508 11221 29560
rect 11221 29508 11227 29560
rect 11109 29441 11115 29493
rect 11115 29441 11161 29493
rect 11175 29441 11221 29493
rect 11221 29441 11227 29493
rect 11109 29380 11115 29426
rect 11115 29380 11161 29426
rect 11175 29380 11221 29426
rect 11221 29380 11227 29426
rect 11109 29374 11161 29380
rect 11175 29374 11227 29380
rect 11109 27840 11115 27892
rect 11115 27840 11161 27892
rect 11175 27840 11221 27892
rect 11221 27840 11227 27892
rect 11109 27774 11115 27826
rect 11115 27774 11161 27826
rect 11175 27774 11221 27826
rect 11221 27774 11227 27826
rect 11109 27708 11115 27760
rect 11115 27708 11161 27760
rect 11175 27708 11221 27760
rect 11221 27708 11227 27760
rect 11109 27642 11115 27694
rect 11115 27642 11161 27694
rect 11175 27642 11221 27694
rect 11221 27642 11227 27694
rect 11109 27575 11115 27627
rect 11115 27575 11161 27627
rect 11175 27575 11221 27627
rect 11221 27575 11227 27627
rect 11109 27508 11115 27560
rect 11115 27508 11161 27560
rect 11175 27508 11221 27560
rect 11221 27508 11227 27560
rect 11109 27441 11115 27493
rect 11115 27441 11161 27493
rect 11175 27441 11221 27493
rect 11221 27441 11227 27493
rect 11109 27380 11115 27426
rect 11115 27380 11161 27426
rect 11175 27380 11221 27426
rect 11221 27380 11227 27426
rect 11109 27374 11161 27380
rect 11175 27374 11227 27380
rect 11109 25857 11161 25891
rect 11109 25839 11115 25857
rect 11115 25839 11149 25857
rect 11149 25839 11161 25857
rect 11175 25857 11227 25891
rect 11175 25839 11187 25857
rect 11187 25839 11221 25857
rect 11221 25839 11227 25857
rect 11109 25823 11115 25825
rect 11115 25823 11149 25825
rect 11149 25823 11161 25825
rect 11109 25780 11161 25823
rect 11109 25773 11115 25780
rect 11115 25773 11149 25780
rect 11149 25773 11161 25780
rect 11175 25823 11187 25825
rect 11187 25823 11221 25825
rect 11221 25823 11227 25825
rect 11175 25780 11227 25823
rect 11175 25773 11187 25780
rect 11187 25773 11221 25780
rect 11221 25773 11227 25780
rect 11109 25746 11115 25759
rect 11115 25746 11149 25759
rect 11149 25746 11161 25759
rect 10273 25641 10325 25693
rect 10339 25641 10391 25693
rect 10273 25574 10325 25626
rect 10339 25574 10391 25626
rect 10273 25507 10325 25559
rect 10339 25507 10391 25559
rect 10273 25440 10325 25492
rect 10339 25440 10391 25492
rect 10273 25373 10325 25425
rect 10339 25373 10391 25425
rect 11109 25707 11161 25746
rect 11175 25746 11187 25759
rect 11187 25746 11221 25759
rect 11221 25746 11227 25759
rect 11175 25707 11227 25746
rect 11527 34714 11579 34720
rect 11527 34680 11533 34714
rect 11533 34680 11567 34714
rect 11567 34680 11579 34714
rect 11527 34668 11579 34680
rect 11593 34714 11645 34720
rect 11593 34680 11605 34714
rect 11605 34680 11639 34714
rect 11639 34680 11645 34714
rect 11593 34668 11645 34680
rect 11527 34641 11579 34654
rect 11527 34607 11533 34641
rect 11533 34607 11567 34641
rect 11567 34607 11579 34641
rect 11527 34602 11579 34607
rect 11593 34641 11645 34654
rect 11593 34607 11605 34641
rect 11605 34607 11639 34641
rect 11639 34607 11645 34641
rect 11593 34602 11645 34607
rect 11527 34568 11579 34588
rect 11527 34536 11533 34568
rect 11533 34536 11567 34568
rect 11567 34536 11579 34568
rect 11593 34568 11645 34588
rect 11593 34536 11605 34568
rect 11605 34536 11639 34568
rect 11639 34536 11645 34568
rect 11527 34495 11579 34522
rect 11527 34470 11533 34495
rect 11533 34470 11567 34495
rect 11567 34470 11579 34495
rect 11593 34495 11645 34522
rect 11593 34470 11605 34495
rect 11605 34470 11639 34495
rect 11639 34470 11645 34495
rect 11527 34422 11579 34456
rect 11593 34422 11645 34456
rect 11527 34404 11533 34422
rect 11533 34404 11579 34422
rect 11593 34404 11639 34422
rect 11639 34404 11645 34422
rect 11527 34338 11533 34390
rect 11533 34338 11579 34390
rect 11593 34338 11639 34390
rect 11639 34338 11645 34390
rect 11527 34271 11533 34323
rect 11533 34271 11579 34323
rect 11593 34271 11639 34323
rect 11639 34271 11645 34323
rect 11527 34204 11533 34256
rect 11533 34204 11579 34256
rect 11593 34204 11639 34256
rect 11639 34204 11645 34256
rect 11527 32714 11579 32720
rect 11527 32680 11533 32714
rect 11533 32680 11567 32714
rect 11567 32680 11579 32714
rect 11527 32668 11579 32680
rect 11593 32714 11645 32720
rect 11593 32680 11605 32714
rect 11605 32680 11639 32714
rect 11639 32680 11645 32714
rect 11593 32668 11645 32680
rect 11527 32641 11579 32654
rect 11527 32607 11533 32641
rect 11533 32607 11567 32641
rect 11567 32607 11579 32641
rect 11527 32602 11579 32607
rect 11593 32641 11645 32654
rect 11593 32607 11605 32641
rect 11605 32607 11639 32641
rect 11639 32607 11645 32641
rect 11593 32602 11645 32607
rect 11527 32568 11579 32588
rect 11527 32536 11533 32568
rect 11533 32536 11567 32568
rect 11567 32536 11579 32568
rect 11593 32568 11645 32588
rect 11593 32536 11605 32568
rect 11605 32536 11639 32568
rect 11639 32536 11645 32568
rect 11527 32495 11579 32522
rect 11527 32470 11533 32495
rect 11533 32470 11567 32495
rect 11567 32470 11579 32495
rect 11593 32495 11645 32522
rect 11593 32470 11605 32495
rect 11605 32470 11639 32495
rect 11639 32470 11645 32495
rect 11527 32422 11579 32456
rect 11593 32422 11645 32456
rect 11527 32404 11533 32422
rect 11533 32404 11579 32422
rect 11593 32404 11639 32422
rect 11639 32404 11645 32422
rect 11527 32338 11533 32390
rect 11533 32338 11579 32390
rect 11593 32338 11639 32390
rect 11639 32338 11645 32390
rect 11527 32271 11533 32323
rect 11533 32271 11579 32323
rect 11593 32271 11639 32323
rect 11639 32271 11645 32323
rect 11527 32204 11533 32256
rect 11533 32204 11579 32256
rect 11593 32204 11639 32256
rect 11639 32204 11645 32256
rect 11527 30714 11579 30720
rect 11527 30680 11533 30714
rect 11533 30680 11567 30714
rect 11567 30680 11579 30714
rect 11527 30668 11579 30680
rect 11593 30714 11645 30720
rect 11593 30680 11605 30714
rect 11605 30680 11639 30714
rect 11639 30680 11645 30714
rect 11593 30668 11645 30680
rect 11527 30641 11579 30654
rect 11527 30607 11533 30641
rect 11533 30607 11567 30641
rect 11567 30607 11579 30641
rect 11527 30602 11579 30607
rect 11593 30641 11645 30654
rect 11593 30607 11605 30641
rect 11605 30607 11639 30641
rect 11639 30607 11645 30641
rect 11593 30602 11645 30607
rect 11527 30568 11579 30588
rect 11527 30536 11533 30568
rect 11533 30536 11567 30568
rect 11567 30536 11579 30568
rect 11593 30568 11645 30588
rect 11593 30536 11605 30568
rect 11605 30536 11639 30568
rect 11639 30536 11645 30568
rect 11527 30495 11579 30522
rect 11527 30470 11533 30495
rect 11533 30470 11567 30495
rect 11567 30470 11579 30495
rect 11593 30495 11645 30522
rect 11593 30470 11605 30495
rect 11605 30470 11639 30495
rect 11639 30470 11645 30495
rect 11527 30422 11579 30456
rect 11593 30422 11645 30456
rect 11527 30404 11533 30422
rect 11533 30404 11579 30422
rect 11593 30404 11639 30422
rect 11639 30404 11645 30422
rect 11527 30338 11533 30390
rect 11533 30338 11579 30390
rect 11593 30338 11639 30390
rect 11639 30338 11645 30390
rect 11527 30271 11533 30323
rect 11533 30271 11579 30323
rect 11593 30271 11639 30323
rect 11639 30271 11645 30323
rect 11527 30204 11533 30256
rect 11533 30204 11579 30256
rect 11593 30204 11639 30256
rect 11639 30204 11645 30256
rect 11527 28714 11579 28720
rect 11527 28680 11533 28714
rect 11533 28680 11567 28714
rect 11567 28680 11579 28714
rect 11527 28668 11579 28680
rect 11593 28714 11645 28720
rect 11593 28680 11605 28714
rect 11605 28680 11639 28714
rect 11639 28680 11645 28714
rect 11593 28668 11645 28680
rect 11527 28641 11579 28654
rect 11527 28607 11533 28641
rect 11533 28607 11567 28641
rect 11567 28607 11579 28641
rect 11527 28602 11579 28607
rect 11593 28641 11645 28654
rect 11593 28607 11605 28641
rect 11605 28607 11639 28641
rect 11639 28607 11645 28641
rect 11593 28602 11645 28607
rect 11527 28568 11579 28588
rect 11527 28536 11533 28568
rect 11533 28536 11567 28568
rect 11567 28536 11579 28568
rect 11593 28568 11645 28588
rect 11593 28536 11605 28568
rect 11605 28536 11639 28568
rect 11639 28536 11645 28568
rect 11527 28495 11579 28522
rect 11527 28470 11533 28495
rect 11533 28470 11567 28495
rect 11567 28470 11579 28495
rect 11593 28495 11645 28522
rect 11593 28470 11605 28495
rect 11605 28470 11639 28495
rect 11639 28470 11645 28495
rect 11527 28422 11579 28456
rect 11593 28422 11645 28456
rect 11527 28404 11533 28422
rect 11533 28404 11579 28422
rect 11593 28404 11639 28422
rect 11639 28404 11645 28422
rect 11527 28338 11533 28390
rect 11533 28338 11579 28390
rect 11593 28338 11639 28390
rect 11639 28338 11645 28390
rect 11527 28271 11533 28323
rect 11533 28271 11579 28323
rect 11593 28271 11639 28323
rect 11639 28271 11645 28323
rect 11527 28204 11533 28256
rect 11533 28204 11579 28256
rect 11593 28204 11639 28256
rect 11639 28204 11645 28256
rect 11527 26717 11533 26720
rect 11533 26717 11567 26720
rect 11567 26717 11579 26720
rect 11527 26676 11579 26717
rect 11527 26668 11533 26676
rect 11533 26668 11567 26676
rect 11567 26668 11579 26676
rect 11593 26717 11605 26720
rect 11605 26717 11639 26720
rect 11639 26717 11645 26720
rect 11593 26676 11645 26717
rect 11593 26668 11605 26676
rect 11605 26668 11639 26676
rect 11639 26668 11645 26676
rect 11527 26642 11533 26654
rect 11533 26642 11567 26654
rect 11567 26642 11579 26654
rect 11527 26602 11579 26642
rect 11593 26642 11605 26654
rect 11605 26642 11639 26654
rect 11639 26642 11645 26654
rect 11593 26602 11645 26642
rect 11527 26567 11533 26588
rect 11533 26567 11567 26588
rect 11567 26567 11579 26588
rect 11527 26536 11579 26567
rect 11593 26567 11605 26588
rect 11605 26567 11639 26588
rect 11639 26567 11645 26588
rect 11593 26536 11645 26567
rect 11527 26492 11533 26522
rect 11533 26492 11567 26522
rect 11567 26492 11579 26522
rect 11527 26470 11579 26492
rect 11593 26492 11605 26522
rect 11605 26492 11639 26522
rect 11639 26492 11645 26522
rect 11593 26470 11645 26492
rect 11527 26451 11579 26456
rect 11527 26417 11533 26451
rect 11533 26417 11567 26451
rect 11567 26417 11579 26451
rect 11527 26404 11579 26417
rect 11593 26451 11645 26456
rect 11593 26417 11605 26451
rect 11605 26417 11639 26451
rect 11639 26417 11645 26451
rect 11593 26404 11645 26417
rect 11527 26376 11579 26389
rect 11527 26342 11533 26376
rect 11533 26342 11567 26376
rect 11567 26342 11579 26376
rect 11527 26337 11579 26342
rect 11593 26376 11645 26389
rect 11593 26342 11605 26376
rect 11605 26342 11639 26376
rect 11639 26342 11645 26376
rect 11593 26337 11645 26342
rect 11527 26301 11579 26322
rect 11527 26270 11533 26301
rect 11533 26270 11567 26301
rect 11567 26270 11579 26301
rect 11593 26301 11645 26322
rect 11593 26270 11605 26301
rect 11605 26270 11639 26301
rect 11639 26270 11645 26301
rect 11527 26226 11579 26255
rect 11527 26203 11533 26226
rect 11533 26203 11567 26226
rect 11567 26203 11579 26226
rect 11593 26226 11645 26255
rect 11593 26203 11605 26226
rect 11605 26203 11639 26226
rect 11639 26203 11645 26226
rect 11945 33840 11951 33892
rect 11951 33840 11997 33892
rect 12011 33840 12057 33892
rect 12057 33840 12063 33892
rect 11945 33774 11951 33826
rect 11951 33774 11997 33826
rect 12011 33774 12057 33826
rect 12057 33774 12063 33826
rect 11945 33708 11951 33760
rect 11951 33708 11997 33760
rect 12011 33708 12057 33760
rect 12057 33708 12063 33760
rect 11945 33642 11951 33694
rect 11951 33642 11997 33694
rect 12011 33642 12057 33694
rect 12057 33642 12063 33694
rect 11945 33575 11951 33627
rect 11951 33575 11997 33627
rect 12011 33575 12057 33627
rect 12057 33575 12063 33627
rect 11945 33508 11951 33560
rect 11951 33508 11997 33560
rect 12011 33508 12057 33560
rect 12057 33508 12063 33560
rect 11945 33441 11951 33493
rect 11951 33441 11997 33493
rect 12011 33441 12057 33493
rect 12057 33441 12063 33493
rect 11945 33380 11951 33426
rect 11951 33380 11997 33426
rect 12011 33380 12057 33426
rect 12057 33380 12063 33426
rect 11945 33374 11997 33380
rect 12011 33374 12063 33380
rect 11945 31840 11951 31892
rect 11951 31840 11997 31892
rect 12011 31840 12057 31892
rect 12057 31840 12063 31892
rect 11945 31774 11951 31826
rect 11951 31774 11997 31826
rect 12011 31774 12057 31826
rect 12057 31774 12063 31826
rect 11945 31708 11951 31760
rect 11951 31708 11997 31760
rect 12011 31708 12057 31760
rect 12057 31708 12063 31760
rect 11945 31642 11951 31694
rect 11951 31642 11997 31694
rect 12011 31642 12057 31694
rect 12057 31642 12063 31694
rect 11945 31575 11951 31627
rect 11951 31575 11997 31627
rect 12011 31575 12057 31627
rect 12057 31575 12063 31627
rect 11945 31508 11951 31560
rect 11951 31508 11997 31560
rect 12011 31508 12057 31560
rect 12057 31508 12063 31560
rect 11945 31441 11951 31493
rect 11951 31441 11997 31493
rect 12011 31441 12057 31493
rect 12057 31441 12063 31493
rect 11945 31380 11951 31426
rect 11951 31380 11997 31426
rect 12011 31380 12057 31426
rect 12057 31380 12063 31426
rect 11945 31374 11997 31380
rect 12011 31374 12063 31380
rect 11945 29840 11951 29892
rect 11951 29840 11997 29892
rect 12011 29840 12057 29892
rect 12057 29840 12063 29892
rect 11945 29774 11951 29826
rect 11951 29774 11997 29826
rect 12011 29774 12057 29826
rect 12057 29774 12063 29826
rect 11945 29708 11951 29760
rect 11951 29708 11997 29760
rect 12011 29708 12057 29760
rect 12057 29708 12063 29760
rect 11945 29642 11951 29694
rect 11951 29642 11997 29694
rect 12011 29642 12057 29694
rect 12057 29642 12063 29694
rect 11945 29575 11951 29627
rect 11951 29575 11997 29627
rect 12011 29575 12057 29627
rect 12057 29575 12063 29627
rect 11945 29508 11951 29560
rect 11951 29508 11997 29560
rect 12011 29508 12057 29560
rect 12057 29508 12063 29560
rect 11945 29441 11951 29493
rect 11951 29441 11997 29493
rect 12011 29441 12057 29493
rect 12057 29441 12063 29493
rect 11945 29380 11951 29426
rect 11951 29380 11997 29426
rect 12011 29380 12057 29426
rect 12057 29380 12063 29426
rect 11945 29374 11997 29380
rect 12011 29374 12063 29380
rect 11945 27840 11951 27892
rect 11951 27840 11997 27892
rect 12011 27840 12057 27892
rect 12057 27840 12063 27892
rect 11945 27774 11951 27826
rect 11951 27774 11997 27826
rect 12011 27774 12057 27826
rect 12057 27774 12063 27826
rect 11945 27708 11951 27760
rect 11951 27708 11997 27760
rect 12011 27708 12057 27760
rect 12057 27708 12063 27760
rect 11945 27642 11951 27694
rect 11951 27642 11997 27694
rect 12011 27642 12057 27694
rect 12057 27642 12063 27694
rect 11945 27575 11951 27627
rect 11951 27575 11997 27627
rect 12011 27575 12057 27627
rect 12057 27575 12063 27627
rect 11945 27508 11951 27560
rect 11951 27508 11997 27560
rect 12011 27508 12057 27560
rect 12057 27508 12063 27560
rect 11945 27441 11951 27493
rect 11951 27441 11997 27493
rect 12011 27441 12057 27493
rect 12057 27441 12063 27493
rect 11945 27380 11951 27426
rect 11951 27380 11997 27426
rect 12011 27380 12057 27426
rect 12057 27380 12063 27426
rect 11945 27374 11997 27380
rect 12011 27374 12063 27380
rect 11945 25857 11997 25891
rect 11945 25839 11951 25857
rect 11951 25839 11985 25857
rect 11985 25839 11997 25857
rect 12011 25857 12063 25891
rect 12011 25839 12023 25857
rect 12023 25839 12057 25857
rect 12057 25839 12063 25857
rect 11945 25823 11951 25825
rect 11951 25823 11985 25825
rect 11985 25823 11997 25825
rect 11945 25780 11997 25823
rect 11945 25773 11951 25780
rect 11951 25773 11985 25780
rect 11985 25773 11997 25780
rect 12011 25823 12023 25825
rect 12023 25823 12057 25825
rect 12057 25823 12063 25825
rect 12011 25780 12063 25823
rect 12011 25773 12023 25780
rect 12023 25773 12057 25780
rect 12057 25773 12063 25780
rect 11945 25746 11951 25759
rect 11951 25746 11985 25759
rect 11985 25746 11997 25759
rect 11109 25641 11161 25693
rect 11175 25641 11227 25693
rect 11109 25574 11161 25626
rect 11175 25574 11227 25626
rect 11109 25507 11161 25559
rect 11175 25507 11227 25559
rect 11109 25440 11161 25492
rect 11175 25440 11227 25492
rect 11109 25373 11161 25425
rect 11175 25373 11227 25425
rect 11945 25707 11997 25746
rect 12011 25746 12023 25759
rect 12023 25746 12057 25759
rect 12057 25746 12063 25759
rect 12011 25707 12063 25746
rect 12363 34714 12415 34720
rect 12363 34680 12369 34714
rect 12369 34680 12403 34714
rect 12403 34680 12415 34714
rect 12363 34668 12415 34680
rect 12429 34714 12481 34720
rect 12429 34680 12441 34714
rect 12441 34680 12475 34714
rect 12475 34680 12481 34714
rect 12429 34668 12481 34680
rect 12363 34641 12415 34654
rect 12363 34607 12369 34641
rect 12369 34607 12403 34641
rect 12403 34607 12415 34641
rect 12363 34602 12415 34607
rect 12429 34641 12481 34654
rect 12429 34607 12441 34641
rect 12441 34607 12475 34641
rect 12475 34607 12481 34641
rect 12429 34602 12481 34607
rect 12363 34568 12415 34588
rect 12363 34536 12369 34568
rect 12369 34536 12403 34568
rect 12403 34536 12415 34568
rect 12429 34568 12481 34588
rect 12429 34536 12441 34568
rect 12441 34536 12475 34568
rect 12475 34536 12481 34568
rect 12363 34495 12415 34522
rect 12363 34470 12369 34495
rect 12369 34470 12403 34495
rect 12403 34470 12415 34495
rect 12429 34495 12481 34522
rect 12429 34470 12441 34495
rect 12441 34470 12475 34495
rect 12475 34470 12481 34495
rect 12363 34422 12415 34456
rect 12429 34422 12481 34456
rect 12363 34404 12369 34422
rect 12369 34404 12415 34422
rect 12429 34404 12475 34422
rect 12475 34404 12481 34422
rect 12363 34338 12369 34390
rect 12369 34338 12415 34390
rect 12429 34338 12475 34390
rect 12475 34338 12481 34390
rect 12363 34271 12369 34323
rect 12369 34271 12415 34323
rect 12429 34271 12475 34323
rect 12475 34271 12481 34323
rect 12363 34204 12369 34256
rect 12369 34204 12415 34256
rect 12429 34204 12475 34256
rect 12475 34204 12481 34256
rect 12363 32714 12415 32720
rect 12363 32680 12369 32714
rect 12369 32680 12403 32714
rect 12403 32680 12415 32714
rect 12363 32668 12415 32680
rect 12429 32714 12481 32720
rect 12429 32680 12441 32714
rect 12441 32680 12475 32714
rect 12475 32680 12481 32714
rect 12429 32668 12481 32680
rect 12363 32641 12415 32654
rect 12363 32607 12369 32641
rect 12369 32607 12403 32641
rect 12403 32607 12415 32641
rect 12363 32602 12415 32607
rect 12429 32641 12481 32654
rect 12429 32607 12441 32641
rect 12441 32607 12475 32641
rect 12475 32607 12481 32641
rect 12429 32602 12481 32607
rect 12363 32568 12415 32588
rect 12363 32536 12369 32568
rect 12369 32536 12403 32568
rect 12403 32536 12415 32568
rect 12429 32568 12481 32588
rect 12429 32536 12441 32568
rect 12441 32536 12475 32568
rect 12475 32536 12481 32568
rect 12363 32495 12415 32522
rect 12363 32470 12369 32495
rect 12369 32470 12403 32495
rect 12403 32470 12415 32495
rect 12429 32495 12481 32522
rect 12429 32470 12441 32495
rect 12441 32470 12475 32495
rect 12475 32470 12481 32495
rect 12363 32422 12415 32456
rect 12429 32422 12481 32456
rect 12363 32404 12369 32422
rect 12369 32404 12415 32422
rect 12429 32404 12475 32422
rect 12475 32404 12481 32422
rect 12363 32338 12369 32390
rect 12369 32338 12415 32390
rect 12429 32338 12475 32390
rect 12475 32338 12481 32390
rect 12363 32271 12369 32323
rect 12369 32271 12415 32323
rect 12429 32271 12475 32323
rect 12475 32271 12481 32323
rect 12363 32204 12369 32256
rect 12369 32204 12415 32256
rect 12429 32204 12475 32256
rect 12475 32204 12481 32256
rect 12363 30714 12415 30720
rect 12363 30680 12369 30714
rect 12369 30680 12403 30714
rect 12403 30680 12415 30714
rect 12363 30668 12415 30680
rect 12429 30714 12481 30720
rect 12429 30680 12441 30714
rect 12441 30680 12475 30714
rect 12475 30680 12481 30714
rect 12429 30668 12481 30680
rect 12363 30641 12415 30654
rect 12363 30607 12369 30641
rect 12369 30607 12403 30641
rect 12403 30607 12415 30641
rect 12363 30602 12415 30607
rect 12429 30641 12481 30654
rect 12429 30607 12441 30641
rect 12441 30607 12475 30641
rect 12475 30607 12481 30641
rect 12429 30602 12481 30607
rect 12363 30568 12415 30588
rect 12363 30536 12369 30568
rect 12369 30536 12403 30568
rect 12403 30536 12415 30568
rect 12429 30568 12481 30588
rect 12429 30536 12441 30568
rect 12441 30536 12475 30568
rect 12475 30536 12481 30568
rect 12363 30495 12415 30522
rect 12363 30470 12369 30495
rect 12369 30470 12403 30495
rect 12403 30470 12415 30495
rect 12429 30495 12481 30522
rect 12429 30470 12441 30495
rect 12441 30470 12475 30495
rect 12475 30470 12481 30495
rect 12363 30422 12415 30456
rect 12429 30422 12481 30456
rect 12363 30404 12369 30422
rect 12369 30404 12415 30422
rect 12429 30404 12475 30422
rect 12475 30404 12481 30422
rect 12363 30338 12369 30390
rect 12369 30338 12415 30390
rect 12429 30338 12475 30390
rect 12475 30338 12481 30390
rect 12363 30271 12369 30323
rect 12369 30271 12415 30323
rect 12429 30271 12475 30323
rect 12475 30271 12481 30323
rect 12363 30204 12369 30256
rect 12369 30204 12415 30256
rect 12429 30204 12475 30256
rect 12475 30204 12481 30256
rect 12363 28714 12415 28720
rect 12363 28680 12369 28714
rect 12369 28680 12403 28714
rect 12403 28680 12415 28714
rect 12363 28668 12415 28680
rect 12429 28714 12481 28720
rect 12429 28680 12441 28714
rect 12441 28680 12475 28714
rect 12475 28680 12481 28714
rect 12429 28668 12481 28680
rect 12363 28641 12415 28654
rect 12363 28607 12369 28641
rect 12369 28607 12403 28641
rect 12403 28607 12415 28641
rect 12363 28602 12415 28607
rect 12429 28641 12481 28654
rect 12429 28607 12441 28641
rect 12441 28607 12475 28641
rect 12475 28607 12481 28641
rect 12429 28602 12481 28607
rect 12363 28568 12415 28588
rect 12363 28536 12369 28568
rect 12369 28536 12403 28568
rect 12403 28536 12415 28568
rect 12429 28568 12481 28588
rect 12429 28536 12441 28568
rect 12441 28536 12475 28568
rect 12475 28536 12481 28568
rect 12363 28495 12415 28522
rect 12363 28470 12369 28495
rect 12369 28470 12403 28495
rect 12403 28470 12415 28495
rect 12429 28495 12481 28522
rect 12429 28470 12441 28495
rect 12441 28470 12475 28495
rect 12475 28470 12481 28495
rect 12363 28422 12415 28456
rect 12429 28422 12481 28456
rect 12363 28404 12369 28422
rect 12369 28404 12415 28422
rect 12429 28404 12475 28422
rect 12475 28404 12481 28422
rect 12363 28338 12369 28390
rect 12369 28338 12415 28390
rect 12429 28338 12475 28390
rect 12475 28338 12481 28390
rect 12363 28271 12369 28323
rect 12369 28271 12415 28323
rect 12429 28271 12475 28323
rect 12475 28271 12481 28323
rect 12363 28204 12369 28256
rect 12369 28204 12415 28256
rect 12429 28204 12475 28256
rect 12475 28204 12481 28256
rect 12363 26717 12369 26720
rect 12369 26717 12403 26720
rect 12403 26717 12415 26720
rect 12363 26676 12415 26717
rect 12363 26668 12369 26676
rect 12369 26668 12403 26676
rect 12403 26668 12415 26676
rect 12429 26717 12441 26720
rect 12441 26717 12475 26720
rect 12475 26717 12481 26720
rect 12429 26676 12481 26717
rect 12429 26668 12441 26676
rect 12441 26668 12475 26676
rect 12475 26668 12481 26676
rect 12363 26642 12369 26654
rect 12369 26642 12403 26654
rect 12403 26642 12415 26654
rect 12363 26602 12415 26642
rect 12429 26642 12441 26654
rect 12441 26642 12475 26654
rect 12475 26642 12481 26654
rect 12429 26602 12481 26642
rect 12363 26567 12369 26588
rect 12369 26567 12403 26588
rect 12403 26567 12415 26588
rect 12363 26536 12415 26567
rect 12429 26567 12441 26588
rect 12441 26567 12475 26588
rect 12475 26567 12481 26588
rect 12429 26536 12481 26567
rect 12363 26492 12369 26522
rect 12369 26492 12403 26522
rect 12403 26492 12415 26522
rect 12363 26470 12415 26492
rect 12429 26492 12441 26522
rect 12441 26492 12475 26522
rect 12475 26492 12481 26522
rect 12429 26470 12481 26492
rect 12363 26451 12415 26456
rect 12363 26417 12369 26451
rect 12369 26417 12403 26451
rect 12403 26417 12415 26451
rect 12363 26404 12415 26417
rect 12429 26451 12481 26456
rect 12429 26417 12441 26451
rect 12441 26417 12475 26451
rect 12475 26417 12481 26451
rect 12429 26404 12481 26417
rect 12363 26376 12415 26389
rect 12363 26342 12369 26376
rect 12369 26342 12403 26376
rect 12403 26342 12415 26376
rect 12363 26337 12415 26342
rect 12429 26376 12481 26389
rect 12429 26342 12441 26376
rect 12441 26342 12475 26376
rect 12475 26342 12481 26376
rect 12429 26337 12481 26342
rect 12363 26301 12415 26322
rect 12363 26270 12369 26301
rect 12369 26270 12403 26301
rect 12403 26270 12415 26301
rect 12429 26301 12481 26322
rect 12429 26270 12441 26301
rect 12441 26270 12475 26301
rect 12475 26270 12481 26301
rect 12363 26226 12415 26255
rect 12363 26203 12369 26226
rect 12369 26203 12403 26226
rect 12403 26203 12415 26226
rect 12429 26226 12481 26255
rect 12429 26203 12441 26226
rect 12441 26203 12475 26226
rect 12475 26203 12481 26226
rect 12781 33840 12787 33892
rect 12787 33840 12833 33892
rect 12847 33840 12893 33892
rect 12893 33840 12899 33892
rect 12781 33774 12787 33826
rect 12787 33774 12833 33826
rect 12847 33774 12893 33826
rect 12893 33774 12899 33826
rect 12781 33708 12787 33760
rect 12787 33708 12833 33760
rect 12847 33708 12893 33760
rect 12893 33708 12899 33760
rect 12781 33642 12787 33694
rect 12787 33642 12833 33694
rect 12847 33642 12893 33694
rect 12893 33642 12899 33694
rect 12781 33575 12787 33627
rect 12787 33575 12833 33627
rect 12847 33575 12893 33627
rect 12893 33575 12899 33627
rect 12781 33508 12787 33560
rect 12787 33508 12833 33560
rect 12847 33508 12893 33560
rect 12893 33508 12899 33560
rect 12781 33441 12787 33493
rect 12787 33441 12833 33493
rect 12847 33441 12893 33493
rect 12893 33441 12899 33493
rect 12781 33380 12787 33426
rect 12787 33380 12833 33426
rect 12847 33380 12893 33426
rect 12893 33380 12899 33426
rect 12781 33374 12833 33380
rect 12847 33374 12899 33380
rect 12781 31840 12787 31892
rect 12787 31840 12833 31892
rect 12847 31840 12893 31892
rect 12893 31840 12899 31892
rect 12781 31774 12787 31826
rect 12787 31774 12833 31826
rect 12847 31774 12893 31826
rect 12893 31774 12899 31826
rect 12781 31708 12787 31760
rect 12787 31708 12833 31760
rect 12847 31708 12893 31760
rect 12893 31708 12899 31760
rect 12781 31642 12787 31694
rect 12787 31642 12833 31694
rect 12847 31642 12893 31694
rect 12893 31642 12899 31694
rect 12781 31575 12787 31627
rect 12787 31575 12833 31627
rect 12847 31575 12893 31627
rect 12893 31575 12899 31627
rect 12781 31508 12787 31560
rect 12787 31508 12833 31560
rect 12847 31508 12893 31560
rect 12893 31508 12899 31560
rect 12781 31441 12787 31493
rect 12787 31441 12833 31493
rect 12847 31441 12893 31493
rect 12893 31441 12899 31493
rect 12781 31380 12787 31426
rect 12787 31380 12833 31426
rect 12847 31380 12893 31426
rect 12893 31380 12899 31426
rect 12781 31374 12833 31380
rect 12847 31374 12899 31380
rect 12781 29840 12787 29892
rect 12787 29840 12833 29892
rect 12847 29840 12893 29892
rect 12893 29840 12899 29892
rect 12781 29774 12787 29826
rect 12787 29774 12833 29826
rect 12847 29774 12893 29826
rect 12893 29774 12899 29826
rect 12781 29708 12787 29760
rect 12787 29708 12833 29760
rect 12847 29708 12893 29760
rect 12893 29708 12899 29760
rect 12781 29642 12787 29694
rect 12787 29642 12833 29694
rect 12847 29642 12893 29694
rect 12893 29642 12899 29694
rect 12781 29575 12787 29627
rect 12787 29575 12833 29627
rect 12847 29575 12893 29627
rect 12893 29575 12899 29627
rect 12781 29508 12787 29560
rect 12787 29508 12833 29560
rect 12847 29508 12893 29560
rect 12893 29508 12899 29560
rect 12781 29441 12787 29493
rect 12787 29441 12833 29493
rect 12847 29441 12893 29493
rect 12893 29441 12899 29493
rect 12781 29380 12787 29426
rect 12787 29380 12833 29426
rect 12847 29380 12893 29426
rect 12893 29380 12899 29426
rect 12781 29374 12833 29380
rect 12847 29374 12899 29380
rect 12781 27840 12787 27892
rect 12787 27840 12833 27892
rect 12847 27840 12893 27892
rect 12893 27840 12899 27892
rect 12781 27774 12787 27826
rect 12787 27774 12833 27826
rect 12847 27774 12893 27826
rect 12893 27774 12899 27826
rect 12781 27708 12787 27760
rect 12787 27708 12833 27760
rect 12847 27708 12893 27760
rect 12893 27708 12899 27760
rect 12781 27642 12787 27694
rect 12787 27642 12833 27694
rect 12847 27642 12893 27694
rect 12893 27642 12899 27694
rect 12781 27575 12787 27627
rect 12787 27575 12833 27627
rect 12847 27575 12893 27627
rect 12893 27575 12899 27627
rect 12781 27508 12787 27560
rect 12787 27508 12833 27560
rect 12847 27508 12893 27560
rect 12893 27508 12899 27560
rect 12781 27441 12787 27493
rect 12787 27441 12833 27493
rect 12847 27441 12893 27493
rect 12893 27441 12899 27493
rect 12781 27380 12787 27426
rect 12787 27380 12833 27426
rect 12847 27380 12893 27426
rect 12893 27380 12899 27426
rect 12781 27374 12833 27380
rect 12847 27374 12899 27380
rect 12781 25857 12833 25891
rect 12781 25839 12787 25857
rect 12787 25839 12821 25857
rect 12821 25839 12833 25857
rect 12847 25857 12899 25891
rect 12847 25839 12859 25857
rect 12859 25839 12893 25857
rect 12893 25839 12899 25857
rect 12781 25823 12787 25825
rect 12787 25823 12821 25825
rect 12821 25823 12833 25825
rect 12781 25780 12833 25823
rect 12781 25773 12787 25780
rect 12787 25773 12821 25780
rect 12821 25773 12833 25780
rect 12847 25823 12859 25825
rect 12859 25823 12893 25825
rect 12893 25823 12899 25825
rect 12847 25780 12899 25823
rect 12847 25773 12859 25780
rect 12859 25773 12893 25780
rect 12893 25773 12899 25780
rect 12781 25746 12787 25759
rect 12787 25746 12821 25759
rect 12821 25746 12833 25759
rect 11945 25641 11997 25693
rect 12011 25641 12063 25693
rect 11945 25574 11997 25626
rect 12011 25574 12063 25626
rect 11945 25507 11997 25559
rect 12011 25507 12063 25559
rect 11945 25440 11997 25492
rect 12011 25440 12063 25492
rect 11945 25373 11997 25425
rect 12011 25373 12063 25425
rect 12781 25707 12833 25746
rect 12847 25746 12859 25759
rect 12859 25746 12893 25759
rect 12893 25746 12899 25759
rect 12847 25707 12899 25746
rect 12781 25641 12833 25693
rect 12847 25641 12899 25693
rect 12781 25574 12833 25626
rect 12847 25574 12899 25626
rect 12781 25507 12833 25559
rect 12847 25507 12899 25559
rect 12781 25440 12833 25492
rect 12847 25440 12899 25492
rect 12781 25373 12833 25425
rect 12847 25373 12899 25425
rect 13200 34714 13252 34720
rect 13200 34680 13205 34714
rect 13205 34680 13239 34714
rect 13239 34680 13252 34714
rect 13200 34668 13252 34680
rect 13270 34714 13322 34720
rect 13270 34680 13277 34714
rect 13277 34680 13311 34714
rect 13311 34680 13322 34714
rect 13270 34668 13322 34680
rect 13340 34668 13392 34720
rect 13410 34668 13462 34720
rect 13480 34668 13521 34720
rect 13521 34668 13532 34720
rect 13550 34668 13602 34720
rect 13200 34641 13252 34654
rect 13200 34607 13205 34641
rect 13205 34607 13239 34641
rect 13239 34607 13252 34641
rect 13200 34602 13252 34607
rect 13270 34641 13322 34654
rect 13270 34607 13277 34641
rect 13277 34607 13311 34641
rect 13311 34607 13322 34641
rect 13270 34602 13322 34607
rect 13340 34602 13392 34654
rect 13410 34602 13462 34654
rect 13480 34602 13521 34654
rect 13521 34602 13532 34654
rect 13550 34602 13602 34654
rect 13200 34568 13252 34588
rect 13200 34536 13205 34568
rect 13205 34536 13239 34568
rect 13239 34536 13252 34568
rect 13270 34568 13322 34588
rect 13270 34536 13277 34568
rect 13277 34536 13311 34568
rect 13311 34536 13322 34568
rect 13340 34536 13392 34588
rect 13410 34536 13462 34588
rect 13480 34536 13521 34588
rect 13521 34536 13532 34588
rect 13550 34536 13602 34588
rect 13200 34495 13252 34522
rect 13200 34470 13205 34495
rect 13205 34470 13239 34495
rect 13239 34470 13252 34495
rect 13270 34495 13322 34522
rect 13270 34470 13277 34495
rect 13277 34470 13311 34495
rect 13311 34470 13322 34495
rect 13340 34470 13392 34522
rect 13410 34470 13462 34522
rect 13480 34470 13521 34522
rect 13521 34470 13532 34522
rect 13550 34470 13602 34522
rect 13200 34422 13252 34456
rect 13270 34422 13322 34456
rect 13200 34404 13205 34422
rect 13205 34404 13252 34422
rect 13270 34404 13311 34422
rect 13311 34404 13322 34422
rect 13340 34404 13392 34456
rect 13410 34404 13462 34456
rect 13480 34404 13521 34456
rect 13521 34404 13532 34456
rect 13550 34404 13602 34456
rect 13200 34338 13205 34390
rect 13205 34338 13252 34390
rect 13270 34338 13311 34390
rect 13311 34338 13322 34390
rect 13340 34338 13392 34390
rect 13410 34338 13462 34390
rect 13480 34338 13521 34390
rect 13521 34338 13532 34390
rect 13550 34338 13602 34390
rect 13200 34271 13205 34323
rect 13205 34271 13252 34323
rect 13270 34271 13311 34323
rect 13311 34271 13322 34323
rect 13340 34271 13392 34323
rect 13410 34271 13462 34323
rect 13480 34271 13521 34323
rect 13521 34271 13532 34323
rect 13550 34271 13602 34323
rect 13200 34204 13205 34256
rect 13205 34204 13252 34256
rect 13270 34204 13311 34256
rect 13311 34204 13322 34256
rect 13340 34204 13392 34256
rect 13410 34204 13462 34256
rect 13480 34204 13521 34256
rect 13521 34204 13532 34256
rect 13550 34204 13602 34256
rect 13200 32714 13252 32720
rect 13200 32680 13205 32714
rect 13205 32680 13239 32714
rect 13239 32680 13252 32714
rect 13200 32668 13252 32680
rect 13270 32714 13322 32720
rect 13270 32680 13277 32714
rect 13277 32680 13311 32714
rect 13311 32680 13322 32714
rect 13270 32668 13322 32680
rect 13340 32668 13392 32720
rect 13410 32668 13462 32720
rect 13480 32668 13521 32720
rect 13521 32668 13532 32720
rect 13550 32668 13602 32720
rect 13200 32641 13252 32654
rect 13200 32607 13205 32641
rect 13205 32607 13239 32641
rect 13239 32607 13252 32641
rect 13200 32602 13252 32607
rect 13270 32641 13322 32654
rect 13270 32607 13277 32641
rect 13277 32607 13311 32641
rect 13311 32607 13322 32641
rect 13270 32602 13322 32607
rect 13340 32602 13392 32654
rect 13410 32602 13462 32654
rect 13480 32602 13521 32654
rect 13521 32602 13532 32654
rect 13550 32602 13602 32654
rect 13200 32568 13252 32588
rect 13200 32536 13205 32568
rect 13205 32536 13239 32568
rect 13239 32536 13252 32568
rect 13270 32568 13322 32588
rect 13270 32536 13277 32568
rect 13277 32536 13311 32568
rect 13311 32536 13322 32568
rect 13340 32536 13392 32588
rect 13410 32536 13462 32588
rect 13480 32536 13521 32588
rect 13521 32536 13532 32588
rect 13550 32536 13602 32588
rect 13200 32495 13252 32522
rect 13200 32470 13205 32495
rect 13205 32470 13239 32495
rect 13239 32470 13252 32495
rect 13270 32495 13322 32522
rect 13270 32470 13277 32495
rect 13277 32470 13311 32495
rect 13311 32470 13322 32495
rect 13340 32470 13392 32522
rect 13410 32470 13462 32522
rect 13480 32470 13521 32522
rect 13521 32470 13532 32522
rect 13550 32470 13602 32522
rect 13200 32422 13252 32456
rect 13270 32422 13322 32456
rect 13200 32404 13205 32422
rect 13205 32404 13252 32422
rect 13270 32404 13311 32422
rect 13311 32404 13322 32422
rect 13340 32404 13392 32456
rect 13410 32404 13462 32456
rect 13480 32404 13521 32456
rect 13521 32404 13532 32456
rect 13550 32404 13602 32456
rect 13200 32338 13205 32390
rect 13205 32338 13252 32390
rect 13270 32338 13311 32390
rect 13311 32338 13322 32390
rect 13340 32338 13392 32390
rect 13410 32338 13462 32390
rect 13480 32338 13521 32390
rect 13521 32338 13532 32390
rect 13550 32338 13602 32390
rect 13200 32271 13205 32323
rect 13205 32271 13252 32323
rect 13270 32271 13311 32323
rect 13311 32271 13322 32323
rect 13340 32271 13392 32323
rect 13410 32271 13462 32323
rect 13480 32271 13521 32323
rect 13521 32271 13532 32323
rect 13550 32271 13602 32323
rect 13200 32204 13205 32256
rect 13205 32204 13252 32256
rect 13270 32204 13311 32256
rect 13311 32204 13322 32256
rect 13340 32204 13392 32256
rect 13410 32204 13462 32256
rect 13480 32204 13521 32256
rect 13521 32204 13532 32256
rect 13550 32204 13602 32256
rect 13200 30714 13252 30720
rect 13200 30680 13205 30714
rect 13205 30680 13239 30714
rect 13239 30680 13252 30714
rect 13200 30668 13252 30680
rect 13270 30714 13322 30720
rect 13270 30680 13277 30714
rect 13277 30680 13311 30714
rect 13311 30680 13322 30714
rect 13270 30668 13322 30680
rect 13340 30668 13392 30720
rect 13410 30668 13462 30720
rect 13480 30668 13521 30720
rect 13521 30668 13532 30720
rect 13550 30668 13602 30720
rect 13200 30641 13252 30654
rect 13200 30607 13205 30641
rect 13205 30607 13239 30641
rect 13239 30607 13252 30641
rect 13200 30602 13252 30607
rect 13270 30641 13322 30654
rect 13270 30607 13277 30641
rect 13277 30607 13311 30641
rect 13311 30607 13322 30641
rect 13270 30602 13322 30607
rect 13340 30602 13392 30654
rect 13410 30602 13462 30654
rect 13480 30602 13521 30654
rect 13521 30602 13532 30654
rect 13550 30602 13602 30654
rect 13200 30568 13252 30588
rect 13200 30536 13205 30568
rect 13205 30536 13239 30568
rect 13239 30536 13252 30568
rect 13270 30568 13322 30588
rect 13270 30536 13277 30568
rect 13277 30536 13311 30568
rect 13311 30536 13322 30568
rect 13340 30536 13392 30588
rect 13410 30536 13462 30588
rect 13480 30536 13521 30588
rect 13521 30536 13532 30588
rect 13550 30536 13602 30588
rect 13200 30495 13252 30522
rect 13200 30470 13205 30495
rect 13205 30470 13239 30495
rect 13239 30470 13252 30495
rect 13270 30495 13322 30522
rect 13270 30470 13277 30495
rect 13277 30470 13311 30495
rect 13311 30470 13322 30495
rect 13340 30470 13392 30522
rect 13410 30470 13462 30522
rect 13480 30470 13521 30522
rect 13521 30470 13532 30522
rect 13550 30470 13602 30522
rect 13200 30422 13252 30456
rect 13270 30422 13322 30456
rect 13200 30404 13205 30422
rect 13205 30404 13252 30422
rect 13270 30404 13311 30422
rect 13311 30404 13322 30422
rect 13340 30404 13392 30456
rect 13410 30404 13462 30456
rect 13480 30404 13521 30456
rect 13521 30404 13532 30456
rect 13550 30404 13602 30456
rect 13200 30338 13205 30390
rect 13205 30338 13252 30390
rect 13270 30338 13311 30390
rect 13311 30338 13322 30390
rect 13340 30338 13392 30390
rect 13410 30338 13462 30390
rect 13480 30338 13521 30390
rect 13521 30338 13532 30390
rect 13550 30338 13602 30390
rect 13200 30271 13205 30323
rect 13205 30271 13252 30323
rect 13270 30271 13311 30323
rect 13311 30271 13322 30323
rect 13340 30271 13392 30323
rect 13410 30271 13462 30323
rect 13480 30271 13521 30323
rect 13521 30271 13532 30323
rect 13550 30271 13602 30323
rect 13200 30204 13205 30256
rect 13205 30204 13252 30256
rect 13270 30204 13311 30256
rect 13311 30204 13322 30256
rect 13340 30204 13392 30256
rect 13410 30204 13462 30256
rect 13480 30204 13521 30256
rect 13521 30204 13532 30256
rect 13550 30204 13602 30256
rect 13200 28714 13252 28720
rect 13200 28680 13205 28714
rect 13205 28680 13239 28714
rect 13239 28680 13252 28714
rect 13200 28668 13252 28680
rect 13270 28714 13322 28720
rect 13270 28680 13277 28714
rect 13277 28680 13311 28714
rect 13311 28680 13322 28714
rect 13270 28668 13322 28680
rect 13340 28668 13392 28720
rect 13410 28668 13462 28720
rect 13480 28668 13521 28720
rect 13521 28668 13532 28720
rect 13550 28668 13602 28720
rect 13200 28641 13252 28654
rect 13200 28607 13205 28641
rect 13205 28607 13239 28641
rect 13239 28607 13252 28641
rect 13200 28602 13252 28607
rect 13270 28641 13322 28654
rect 13270 28607 13277 28641
rect 13277 28607 13311 28641
rect 13311 28607 13322 28641
rect 13270 28602 13322 28607
rect 13340 28602 13392 28654
rect 13410 28602 13462 28654
rect 13480 28602 13521 28654
rect 13521 28602 13532 28654
rect 13550 28602 13602 28654
rect 13200 28568 13252 28588
rect 13200 28536 13205 28568
rect 13205 28536 13239 28568
rect 13239 28536 13252 28568
rect 13270 28568 13322 28588
rect 13270 28536 13277 28568
rect 13277 28536 13311 28568
rect 13311 28536 13322 28568
rect 13340 28536 13392 28588
rect 13410 28536 13462 28588
rect 13480 28536 13521 28588
rect 13521 28536 13532 28588
rect 13550 28536 13602 28588
rect 13200 28495 13252 28522
rect 13200 28470 13205 28495
rect 13205 28470 13239 28495
rect 13239 28470 13252 28495
rect 13270 28495 13322 28522
rect 13270 28470 13277 28495
rect 13277 28470 13311 28495
rect 13311 28470 13322 28495
rect 13340 28470 13392 28522
rect 13410 28470 13462 28522
rect 13480 28470 13521 28522
rect 13521 28470 13532 28522
rect 13550 28470 13602 28522
rect 13200 28422 13252 28456
rect 13270 28422 13322 28456
rect 13200 28404 13205 28422
rect 13205 28404 13252 28422
rect 13270 28404 13311 28422
rect 13311 28404 13322 28422
rect 13340 28404 13392 28456
rect 13410 28404 13462 28456
rect 13480 28404 13521 28456
rect 13521 28404 13532 28456
rect 13550 28404 13602 28456
rect 13200 28338 13205 28390
rect 13205 28338 13252 28390
rect 13270 28338 13311 28390
rect 13311 28338 13322 28390
rect 13340 28338 13392 28390
rect 13410 28338 13462 28390
rect 13480 28338 13521 28390
rect 13521 28338 13532 28390
rect 13550 28338 13602 28390
rect 13200 28271 13205 28323
rect 13205 28271 13252 28323
rect 13270 28271 13311 28323
rect 13311 28271 13322 28323
rect 13340 28271 13392 28323
rect 13410 28271 13462 28323
rect 13480 28271 13521 28323
rect 13521 28271 13532 28323
rect 13550 28271 13602 28323
rect 13200 28204 13205 28256
rect 13205 28204 13252 28256
rect 13270 28204 13311 28256
rect 13311 28204 13322 28256
rect 13340 28204 13392 28256
rect 13410 28204 13462 28256
rect 13480 28204 13521 28256
rect 13521 28204 13532 28256
rect 13550 28204 13602 28256
rect 13200 26717 13205 26720
rect 13205 26717 13239 26720
rect 13239 26717 13252 26720
rect 13200 26676 13252 26717
rect 13200 26668 13205 26676
rect 13205 26668 13239 26676
rect 13239 26668 13252 26676
rect 13270 26717 13277 26720
rect 13277 26717 13311 26720
rect 13311 26717 13322 26720
rect 13270 26676 13322 26717
rect 13270 26668 13277 26676
rect 13277 26668 13311 26676
rect 13311 26668 13322 26676
rect 13340 26668 13392 26720
rect 13410 26668 13462 26720
rect 13480 26668 13521 26720
rect 13521 26668 13532 26720
rect 13550 26668 13602 26720
rect 13200 26642 13205 26654
rect 13205 26642 13239 26654
rect 13239 26642 13252 26654
rect 13200 26602 13252 26642
rect 13270 26642 13277 26654
rect 13277 26642 13311 26654
rect 13311 26642 13322 26654
rect 13270 26602 13322 26642
rect 13340 26602 13392 26654
rect 13410 26602 13462 26654
rect 13480 26602 13521 26654
rect 13521 26602 13532 26654
rect 13550 26602 13602 26654
rect 13200 26567 13205 26588
rect 13205 26567 13239 26588
rect 13239 26567 13252 26588
rect 13200 26536 13252 26567
rect 13270 26567 13277 26588
rect 13277 26567 13311 26588
rect 13311 26567 13322 26588
rect 13270 26536 13322 26567
rect 13340 26536 13392 26588
rect 13410 26536 13462 26588
rect 13480 26536 13521 26588
rect 13521 26536 13532 26588
rect 13550 26536 13602 26588
rect 13200 26492 13205 26522
rect 13205 26492 13239 26522
rect 13239 26492 13252 26522
rect 13200 26470 13252 26492
rect 13270 26492 13277 26522
rect 13277 26492 13311 26522
rect 13311 26492 13322 26522
rect 13270 26470 13322 26492
rect 13340 26470 13392 26522
rect 13410 26470 13462 26522
rect 13480 26470 13521 26522
rect 13521 26470 13532 26522
rect 13550 26470 13602 26522
rect 13200 26451 13252 26456
rect 13200 26417 13205 26451
rect 13205 26417 13239 26451
rect 13239 26417 13252 26451
rect 13200 26404 13252 26417
rect 13270 26451 13322 26456
rect 13270 26417 13277 26451
rect 13277 26417 13311 26451
rect 13311 26417 13322 26451
rect 13270 26404 13322 26417
rect 13340 26404 13392 26456
rect 13410 26404 13462 26456
rect 13480 26404 13521 26456
rect 13521 26404 13532 26456
rect 13550 26404 13602 26456
rect 13200 26376 13252 26389
rect 13200 26342 13205 26376
rect 13205 26342 13239 26376
rect 13239 26342 13252 26376
rect 13200 26337 13252 26342
rect 13270 26376 13322 26389
rect 13270 26342 13277 26376
rect 13277 26342 13311 26376
rect 13311 26342 13322 26376
rect 13270 26337 13322 26342
rect 13340 26337 13392 26389
rect 13410 26337 13462 26389
rect 13480 26337 13521 26389
rect 13521 26337 13532 26389
rect 13550 26337 13602 26389
rect 13200 26301 13252 26322
rect 13200 26270 13205 26301
rect 13205 26270 13239 26301
rect 13239 26270 13252 26301
rect 13270 26301 13322 26322
rect 13270 26270 13277 26301
rect 13277 26270 13311 26301
rect 13311 26270 13322 26301
rect 13340 26270 13392 26322
rect 13410 26270 13462 26322
rect 13480 26270 13521 26322
rect 13521 26270 13532 26322
rect 13550 26270 13602 26322
rect 13200 26226 13252 26255
rect 13200 26203 13205 26226
rect 13205 26203 13239 26226
rect 13239 26203 13252 26226
rect 13270 26226 13322 26255
rect 13270 26203 13277 26226
rect 13277 26203 13311 26226
rect 13311 26203 13322 26226
rect 13340 26203 13392 26255
rect 13410 26203 13462 26255
rect 13480 26203 13521 26255
rect 13521 26203 13532 26255
rect 13550 26203 13602 26255
rect 5075 23697 5127 23703
rect 5075 23663 5081 23697
rect 5081 23663 5115 23697
rect 5115 23663 5127 23697
rect 5075 23651 5127 23663
rect 5151 23697 5203 23703
rect 5151 23663 5154 23697
rect 5154 23663 5188 23697
rect 5188 23663 5203 23697
rect 5151 23651 5203 23663
rect 5226 23697 5278 23703
rect 5301 23697 5353 23703
rect 5376 23697 5428 23703
rect 5451 23697 5503 23703
rect 5226 23663 5227 23697
rect 5227 23663 5261 23697
rect 5261 23663 5278 23697
rect 5301 23663 5334 23697
rect 5334 23663 5353 23697
rect 5376 23663 5407 23697
rect 5407 23663 5428 23697
rect 5451 23663 5480 23697
rect 5480 23663 5503 23697
rect 5226 23651 5278 23663
rect 5301 23651 5353 23663
rect 5376 23651 5428 23663
rect 5451 23651 5503 23663
rect 5075 23575 5127 23627
rect 5151 23575 5203 23627
rect 5226 23575 5278 23627
rect 5301 23575 5353 23627
rect 5376 23575 5428 23627
rect 5451 23575 5503 23627
rect 5075 23499 5127 23551
rect 5151 23499 5203 23551
rect 5226 23499 5278 23551
rect 5301 23499 5353 23551
rect 5376 23499 5428 23551
rect 5451 23499 5503 23551
rect 5075 23462 5127 23475
rect 5075 23428 5081 23462
rect 5081 23428 5115 23462
rect 5115 23428 5127 23462
rect 5075 23423 5127 23428
rect 5151 23462 5203 23475
rect 5151 23428 5154 23462
rect 5154 23428 5188 23462
rect 5188 23428 5203 23462
rect 5151 23423 5203 23428
rect 5226 23462 5278 23475
rect 5301 23462 5353 23475
rect 5376 23462 5428 23475
rect 5451 23462 5503 23475
rect 5226 23428 5227 23462
rect 5227 23428 5261 23462
rect 5261 23428 5278 23462
rect 5301 23428 5334 23462
rect 5334 23428 5353 23462
rect 5376 23428 5407 23462
rect 5407 23428 5428 23462
rect 5451 23428 5480 23462
rect 5480 23428 5503 23462
rect 5226 23423 5278 23428
rect 5301 23423 5353 23428
rect 5376 23423 5428 23428
rect 5451 23423 5503 23428
rect 5073 21763 5125 21775
rect 5073 21729 5079 21763
rect 5079 21729 5113 21763
rect 5113 21729 5125 21763
rect 5073 21723 5125 21729
rect 5140 21763 5192 21775
rect 5140 21729 5152 21763
rect 5152 21729 5186 21763
rect 5186 21729 5192 21763
rect 5140 21723 5192 21729
rect 5206 21763 5258 21775
rect 5272 21763 5324 21775
rect 5206 21729 5225 21763
rect 5225 21729 5258 21763
rect 5272 21729 5298 21763
rect 5298 21729 5324 21763
rect 5206 21723 5258 21729
rect 5272 21723 5324 21729
rect 4917 19742 4969 19754
rect 4917 19708 4923 19742
rect 4923 19708 4957 19742
rect 4957 19708 4969 19742
rect 4917 19702 4969 19708
rect 4981 19742 5033 19754
rect 4981 19708 4996 19742
rect 4996 19708 5030 19742
rect 5030 19708 5033 19742
rect 4981 19702 5033 19708
rect 13200 19654 13252 19706
rect 13270 19654 13322 19706
rect 13340 19654 13392 19706
rect 13410 19654 13462 19706
rect 13480 19654 13490 19706
rect 13490 19654 13532 19706
rect 13550 19654 13596 19706
rect 13596 19654 13602 19706
rect 4481 16643 4533 16657
rect 4481 16609 4486 16643
rect 4486 16609 4520 16643
rect 4520 16609 4533 16643
rect 4481 16605 4533 16609
rect 4545 16605 4597 16657
rect 4609 16643 4661 16657
rect 4609 16609 4622 16643
rect 4622 16609 4656 16643
rect 4656 16609 4661 16643
rect 4609 16605 4661 16609
rect 13200 19590 13252 19642
rect 13270 19590 13322 19642
rect 13340 19590 13392 19642
rect 13410 19590 13462 19642
rect 13480 19590 13490 19642
rect 13490 19590 13532 19642
rect 13550 19590 13596 19642
rect 13596 19590 13602 19642
rect 13200 19526 13252 19578
rect 13270 19526 13322 19578
rect 13340 19574 13392 19578
rect 13340 19540 13342 19574
rect 13342 19540 13376 19574
rect 13376 19540 13392 19574
rect 13340 19526 13392 19540
rect 13410 19526 13462 19578
rect 13480 19526 13490 19578
rect 13490 19526 13532 19578
rect 13550 19526 13596 19578
rect 13596 19526 13602 19578
rect 13200 19462 13252 19514
rect 13270 19462 13322 19514
rect 13340 19498 13392 19514
rect 13340 19464 13342 19498
rect 13342 19464 13376 19498
rect 13376 19464 13392 19498
rect 13340 19462 13392 19464
rect 13410 19462 13462 19514
rect 13480 19462 13490 19514
rect 13490 19462 13532 19514
rect 13550 19462 13596 19514
rect 13596 19462 13602 19514
rect 13200 19398 13252 19450
rect 13270 19398 13322 19450
rect 13340 19422 13392 19450
rect 13340 19398 13342 19422
rect 13342 19398 13376 19422
rect 13376 19398 13392 19422
rect 13410 19398 13462 19450
rect 13480 19398 13490 19450
rect 13490 19398 13532 19450
rect 13550 19398 13596 19450
rect 13596 19398 13602 19450
rect 13200 19334 13252 19386
rect 13270 19334 13322 19386
rect 13340 19346 13392 19386
rect 13340 19334 13342 19346
rect 13342 19334 13376 19346
rect 13376 19334 13392 19346
rect 13410 19334 13462 19386
rect 13480 19334 13490 19386
rect 13490 19334 13532 19386
rect 13550 19334 13596 19386
rect 13596 19334 13602 19386
rect 13200 19270 13252 19322
rect 13270 19270 13322 19322
rect 13340 19312 13342 19322
rect 13342 19312 13376 19322
rect 13376 19312 13392 19322
rect 13340 19270 13392 19312
rect 13410 19270 13462 19322
rect 13480 19270 13490 19322
rect 13490 19270 13532 19322
rect 13550 19270 13596 19322
rect 13596 19270 13602 19322
rect 13200 19206 13252 19258
rect 13270 19206 13322 19258
rect 13340 19236 13342 19258
rect 13342 19236 13376 19258
rect 13376 19236 13392 19258
rect 13340 19206 13392 19236
rect 13410 19206 13462 19258
rect 13480 19206 13490 19258
rect 13490 19206 13532 19258
rect 13550 19206 13596 19258
rect 13596 19206 13602 19258
rect 13200 19142 13252 19194
rect 13270 19142 13322 19194
rect 13340 19160 13342 19194
rect 13342 19160 13376 19194
rect 13376 19160 13392 19194
rect 13340 19142 13392 19160
rect 13410 19142 13462 19194
rect 13480 19142 13490 19194
rect 13490 19142 13532 19194
rect 13550 19142 13596 19194
rect 13596 19142 13602 19194
rect 13200 19078 13252 19130
rect 13270 19078 13322 19130
rect 13340 19118 13392 19130
rect 13340 19084 13342 19118
rect 13342 19084 13376 19118
rect 13376 19084 13392 19118
rect 13340 19078 13392 19084
rect 13410 19078 13462 19130
rect 13480 19078 13490 19130
rect 13490 19078 13532 19130
rect 13550 19078 13596 19130
rect 13596 19078 13602 19130
rect 13200 19014 13252 19066
rect 13270 19014 13322 19066
rect 13340 19042 13392 19066
rect 13340 19014 13342 19042
rect 13342 19014 13376 19042
rect 13376 19014 13392 19042
rect 13410 19014 13462 19066
rect 13480 19014 13490 19066
rect 13490 19014 13532 19066
rect 13550 19014 13596 19066
rect 13596 19014 13602 19066
rect 13200 18950 13252 19002
rect 13270 18950 13322 19002
rect 13340 18966 13392 19002
rect 13340 18950 13342 18966
rect 13342 18950 13376 18966
rect 13376 18950 13392 18966
rect 13410 18950 13462 19002
rect 13480 18950 13490 19002
rect 13490 18950 13532 19002
rect 13550 18950 13596 19002
rect 13596 18950 13602 19002
rect 13200 18886 13252 18938
rect 13270 18886 13322 18938
rect 13340 18932 13342 18938
rect 13342 18932 13376 18938
rect 13376 18932 13392 18938
rect 13340 18890 13392 18932
rect 13340 18886 13342 18890
rect 13342 18886 13376 18890
rect 13376 18886 13392 18890
rect 13410 18886 13462 18938
rect 13480 18886 13490 18938
rect 13490 18886 13532 18938
rect 13550 18886 13596 18938
rect 13596 18886 13602 18938
rect 13200 18822 13252 18874
rect 13270 18822 13322 18874
rect 13340 18856 13342 18874
rect 13342 18856 13376 18874
rect 13376 18856 13392 18874
rect 13340 18822 13392 18856
rect 13410 18822 13462 18874
rect 13480 18822 13490 18874
rect 13490 18822 13532 18874
rect 13550 18822 13596 18874
rect 13596 18822 13602 18874
rect 13200 18758 13252 18810
rect 13270 18758 13322 18810
rect 13340 18781 13342 18810
rect 13342 18781 13376 18810
rect 13376 18781 13392 18810
rect 13340 18758 13392 18781
rect 13410 18758 13462 18810
rect 13480 18758 13490 18810
rect 13490 18758 13532 18810
rect 13550 18758 13596 18810
rect 13596 18758 13602 18810
rect 13200 18694 13252 18746
rect 13270 18694 13322 18746
rect 13340 18740 13392 18746
rect 13340 18706 13342 18740
rect 13342 18706 13376 18740
rect 13376 18706 13392 18740
rect 13340 18694 13392 18706
rect 13410 18694 13462 18746
rect 13480 18694 13490 18746
rect 13490 18694 13532 18746
rect 13550 18694 13596 18746
rect 13596 18694 13602 18746
rect 13200 18630 13252 18682
rect 13270 18630 13322 18682
rect 13340 18665 13392 18682
rect 13340 18631 13342 18665
rect 13342 18631 13376 18665
rect 13376 18631 13392 18665
rect 13340 18630 13392 18631
rect 13410 18630 13462 18682
rect 13480 18630 13490 18682
rect 13490 18630 13532 18682
rect 13550 18630 13596 18682
rect 13596 18630 13602 18682
rect 13200 18566 13252 18618
rect 13270 18566 13322 18618
rect 13340 18590 13392 18618
rect 13340 18566 13342 18590
rect 13342 18566 13376 18590
rect 13376 18566 13392 18590
rect 13410 18566 13462 18618
rect 13480 18566 13490 18618
rect 13490 18566 13532 18618
rect 13550 18566 13596 18618
rect 13596 18566 13602 18618
rect 13200 18502 13252 18554
rect 13270 18502 13322 18554
rect 13340 18515 13392 18554
rect 13340 18502 13342 18515
rect 13342 18502 13376 18515
rect 13376 18502 13392 18515
rect 13410 18502 13462 18554
rect 13480 18502 13490 18554
rect 13490 18502 13532 18554
rect 13550 18502 13596 18554
rect 13596 18502 13602 18554
rect 13200 18438 13252 18490
rect 13270 18438 13322 18490
rect 13340 18481 13342 18490
rect 13342 18481 13376 18490
rect 13376 18481 13392 18490
rect 13340 18440 13392 18481
rect 13340 18438 13342 18440
rect 13342 18438 13376 18440
rect 13376 18438 13392 18440
rect 13410 18438 13462 18490
rect 13480 18438 13490 18490
rect 13490 18438 13532 18490
rect 13550 18438 13596 18490
rect 13596 18438 13602 18490
rect 13200 18374 13252 18426
rect 13270 18374 13322 18426
rect 13340 18406 13342 18426
rect 13342 18406 13376 18426
rect 13376 18406 13392 18426
rect 13340 18374 13392 18406
rect 13410 18374 13462 18426
rect 13480 18374 13490 18426
rect 13490 18374 13532 18426
rect 13550 18374 13596 18426
rect 13596 18374 13602 18426
rect 13200 18310 13252 18362
rect 13270 18310 13322 18362
rect 13340 18331 13342 18362
rect 13342 18331 13376 18362
rect 13376 18331 13392 18362
rect 13340 18310 13392 18331
rect 13410 18310 13462 18362
rect 13480 18310 13490 18362
rect 13490 18310 13532 18362
rect 13550 18310 13596 18362
rect 13596 18310 13602 18362
rect 13200 18246 13252 18298
rect 13270 18246 13322 18298
rect 13340 18290 13392 18298
rect 13340 18256 13342 18290
rect 13342 18256 13376 18290
rect 13376 18256 13392 18290
rect 13340 18246 13392 18256
rect 13410 18246 13462 18298
rect 13480 18246 13490 18298
rect 13490 18246 13532 18298
rect 13550 18246 13596 18298
rect 13596 18246 13602 18298
rect 13200 18182 13252 18234
rect 13270 18182 13322 18234
rect 13340 18182 13392 18234
rect 13410 18182 13462 18234
rect 13480 18182 13490 18234
rect 13490 18182 13532 18234
rect 13550 18182 13596 18234
rect 13596 18182 13602 18234
rect 13200 18118 13252 18170
rect 13270 18118 13322 18170
rect 13340 18118 13392 18170
rect 13410 18118 13462 18170
rect 13480 18118 13490 18170
rect 13490 18118 13532 18170
rect 13550 18118 13596 18170
rect 13596 18118 13602 18170
rect 4917 18043 4969 18055
rect 4917 18009 4923 18043
rect 4923 18009 4957 18043
rect 4957 18009 4969 18043
rect 4917 18003 4969 18009
rect 4981 18043 5033 18055
rect 13200 18054 13252 18106
rect 13270 18054 13322 18106
rect 13340 18054 13392 18106
rect 13410 18054 13462 18106
rect 13480 18054 13490 18106
rect 13490 18054 13532 18106
rect 13550 18054 13596 18106
rect 13596 18054 13602 18106
rect 4981 18009 4996 18043
rect 4996 18009 5030 18043
rect 5030 18009 5033 18043
rect 4981 18003 5033 18009
rect 13200 17990 13252 18042
rect 13270 17990 13322 18042
rect 13340 17990 13392 18042
rect 13410 17990 13462 18042
rect 13480 17990 13490 18042
rect 13490 17990 13532 18042
rect 13550 17990 13596 18042
rect 13596 17990 13602 18042
rect 13200 17926 13252 17978
rect 13270 17926 13322 17978
rect 13340 17926 13392 17978
rect 13410 17926 13462 17978
rect 13480 17926 13490 17978
rect 13490 17926 13532 17978
rect 13550 17926 13596 17978
rect 13596 17926 13602 17978
rect 13200 17862 13252 17914
rect 13270 17862 13322 17914
rect 13340 17875 13392 17914
rect 13340 17862 13342 17875
rect 13342 17862 13376 17875
rect 13376 17862 13392 17875
rect 13410 17862 13462 17914
rect 13480 17862 13490 17914
rect 13490 17862 13532 17914
rect 13550 17862 13596 17914
rect 13596 17862 13602 17914
rect 4731 16776 4737 16809
rect 4737 16776 4771 16809
rect 4771 16776 4783 16809
rect 4731 16757 4783 16776
rect 4797 16776 4809 16809
rect 4809 16776 4843 16809
rect 4843 16776 4849 16809
rect 4797 16757 4849 16776
rect 4731 16703 4737 16706
rect 4737 16703 4771 16706
rect 4771 16703 4783 16706
rect 4731 16664 4783 16703
rect 4731 16654 4737 16664
rect 4737 16654 4771 16664
rect 4771 16654 4783 16664
rect 4797 16703 4809 16706
rect 4809 16703 4843 16706
rect 4843 16703 4849 16706
rect 4797 16664 4849 16703
rect 4797 16654 4809 16664
rect 4809 16654 4843 16664
rect 4843 16654 4849 16664
rect 4731 16591 4783 16603
rect 4731 16557 4737 16591
rect 4737 16557 4771 16591
rect 4771 16557 4783 16591
rect 4731 16551 4783 16557
rect 4797 16591 4849 16603
rect 4797 16557 4809 16591
rect 4809 16557 4843 16591
rect 4843 16557 4849 16591
rect 13200 17798 13252 17850
rect 13270 17798 13322 17850
rect 13340 17841 13342 17850
rect 13342 17841 13376 17850
rect 13376 17841 13392 17850
rect 13340 17800 13392 17841
rect 13340 17798 13342 17800
rect 13342 17798 13376 17800
rect 13376 17798 13392 17800
rect 13410 17798 13462 17850
rect 13480 17798 13490 17850
rect 13490 17798 13532 17850
rect 13550 17798 13596 17850
rect 13596 17798 13602 17850
rect 13200 17734 13252 17786
rect 13270 17734 13322 17786
rect 13340 17766 13342 17786
rect 13342 17766 13376 17786
rect 13376 17766 13392 17786
rect 13340 17734 13392 17766
rect 13410 17734 13462 17786
rect 13480 17734 13490 17786
rect 13490 17734 13532 17786
rect 13550 17734 13596 17786
rect 13596 17734 13602 17786
rect 13200 17670 13252 17722
rect 13270 17670 13322 17722
rect 13340 17691 13342 17722
rect 13342 17691 13376 17722
rect 13376 17691 13392 17722
rect 13340 17670 13392 17691
rect 13410 17670 13462 17722
rect 13480 17670 13490 17722
rect 13490 17670 13532 17722
rect 13550 17670 13596 17722
rect 13596 17670 13602 17722
rect 13200 17606 13252 17658
rect 13270 17606 13322 17658
rect 13340 17650 13392 17658
rect 13340 17616 13342 17650
rect 13342 17616 13376 17650
rect 13376 17616 13392 17650
rect 13340 17606 13392 17616
rect 13410 17606 13462 17658
rect 13480 17606 13490 17658
rect 13490 17606 13532 17658
rect 13550 17606 13596 17658
rect 13596 17606 13602 17658
rect 13200 17542 13252 17594
rect 13270 17542 13322 17594
rect 13340 17575 13392 17594
rect 13340 17542 13342 17575
rect 13342 17542 13376 17575
rect 13376 17542 13392 17575
rect 13410 17542 13462 17594
rect 13480 17542 13490 17594
rect 13490 17542 13532 17594
rect 13550 17542 13596 17594
rect 13596 17542 13602 17594
rect 13200 17478 13252 17530
rect 13270 17478 13322 17530
rect 13340 17500 13392 17530
rect 13340 17478 13342 17500
rect 13342 17478 13376 17500
rect 13376 17478 13392 17500
rect 13410 17478 13462 17530
rect 13480 17478 13490 17530
rect 13490 17478 13532 17530
rect 13550 17478 13596 17530
rect 13596 17478 13602 17530
rect 13200 17414 13252 17466
rect 13270 17414 13322 17466
rect 13340 17425 13392 17466
rect 13340 17414 13342 17425
rect 13342 17414 13376 17425
rect 13376 17414 13392 17425
rect 13410 17414 13462 17466
rect 13480 17414 13490 17466
rect 13490 17414 13532 17466
rect 13550 17414 13596 17466
rect 13596 17414 13602 17466
rect 13200 17350 13252 17402
rect 13270 17350 13322 17402
rect 13340 17391 13342 17402
rect 13342 17391 13376 17402
rect 13376 17391 13392 17402
rect 13340 17350 13392 17391
rect 13410 17350 13462 17402
rect 13480 17350 13490 17402
rect 13490 17350 13532 17402
rect 13550 17350 13596 17402
rect 13596 17350 13602 17402
rect 13200 17286 13252 17338
rect 13270 17286 13322 17338
rect 13340 17316 13342 17338
rect 13342 17316 13376 17338
rect 13376 17316 13392 17338
rect 13340 17286 13392 17316
rect 13410 17286 13462 17338
rect 13480 17286 13490 17338
rect 13490 17286 13532 17338
rect 13550 17286 13596 17338
rect 13596 17286 13602 17338
rect 13200 17222 13252 17274
rect 13270 17222 13322 17274
rect 13340 17241 13342 17274
rect 13342 17241 13376 17274
rect 13376 17241 13392 17274
rect 13340 17222 13392 17241
rect 13410 17222 13462 17274
rect 13480 17222 13490 17274
rect 13490 17222 13532 17274
rect 13550 17222 13596 17274
rect 13596 17222 13602 17274
rect 13200 17158 13252 17210
rect 13270 17158 13322 17210
rect 13340 17199 13392 17210
rect 13340 17165 13342 17199
rect 13342 17165 13376 17199
rect 13376 17165 13392 17199
rect 13340 17158 13392 17165
rect 13410 17158 13462 17210
rect 13480 17158 13490 17210
rect 13490 17158 13532 17210
rect 13550 17158 13596 17210
rect 13596 17158 13602 17210
rect 13200 17094 13252 17146
rect 13270 17094 13322 17146
rect 13340 17123 13392 17146
rect 13340 17094 13342 17123
rect 13342 17094 13376 17123
rect 13376 17094 13392 17123
rect 13410 17094 13462 17146
rect 13480 17094 13490 17146
rect 13490 17094 13532 17146
rect 13550 17094 13596 17146
rect 13596 17094 13602 17146
rect 13200 17030 13252 17082
rect 13270 17030 13322 17082
rect 13340 17047 13392 17082
rect 13340 17030 13342 17047
rect 13342 17030 13376 17047
rect 13376 17030 13392 17047
rect 13410 17030 13462 17082
rect 13480 17030 13490 17082
rect 13490 17030 13532 17082
rect 13550 17030 13596 17082
rect 13596 17030 13602 17082
rect 13200 16966 13252 17018
rect 13270 16966 13322 17018
rect 13340 17013 13342 17018
rect 13342 17013 13376 17018
rect 13376 17013 13392 17018
rect 13340 16971 13392 17013
rect 13340 16966 13342 16971
rect 13342 16966 13376 16971
rect 13376 16966 13392 16971
rect 13410 16966 13462 17018
rect 13480 16966 13490 17018
rect 13490 16966 13532 17018
rect 13550 16966 13596 17018
rect 13596 16966 13602 17018
rect 13200 16902 13252 16954
rect 13270 16902 13322 16954
rect 13340 16937 13342 16954
rect 13342 16937 13376 16954
rect 13376 16937 13392 16954
rect 13340 16902 13392 16937
rect 13410 16902 13462 16954
rect 13480 16902 13490 16954
rect 13490 16902 13532 16954
rect 13550 16902 13596 16954
rect 13596 16902 13602 16954
rect 13200 16838 13252 16890
rect 13270 16838 13322 16890
rect 13340 16861 13342 16890
rect 13342 16861 13376 16890
rect 13376 16861 13392 16890
rect 13340 16838 13392 16861
rect 13410 16838 13462 16890
rect 13480 16838 13490 16890
rect 13490 16838 13532 16890
rect 13550 16838 13596 16890
rect 13596 16838 13602 16890
rect 13200 16774 13252 16826
rect 13270 16774 13322 16826
rect 13340 16819 13392 16826
rect 13340 16785 13342 16819
rect 13342 16785 13376 16819
rect 13376 16785 13392 16819
rect 13340 16774 13392 16785
rect 13410 16774 13462 16826
rect 13480 16774 13490 16826
rect 13490 16774 13532 16826
rect 13550 16774 13596 16826
rect 13596 16774 13602 16826
rect 13200 16710 13252 16762
rect 13270 16710 13322 16762
rect 13340 16743 13392 16762
rect 13340 16710 13342 16743
rect 13342 16710 13376 16743
rect 13376 16710 13392 16743
rect 13410 16710 13462 16762
rect 13480 16710 13490 16762
rect 13490 16710 13532 16762
rect 13550 16710 13596 16762
rect 13596 16710 13602 16762
rect 13200 16646 13252 16698
rect 13270 16646 13322 16698
rect 13340 16667 13392 16698
rect 13340 16646 13342 16667
rect 13342 16646 13376 16667
rect 13376 16646 13392 16667
rect 13410 16646 13462 16698
rect 13480 16646 13490 16698
rect 13490 16646 13532 16698
rect 13550 16646 13596 16698
rect 13596 16646 13602 16698
rect 13200 16582 13252 16634
rect 13270 16582 13322 16634
rect 13340 16633 13342 16634
rect 13342 16633 13376 16634
rect 13376 16633 13392 16634
rect 13340 16591 13392 16633
rect 13340 16582 13342 16591
rect 13342 16582 13376 16591
rect 13376 16582 13392 16591
rect 13410 16582 13462 16634
rect 13480 16582 13490 16634
rect 13490 16582 13532 16634
rect 13550 16582 13596 16634
rect 13596 16582 13602 16634
rect 4797 16551 4849 16557
rect 4481 16535 4486 16545
rect 4486 16535 4520 16545
rect 4520 16535 4533 16545
rect 4481 16495 4533 16535
rect 4481 16493 4486 16495
rect 4486 16493 4520 16495
rect 4520 16493 4533 16495
rect 4545 16493 4597 16545
rect 4609 16535 4622 16545
rect 4622 16535 4656 16545
rect 4656 16535 4661 16545
rect 4609 16495 4661 16535
rect 4609 16493 4622 16495
rect 4622 16493 4656 16495
rect 4656 16493 4661 16495
rect 4481 16421 4533 16433
rect 4481 16387 4486 16421
rect 4486 16387 4520 16421
rect 4520 16387 4533 16421
rect 4481 16381 4533 16387
rect 4545 16381 4597 16433
rect 4609 16421 4661 16433
rect 4609 16387 4622 16421
rect 4622 16387 4656 16421
rect 4656 16387 4661 16421
rect 4609 16381 4661 16387
rect 13200 16518 13252 16570
rect 13270 16518 13322 16570
rect 13340 16557 13342 16570
rect 13342 16557 13376 16570
rect 13376 16557 13392 16570
rect 13340 16518 13392 16557
rect 13410 16518 13462 16570
rect 13480 16518 13490 16570
rect 13490 16518 13532 16570
rect 13550 16518 13596 16570
rect 13596 16518 13602 16570
rect 13200 16454 13252 16506
rect 13270 16454 13322 16506
rect 13340 16454 13392 16506
rect 13410 16454 13462 16506
rect 13480 16454 13490 16506
rect 13490 16454 13532 16506
rect 13550 16454 13596 16506
rect 13596 16454 13602 16506
rect 13200 16390 13252 16442
rect 13270 16390 13322 16442
rect 13340 16390 13392 16442
rect 13410 16390 13462 16442
rect 13480 16390 13490 16442
rect 13490 16390 13532 16442
rect 13550 16390 13596 16442
rect 13596 16390 13602 16442
rect 13200 16326 13252 16378
rect 13270 16326 13322 16378
rect 13340 16326 13392 16378
rect 13410 16326 13462 16378
rect 13480 16326 13490 16378
rect 13490 16326 13532 16378
rect 13550 16326 13596 16378
rect 13596 16326 13602 16378
rect 4917 16243 4969 16271
rect 4917 16219 4923 16243
rect 4923 16219 4957 16243
rect 4957 16219 4969 16243
rect 4981 16243 5033 16271
rect 4981 16219 4996 16243
rect 4996 16219 5030 16243
rect 5030 16219 5033 16243
rect 13200 16262 13252 16314
rect 13270 16262 13322 16314
rect 13340 16262 13392 16314
rect 13410 16262 13462 16314
rect 13480 16262 13490 16314
rect 13490 16262 13532 16314
rect 13550 16262 13596 16314
rect 13596 16262 13602 16314
rect 13200 16198 13252 16250
rect 13270 16198 13322 16250
rect 13340 16198 13392 16250
rect 13410 16198 13462 16250
rect 13480 16198 13490 16250
rect 13490 16198 13532 16250
rect 13550 16198 13596 16250
rect 13596 16198 13602 16250
rect 13200 16134 13252 16186
rect 13270 16134 13322 16186
rect 13340 16134 13392 16186
rect 13410 16134 13462 16186
rect 13480 16134 13490 16186
rect 13490 16134 13532 16186
rect 13550 16134 13596 16186
rect 13596 16134 13602 16186
rect 13200 16070 13252 16122
rect 13270 16070 13322 16122
rect 13340 16107 13392 16122
rect 13340 16073 13342 16107
rect 13342 16073 13376 16107
rect 13376 16073 13392 16107
rect 13340 16070 13392 16073
rect 13410 16070 13462 16122
rect 13480 16070 13490 16122
rect 13490 16070 13532 16122
rect 13550 16070 13596 16122
rect 13596 16070 13602 16122
rect 4481 16014 4533 16066
rect 4545 16014 4597 16066
rect 4609 16014 4661 16066
rect 13200 16006 13252 16058
rect 13270 16006 13322 16058
rect 13340 16030 13392 16058
rect 13340 16006 13342 16030
rect 13342 16006 13376 16030
rect 13376 16006 13392 16030
rect 13410 16006 13462 16058
rect 13480 16006 13490 16058
rect 13490 16006 13532 16058
rect 13550 16006 13596 16058
rect 13596 16006 13602 16058
rect 13200 15942 13252 15994
rect 13270 15942 13322 15994
rect 13340 15953 13392 15994
rect 13340 15942 13342 15953
rect 13342 15942 13376 15953
rect 13376 15942 13392 15953
rect 13410 15942 13462 15994
rect 13480 15942 13490 15994
rect 13490 15942 13532 15994
rect 13550 15942 13596 15994
rect 13596 15942 13602 15994
rect 4481 15870 4533 15922
rect 4545 15870 4597 15922
rect 4609 15870 4661 15922
rect 13200 15878 13252 15930
rect 13270 15878 13322 15930
rect 13340 15919 13342 15930
rect 13342 15919 13376 15930
rect 13376 15919 13392 15930
rect 13340 15878 13392 15919
rect 13410 15878 13462 15930
rect 13480 15878 13490 15930
rect 13490 15878 13532 15930
rect 13550 15878 13596 15930
rect 13596 15878 13602 15930
rect 13200 15814 13252 15866
rect 13270 15814 13322 15866
rect 13340 15842 13342 15866
rect 13342 15842 13376 15866
rect 13376 15842 13392 15866
rect 13340 15814 13392 15842
rect 13410 15814 13462 15866
rect 13480 15814 13490 15866
rect 13490 15814 13532 15866
rect 13550 15814 13596 15866
rect 13596 15814 13602 15866
rect 4481 15726 4533 15778
rect 4545 15726 4597 15778
rect 4609 15726 4661 15778
rect 13200 15750 13252 15802
rect 13270 15750 13322 15802
rect 13340 15799 13392 15802
rect 13340 15765 13342 15799
rect 13342 15765 13376 15799
rect 13376 15765 13392 15799
rect 13340 15750 13392 15765
rect 13410 15750 13462 15802
rect 13480 15750 13490 15802
rect 13490 15750 13532 15802
rect 13550 15750 13596 15802
rect 13596 15750 13602 15802
rect 13200 15686 13252 15738
rect 13270 15686 13322 15738
rect 13340 15723 13392 15738
rect 13340 15689 13342 15723
rect 13342 15689 13376 15723
rect 13376 15689 13392 15723
rect 13340 15686 13392 15689
rect 13410 15686 13462 15738
rect 13480 15686 13490 15738
rect 13490 15686 13532 15738
rect 13550 15686 13596 15738
rect 13596 15686 13602 15738
rect 4481 15582 4533 15634
rect 4545 15582 4597 15634
rect 4609 15582 4661 15634
rect 13200 15622 13252 15674
rect 13270 15622 13322 15674
rect 13340 15647 13392 15674
rect 13340 15622 13342 15647
rect 13342 15622 13376 15647
rect 13376 15622 13392 15647
rect 13410 15622 13462 15674
rect 13480 15622 13490 15674
rect 13490 15622 13532 15674
rect 13550 15622 13596 15674
rect 13596 15622 13602 15674
rect 13200 15558 13252 15610
rect 13270 15558 13322 15610
rect 13340 15571 13392 15610
rect 13340 15558 13342 15571
rect 13342 15558 13376 15571
rect 13376 15558 13392 15571
rect 13410 15558 13462 15610
rect 13480 15558 13490 15610
rect 13490 15558 13532 15610
rect 13550 15558 13596 15610
rect 13596 15558 13602 15610
rect 13200 15494 13252 15546
rect 13270 15494 13322 15546
rect 13340 15537 13342 15546
rect 13342 15537 13376 15546
rect 13376 15537 13392 15546
rect 13340 15495 13392 15537
rect 13340 15494 13342 15495
rect 13342 15494 13376 15495
rect 13376 15494 13392 15495
rect 13410 15494 13462 15546
rect 13480 15494 13490 15546
rect 13490 15494 13532 15546
rect 13550 15494 13596 15546
rect 13596 15494 13602 15546
rect 4481 15438 4533 15490
rect 4545 15438 4597 15490
rect 4609 15438 4661 15490
rect 13200 15430 13252 15482
rect 13270 15430 13322 15482
rect 13340 15461 13342 15482
rect 13342 15461 13376 15482
rect 13376 15461 13392 15482
rect 13340 15430 13392 15461
rect 13410 15430 13462 15482
rect 13480 15430 13490 15482
rect 13490 15430 13532 15482
rect 13550 15430 13596 15482
rect 13596 15430 13602 15482
rect 13200 15366 13252 15418
rect 13270 15366 13322 15418
rect 13340 15385 13342 15418
rect 13342 15385 13376 15418
rect 13376 15385 13392 15418
rect 13340 15366 13392 15385
rect 13410 15366 13462 15418
rect 13480 15366 13490 15418
rect 13490 15366 13532 15418
rect 13550 15366 13596 15418
rect 13596 15366 13602 15418
rect 4481 15294 4533 15346
rect 4545 15294 4597 15346
rect 4609 15294 4661 15346
rect 13200 15302 13252 15354
rect 13270 15302 13322 15354
rect 13340 15343 13392 15354
rect 13340 15309 13342 15343
rect 13342 15309 13376 15343
rect 13376 15309 13392 15343
rect 13340 15302 13392 15309
rect 13410 15302 13462 15354
rect 13480 15302 13490 15354
rect 13490 15302 13532 15354
rect 13550 15302 13596 15354
rect 13596 15302 13602 15354
rect 13200 15238 13252 15290
rect 13270 15238 13322 15290
rect 13340 15267 13392 15290
rect 13340 15238 13342 15267
rect 13342 15238 13376 15267
rect 13376 15238 13392 15267
rect 13410 15238 13462 15290
rect 13480 15238 13490 15290
rect 13490 15238 13532 15290
rect 13550 15238 13596 15290
rect 13596 15238 13602 15290
rect 4481 15150 4533 15202
rect 4545 15150 4597 15202
rect 4609 15150 4661 15202
rect 13200 15174 13252 15226
rect 13270 15174 13322 15226
rect 13340 15191 13392 15226
rect 13340 15174 13342 15191
rect 13342 15174 13376 15191
rect 13376 15174 13392 15191
rect 13410 15174 13462 15226
rect 13480 15174 13490 15226
rect 13490 15174 13532 15226
rect 13550 15174 13596 15226
rect 13596 15174 13602 15226
rect 13200 15110 13252 15162
rect 13270 15110 13322 15162
rect 13340 15157 13342 15162
rect 13342 15157 13376 15162
rect 13376 15157 13392 15162
rect 13340 15110 13392 15157
rect 13410 15110 13462 15162
rect 13480 15110 13490 15162
rect 13490 15110 13532 15162
rect 13550 15110 13596 15162
rect 13596 15110 13602 15162
rect 4731 14990 4783 15042
rect 4797 14990 4849 15042
rect 13200 15046 13252 15098
rect 13270 15046 13322 15098
rect 13340 15046 13392 15098
rect 13410 15046 13462 15098
rect 13480 15046 13490 15098
rect 13490 15046 13532 15098
rect 13550 15046 13596 15098
rect 13596 15046 13602 15098
rect 13200 14982 13252 15034
rect 13270 14982 13322 15034
rect 13340 14982 13392 15034
rect 13410 14982 13462 15034
rect 13480 14982 13490 15034
rect 13490 14982 13532 15034
rect 13550 14982 13596 15034
rect 13596 14982 13602 15034
rect 4731 14869 4783 14921
rect 4797 14869 4849 14921
rect 13200 14918 13252 14970
rect 13270 14918 13322 14970
rect 13340 14918 13392 14970
rect 13410 14918 13462 14970
rect 13480 14918 13490 14970
rect 13490 14918 13532 14970
rect 13550 14918 13596 14970
rect 13596 14918 13602 14970
rect 13200 14854 13252 14906
rect 13270 14854 13322 14906
rect 13340 14854 13392 14906
rect 13410 14854 13462 14906
rect 13480 14854 13490 14906
rect 13490 14854 13532 14906
rect 13550 14854 13596 14906
rect 13596 14854 13602 14906
rect 13200 14790 13252 14842
rect 13270 14790 13322 14842
rect 13340 14790 13392 14842
rect 13410 14790 13462 14842
rect 13480 14790 13490 14842
rect 13490 14790 13532 14842
rect 13550 14790 13596 14842
rect 13596 14790 13602 14842
rect 13200 14726 13252 14778
rect 13270 14726 13322 14778
rect 13340 14726 13392 14778
rect 13410 14726 13462 14778
rect 13480 14726 13490 14778
rect 13490 14726 13532 14778
rect 13550 14726 13596 14778
rect 13596 14726 13602 14778
rect 3227 14668 3279 14720
rect 3293 14668 3345 14720
rect 3227 14602 3279 14654
rect 3293 14602 3345 14654
rect 3227 14536 3279 14588
rect 3293 14536 3345 14588
rect 3227 14470 3279 14522
rect 3293 14470 3345 14522
rect 3227 14404 3279 14456
rect 3293 14404 3345 14456
rect 2950 13877 3002 13892
rect 2950 13843 2956 13877
rect 2956 13843 2990 13877
rect 2990 13843 3002 13877
rect 2950 13840 3002 13843
rect 3016 13877 3068 13892
rect 3016 13843 3028 13877
rect 3028 13843 3062 13877
rect 3062 13843 3068 13877
rect 3016 13840 3068 13843
rect 2950 13799 3002 13826
rect 2950 13774 2956 13799
rect 2956 13774 2990 13799
rect 2990 13774 3002 13799
rect 3016 13799 3068 13826
rect 3016 13774 3028 13799
rect 3028 13774 3062 13799
rect 3062 13774 3068 13799
rect 2950 13722 3002 13760
rect 2950 13708 2956 13722
rect 2956 13708 2990 13722
rect 2990 13708 3002 13722
rect 3016 13722 3068 13760
rect 3016 13708 3028 13722
rect 3028 13708 3062 13722
rect 3062 13708 3068 13722
rect 2950 13688 2956 13694
rect 2956 13688 2990 13694
rect 2990 13688 3002 13694
rect 2950 13645 3002 13688
rect 2950 13642 2956 13645
rect 2956 13642 2990 13645
rect 2990 13642 3002 13645
rect 3016 13688 3028 13694
rect 3028 13688 3062 13694
rect 3062 13688 3068 13694
rect 3016 13645 3068 13688
rect 3016 13642 3028 13645
rect 3028 13642 3062 13645
rect 3062 13642 3068 13645
rect 2950 13611 2956 13628
rect 2956 13611 2990 13628
rect 2990 13611 3002 13628
rect 2950 13576 3002 13611
rect 3016 13611 3028 13628
rect 3028 13611 3062 13628
rect 3062 13611 3068 13628
rect 3016 13576 3068 13611
rect 2950 13534 2956 13562
rect 2956 13534 2990 13562
rect 2990 13534 3002 13562
rect 2950 13510 3002 13534
rect 3016 13534 3028 13562
rect 3028 13534 3062 13562
rect 3062 13534 3068 13562
rect 3016 13510 3068 13534
rect 2950 13491 3002 13495
rect 2950 13457 2956 13491
rect 2956 13457 2990 13491
rect 2990 13457 3002 13491
rect 2950 13443 3002 13457
rect 3016 13491 3068 13495
rect 3016 13457 3028 13491
rect 3028 13457 3062 13491
rect 3062 13457 3068 13491
rect 3016 13443 3068 13457
rect 2950 13414 3002 13428
rect 2950 13380 2956 13414
rect 2956 13380 2990 13414
rect 2990 13380 3002 13414
rect 2950 13376 3002 13380
rect 3016 13414 3068 13428
rect 3016 13380 3028 13414
rect 3028 13380 3062 13414
rect 3062 13380 3068 13414
rect 3016 13376 3068 13380
rect 2950 11840 2956 11892
rect 2956 11840 3002 11892
rect 3016 11840 3062 11892
rect 3062 11840 3068 11892
rect 2950 11774 2956 11826
rect 2956 11774 3002 11826
rect 3016 11774 3062 11826
rect 3062 11774 3068 11826
rect 2950 11708 2956 11760
rect 2956 11708 3002 11760
rect 3016 11708 3062 11760
rect 3062 11708 3068 11760
rect 2950 11642 2956 11694
rect 2956 11642 3002 11694
rect 3016 11642 3062 11694
rect 3062 11642 3068 11694
rect 2950 11576 2956 11628
rect 2956 11576 3002 11628
rect 3016 11576 3062 11628
rect 3062 11576 3068 11628
rect 2950 11510 2956 11562
rect 2956 11510 3002 11562
rect 3016 11510 3062 11562
rect 3062 11510 3068 11562
rect 2950 11443 2956 11495
rect 2956 11443 3002 11495
rect 3016 11443 3062 11495
rect 3062 11443 3068 11495
rect 2950 11380 2956 11428
rect 2956 11380 3002 11428
rect 3016 11380 3062 11428
rect 3062 11380 3068 11428
rect 2950 11376 3002 11380
rect 3016 11376 3068 11380
rect 2950 9844 2956 9896
rect 2956 9844 3002 9896
rect 3016 9844 3062 9896
rect 3062 9844 3068 9896
rect 2950 9778 2956 9830
rect 2956 9778 3002 9830
rect 3016 9778 3062 9830
rect 3062 9778 3068 9830
rect 2950 9712 2956 9764
rect 2956 9712 3002 9764
rect 3016 9712 3062 9764
rect 3062 9712 3068 9764
rect 2950 9646 2956 9698
rect 2956 9646 3002 9698
rect 3016 9646 3062 9698
rect 3062 9646 3068 9698
rect 2950 9580 2956 9632
rect 2956 9580 3002 9632
rect 3016 9580 3062 9632
rect 3062 9580 3068 9632
rect 2950 9514 2956 9566
rect 2956 9514 3002 9566
rect 3016 9514 3062 9566
rect 3062 9514 3068 9566
rect 2950 9447 2956 9499
rect 2956 9447 3002 9499
rect 3016 9447 3062 9499
rect 3062 9447 3068 9499
rect 2950 9380 2956 9432
rect 2956 9380 3002 9432
rect 3016 9380 3062 9432
rect 3062 9380 3068 9432
rect 2950 7840 2956 7892
rect 2956 7840 3002 7892
rect 3016 7840 3062 7892
rect 3062 7840 3068 7892
rect 2950 7774 2956 7826
rect 2956 7774 3002 7826
rect 3016 7774 3062 7826
rect 3062 7774 3068 7826
rect 2950 7708 2956 7760
rect 2956 7708 3002 7760
rect 3016 7708 3062 7760
rect 3062 7708 3068 7760
rect 2950 7642 2956 7694
rect 2956 7642 3002 7694
rect 3016 7642 3062 7694
rect 3062 7642 3068 7694
rect 2950 7576 2956 7628
rect 2956 7576 3002 7628
rect 3016 7576 3062 7628
rect 3062 7576 3068 7628
rect 2950 7510 2956 7562
rect 2956 7510 3002 7562
rect 3016 7510 3062 7562
rect 3062 7510 3068 7562
rect 2950 7443 2956 7495
rect 2956 7443 3002 7495
rect 3016 7443 3062 7495
rect 3062 7443 3068 7495
rect 2950 7380 2956 7428
rect 2956 7380 3002 7428
rect 3016 7380 3062 7428
rect 3062 7380 3068 7428
rect 2950 7376 3002 7380
rect 3016 7376 3068 7380
rect 2950 5844 2956 5896
rect 2956 5844 3002 5896
rect 3016 5844 3062 5896
rect 3062 5844 3068 5896
rect 2950 5778 2956 5830
rect 2956 5778 3002 5830
rect 3016 5778 3062 5830
rect 3062 5778 3068 5830
rect 2950 5712 2956 5764
rect 2956 5712 3002 5764
rect 3016 5712 3062 5764
rect 3062 5712 3068 5764
rect 2950 5646 2956 5698
rect 2956 5646 3002 5698
rect 3016 5646 3062 5698
rect 3062 5646 3068 5698
rect 2950 5580 2956 5632
rect 2956 5580 3002 5632
rect 3016 5580 3062 5632
rect 3062 5580 3068 5632
rect 2950 5514 2956 5566
rect 2956 5514 3002 5566
rect 3016 5514 3062 5566
rect 3062 5514 3068 5566
rect 2950 5447 2956 5499
rect 2956 5447 3002 5499
rect 3016 5447 3062 5499
rect 3062 5447 3068 5499
rect 2950 5380 2956 5432
rect 2956 5380 3002 5432
rect 3016 5380 3062 5432
rect 3062 5380 3068 5432
rect 3227 14345 3279 14390
rect 3227 14338 3233 14345
rect 3233 14338 3267 14345
rect 3267 14338 3279 14345
rect 3293 14345 3345 14390
rect 3781 14668 3833 14720
rect 3847 14668 3899 14720
rect 3781 14602 3833 14654
rect 3847 14602 3899 14654
rect 3781 14536 3833 14588
rect 3847 14536 3899 14588
rect 3781 14470 3833 14522
rect 3847 14470 3899 14522
rect 3781 14404 3833 14456
rect 3847 14404 3899 14456
rect 3293 14338 3305 14345
rect 3305 14338 3339 14345
rect 3339 14338 3345 14345
rect 3227 14311 3233 14323
rect 3233 14311 3267 14323
rect 3267 14311 3279 14323
rect 3227 14271 3279 14311
rect 3293 14311 3305 14323
rect 3305 14311 3339 14323
rect 3339 14311 3345 14323
rect 3293 14271 3345 14311
rect 3227 14233 3233 14256
rect 3233 14233 3267 14256
rect 3267 14233 3279 14256
rect 3227 14204 3279 14233
rect 3293 14233 3305 14256
rect 3305 14233 3339 14256
rect 3339 14233 3345 14256
rect 3293 14204 3345 14233
rect 3227 12714 3279 12720
rect 3227 12680 3233 12714
rect 3233 12680 3267 12714
rect 3267 12680 3279 12714
rect 3227 12668 3279 12680
rect 3293 12714 3345 12720
rect 3293 12680 3305 12714
rect 3305 12680 3339 12714
rect 3339 12680 3345 12714
rect 3293 12668 3345 12680
rect 3227 12641 3279 12654
rect 3227 12607 3233 12641
rect 3233 12607 3267 12641
rect 3267 12607 3279 12641
rect 3227 12602 3279 12607
rect 3293 12641 3345 12654
rect 3293 12607 3305 12641
rect 3305 12607 3339 12641
rect 3339 12607 3345 12641
rect 3293 12602 3345 12607
rect 3227 12568 3279 12588
rect 3227 12536 3233 12568
rect 3233 12536 3267 12568
rect 3267 12536 3279 12568
rect 3293 12568 3345 12588
rect 3293 12536 3305 12568
rect 3305 12536 3339 12568
rect 3339 12536 3345 12568
rect 3227 12495 3279 12522
rect 3227 12470 3233 12495
rect 3233 12470 3267 12495
rect 3267 12470 3279 12495
rect 3293 12495 3345 12522
rect 3293 12470 3305 12495
rect 3305 12470 3339 12495
rect 3339 12470 3345 12495
rect 3227 12422 3279 12456
rect 3293 12422 3345 12456
rect 3227 12404 3233 12422
rect 3233 12404 3279 12422
rect 3293 12404 3339 12422
rect 3339 12404 3345 12422
rect 3227 12338 3233 12390
rect 3233 12338 3279 12390
rect 3293 12338 3339 12390
rect 3339 12338 3345 12390
rect 3227 12271 3233 12323
rect 3233 12271 3279 12323
rect 3293 12271 3339 12323
rect 3339 12271 3345 12323
rect 3227 12204 3233 12256
rect 3233 12204 3279 12256
rect 3293 12204 3339 12256
rect 3339 12204 3345 12256
rect 3227 10714 3279 10724
rect 3227 10680 3233 10714
rect 3233 10680 3267 10714
rect 3267 10680 3279 10714
rect 3227 10672 3279 10680
rect 3293 10714 3345 10724
rect 3293 10680 3305 10714
rect 3305 10680 3339 10714
rect 3339 10680 3345 10714
rect 3293 10672 3345 10680
rect 3227 10641 3279 10658
rect 3227 10607 3233 10641
rect 3233 10607 3267 10641
rect 3267 10607 3279 10641
rect 3227 10606 3279 10607
rect 3293 10641 3345 10658
rect 3293 10607 3305 10641
rect 3305 10607 3339 10641
rect 3339 10607 3345 10641
rect 3293 10606 3345 10607
rect 3227 10568 3279 10592
rect 3227 10540 3233 10568
rect 3233 10540 3267 10568
rect 3267 10540 3279 10568
rect 3293 10568 3345 10592
rect 3293 10540 3305 10568
rect 3305 10540 3339 10568
rect 3339 10540 3345 10568
rect 3227 10495 3279 10526
rect 3227 10474 3233 10495
rect 3233 10474 3267 10495
rect 3267 10474 3279 10495
rect 3293 10495 3345 10526
rect 3293 10474 3305 10495
rect 3305 10474 3339 10495
rect 3339 10474 3345 10495
rect 3227 10422 3279 10460
rect 3293 10422 3345 10460
rect 3227 10408 3233 10422
rect 3233 10408 3279 10422
rect 3293 10408 3339 10422
rect 3339 10408 3345 10422
rect 3227 10342 3233 10394
rect 3233 10342 3279 10394
rect 3293 10342 3339 10394
rect 3339 10342 3345 10394
rect 3227 10275 3233 10327
rect 3233 10275 3279 10327
rect 3293 10275 3339 10327
rect 3339 10275 3345 10327
rect 3227 10208 3233 10260
rect 3233 10208 3279 10260
rect 3293 10208 3339 10260
rect 3339 10208 3345 10260
rect 3227 8714 3279 8720
rect 3227 8680 3233 8714
rect 3233 8680 3267 8714
rect 3267 8680 3279 8714
rect 3227 8668 3279 8680
rect 3293 8714 3345 8720
rect 3293 8680 3305 8714
rect 3305 8680 3339 8714
rect 3339 8680 3345 8714
rect 3293 8668 3345 8680
rect 3227 8641 3279 8654
rect 3227 8607 3233 8641
rect 3233 8607 3267 8641
rect 3267 8607 3279 8641
rect 3227 8602 3279 8607
rect 3293 8641 3345 8654
rect 3293 8607 3305 8641
rect 3305 8607 3339 8641
rect 3339 8607 3345 8641
rect 3293 8602 3345 8607
rect 3227 8568 3279 8588
rect 3227 8536 3233 8568
rect 3233 8536 3267 8568
rect 3267 8536 3279 8568
rect 3293 8568 3345 8588
rect 3293 8536 3305 8568
rect 3305 8536 3339 8568
rect 3339 8536 3345 8568
rect 3227 8495 3279 8522
rect 3227 8470 3233 8495
rect 3233 8470 3267 8495
rect 3267 8470 3279 8495
rect 3293 8495 3345 8522
rect 3293 8470 3305 8495
rect 3305 8470 3339 8495
rect 3339 8470 3345 8495
rect 3227 8422 3279 8456
rect 3293 8422 3345 8456
rect 3227 8404 3233 8422
rect 3233 8404 3279 8422
rect 3293 8404 3339 8422
rect 3339 8404 3345 8422
rect 3227 8338 3233 8390
rect 3233 8338 3279 8390
rect 3293 8338 3339 8390
rect 3339 8338 3345 8390
rect 3227 8271 3233 8323
rect 3233 8271 3279 8323
rect 3293 8271 3339 8323
rect 3339 8271 3345 8323
rect 3227 8204 3233 8256
rect 3233 8204 3279 8256
rect 3293 8204 3339 8256
rect 3339 8204 3345 8256
rect 3227 6714 3279 6724
rect 3227 6680 3233 6714
rect 3233 6680 3267 6714
rect 3267 6680 3279 6714
rect 3227 6672 3279 6680
rect 3293 6714 3345 6724
rect 3293 6680 3305 6714
rect 3305 6680 3339 6714
rect 3339 6680 3345 6714
rect 3293 6672 3345 6680
rect 3227 6641 3279 6658
rect 3227 6607 3233 6641
rect 3233 6607 3267 6641
rect 3267 6607 3279 6641
rect 3227 6606 3279 6607
rect 3293 6641 3345 6658
rect 3293 6607 3305 6641
rect 3305 6607 3339 6641
rect 3339 6607 3345 6641
rect 3293 6606 3345 6607
rect 3227 6568 3279 6592
rect 3227 6540 3233 6568
rect 3233 6540 3267 6568
rect 3267 6540 3279 6568
rect 3293 6568 3345 6592
rect 3293 6540 3305 6568
rect 3305 6540 3339 6568
rect 3339 6540 3345 6568
rect 3227 6495 3279 6526
rect 3227 6474 3233 6495
rect 3233 6474 3267 6495
rect 3267 6474 3279 6495
rect 3293 6495 3345 6526
rect 3293 6474 3305 6495
rect 3305 6474 3339 6495
rect 3339 6474 3345 6495
rect 3227 6422 3279 6460
rect 3293 6422 3345 6460
rect 3227 6408 3233 6422
rect 3233 6408 3279 6422
rect 3293 6408 3339 6422
rect 3339 6408 3345 6422
rect 3227 6342 3233 6394
rect 3233 6342 3279 6394
rect 3293 6342 3339 6394
rect 3339 6342 3345 6394
rect 3227 6275 3233 6327
rect 3233 6275 3279 6327
rect 3293 6275 3339 6327
rect 3339 6275 3345 6327
rect 3227 6208 3233 6260
rect 3233 6208 3279 6260
rect 3293 6208 3339 6260
rect 3339 6208 3345 6260
rect 3504 13877 3556 13892
rect 3504 13843 3510 13877
rect 3510 13843 3544 13877
rect 3544 13843 3556 13877
rect 3504 13840 3556 13843
rect 3570 13877 3622 13892
rect 3570 13843 3582 13877
rect 3582 13843 3616 13877
rect 3616 13843 3622 13877
rect 3570 13840 3622 13843
rect 3504 13799 3556 13826
rect 3504 13774 3510 13799
rect 3510 13774 3544 13799
rect 3544 13774 3556 13799
rect 3570 13799 3622 13826
rect 3570 13774 3582 13799
rect 3582 13774 3616 13799
rect 3616 13774 3622 13799
rect 3504 13722 3556 13760
rect 3504 13708 3510 13722
rect 3510 13708 3544 13722
rect 3544 13708 3556 13722
rect 3570 13722 3622 13760
rect 3570 13708 3582 13722
rect 3582 13708 3616 13722
rect 3616 13708 3622 13722
rect 3504 13688 3510 13694
rect 3510 13688 3544 13694
rect 3544 13688 3556 13694
rect 3504 13645 3556 13688
rect 3504 13642 3510 13645
rect 3510 13642 3544 13645
rect 3544 13642 3556 13645
rect 3570 13688 3582 13694
rect 3582 13688 3616 13694
rect 3616 13688 3622 13694
rect 3570 13645 3622 13688
rect 3570 13642 3582 13645
rect 3582 13642 3616 13645
rect 3616 13642 3622 13645
rect 3504 13611 3510 13628
rect 3510 13611 3544 13628
rect 3544 13611 3556 13628
rect 3504 13576 3556 13611
rect 3570 13611 3582 13628
rect 3582 13611 3616 13628
rect 3616 13611 3622 13628
rect 3570 13576 3622 13611
rect 3504 13534 3510 13562
rect 3510 13534 3544 13562
rect 3544 13534 3556 13562
rect 3504 13510 3556 13534
rect 3570 13534 3582 13562
rect 3582 13534 3616 13562
rect 3616 13534 3622 13562
rect 3570 13510 3622 13534
rect 3504 13491 3556 13495
rect 3504 13457 3510 13491
rect 3510 13457 3544 13491
rect 3544 13457 3556 13491
rect 3504 13443 3556 13457
rect 3570 13491 3622 13495
rect 3570 13457 3582 13491
rect 3582 13457 3616 13491
rect 3616 13457 3622 13491
rect 3570 13443 3622 13457
rect 3504 13414 3556 13428
rect 3504 13380 3510 13414
rect 3510 13380 3544 13414
rect 3544 13380 3556 13414
rect 3504 13376 3556 13380
rect 3570 13414 3622 13428
rect 3570 13380 3582 13414
rect 3582 13380 3616 13414
rect 3616 13380 3622 13414
rect 3570 13376 3622 13380
rect 3504 11840 3510 11892
rect 3510 11840 3556 11892
rect 3570 11840 3616 11892
rect 3616 11840 3622 11892
rect 3504 11774 3510 11826
rect 3510 11774 3556 11826
rect 3570 11774 3616 11826
rect 3616 11774 3622 11826
rect 3504 11708 3510 11760
rect 3510 11708 3556 11760
rect 3570 11708 3616 11760
rect 3616 11708 3622 11760
rect 3504 11642 3510 11694
rect 3510 11642 3556 11694
rect 3570 11642 3616 11694
rect 3616 11642 3622 11694
rect 3504 11576 3510 11628
rect 3510 11576 3556 11628
rect 3570 11576 3616 11628
rect 3616 11576 3622 11628
rect 3504 11510 3510 11562
rect 3510 11510 3556 11562
rect 3570 11510 3616 11562
rect 3616 11510 3622 11562
rect 3504 11443 3510 11495
rect 3510 11443 3556 11495
rect 3570 11443 3616 11495
rect 3616 11443 3622 11495
rect 3504 11380 3510 11428
rect 3510 11380 3556 11428
rect 3570 11380 3616 11428
rect 3616 11380 3622 11428
rect 3504 11376 3556 11380
rect 3570 11376 3622 11380
rect 3504 9844 3510 9896
rect 3510 9844 3556 9896
rect 3570 9844 3616 9896
rect 3616 9844 3622 9896
rect 3504 9778 3510 9830
rect 3510 9778 3556 9830
rect 3570 9778 3616 9830
rect 3616 9778 3622 9830
rect 3504 9712 3510 9764
rect 3510 9712 3556 9764
rect 3570 9712 3616 9764
rect 3616 9712 3622 9764
rect 3504 9646 3510 9698
rect 3510 9646 3556 9698
rect 3570 9646 3616 9698
rect 3616 9646 3622 9698
rect 3504 9580 3510 9632
rect 3510 9580 3556 9632
rect 3570 9580 3616 9632
rect 3616 9580 3622 9632
rect 3504 9514 3510 9566
rect 3510 9514 3556 9566
rect 3570 9514 3616 9566
rect 3616 9514 3622 9566
rect 3504 9447 3510 9499
rect 3510 9447 3556 9499
rect 3570 9447 3616 9499
rect 3616 9447 3622 9499
rect 3504 9380 3510 9432
rect 3510 9380 3556 9432
rect 3570 9380 3616 9432
rect 3616 9380 3622 9432
rect 3504 7840 3510 7892
rect 3510 7840 3556 7892
rect 3570 7840 3616 7892
rect 3616 7840 3622 7892
rect 3504 7774 3510 7826
rect 3510 7774 3556 7826
rect 3570 7774 3616 7826
rect 3616 7774 3622 7826
rect 3504 7708 3510 7760
rect 3510 7708 3556 7760
rect 3570 7708 3616 7760
rect 3616 7708 3622 7760
rect 3504 7642 3510 7694
rect 3510 7642 3556 7694
rect 3570 7642 3616 7694
rect 3616 7642 3622 7694
rect 3504 7576 3510 7628
rect 3510 7576 3556 7628
rect 3570 7576 3616 7628
rect 3616 7576 3622 7628
rect 3504 7510 3510 7562
rect 3510 7510 3556 7562
rect 3570 7510 3616 7562
rect 3616 7510 3622 7562
rect 3504 7443 3510 7495
rect 3510 7443 3556 7495
rect 3570 7443 3616 7495
rect 3616 7443 3622 7495
rect 3504 7380 3510 7428
rect 3510 7380 3556 7428
rect 3570 7380 3616 7428
rect 3616 7380 3622 7428
rect 3504 7376 3556 7380
rect 3570 7376 3622 7380
rect 3504 5844 3510 5896
rect 3510 5844 3556 5896
rect 3570 5844 3616 5896
rect 3616 5844 3622 5896
rect 3504 5778 3510 5830
rect 3510 5778 3556 5830
rect 3570 5778 3616 5830
rect 3616 5778 3622 5830
rect 3504 5712 3510 5764
rect 3510 5712 3556 5764
rect 3570 5712 3616 5764
rect 3616 5712 3622 5764
rect 3504 5646 3510 5698
rect 3510 5646 3556 5698
rect 3570 5646 3616 5698
rect 3616 5646 3622 5698
rect 3504 5580 3510 5632
rect 3510 5580 3556 5632
rect 3570 5580 3616 5632
rect 3616 5580 3622 5632
rect 3504 5514 3510 5566
rect 3510 5514 3556 5566
rect 3570 5514 3616 5566
rect 3616 5514 3622 5566
rect 3504 5447 3510 5499
rect 3510 5447 3556 5499
rect 3570 5447 3616 5499
rect 3616 5447 3622 5499
rect 3504 5380 3510 5432
rect 3510 5380 3556 5432
rect 3570 5380 3616 5432
rect 3616 5380 3622 5432
rect 3781 14345 3833 14390
rect 3781 14338 3787 14345
rect 3787 14338 3821 14345
rect 3821 14338 3833 14345
rect 3847 14345 3899 14390
rect 4335 14668 4387 14720
rect 4401 14668 4453 14720
rect 4335 14602 4387 14654
rect 4401 14602 4453 14654
rect 4335 14536 4387 14588
rect 4401 14536 4453 14588
rect 4335 14470 4387 14522
rect 4401 14470 4453 14522
rect 4335 14404 4387 14456
rect 4401 14404 4453 14456
rect 3847 14338 3859 14345
rect 3859 14338 3893 14345
rect 3893 14338 3899 14345
rect 3781 14311 3787 14323
rect 3787 14311 3821 14323
rect 3821 14311 3833 14323
rect 3781 14271 3833 14311
rect 3847 14311 3859 14323
rect 3859 14311 3893 14323
rect 3893 14311 3899 14323
rect 3847 14271 3899 14311
rect 3781 14233 3787 14256
rect 3787 14233 3821 14256
rect 3821 14233 3833 14256
rect 3781 14204 3833 14233
rect 3847 14233 3859 14256
rect 3859 14233 3893 14256
rect 3893 14233 3899 14256
rect 3847 14204 3899 14233
rect 3781 12714 3833 12720
rect 3781 12680 3787 12714
rect 3787 12680 3821 12714
rect 3821 12680 3833 12714
rect 3781 12668 3833 12680
rect 3847 12714 3899 12720
rect 3847 12680 3859 12714
rect 3859 12680 3893 12714
rect 3893 12680 3899 12714
rect 3847 12668 3899 12680
rect 3781 12641 3833 12654
rect 3781 12607 3787 12641
rect 3787 12607 3821 12641
rect 3821 12607 3833 12641
rect 3781 12602 3833 12607
rect 3847 12641 3899 12654
rect 3847 12607 3859 12641
rect 3859 12607 3893 12641
rect 3893 12607 3899 12641
rect 3847 12602 3899 12607
rect 3781 12568 3833 12588
rect 3781 12536 3787 12568
rect 3787 12536 3821 12568
rect 3821 12536 3833 12568
rect 3847 12568 3899 12588
rect 3847 12536 3859 12568
rect 3859 12536 3893 12568
rect 3893 12536 3899 12568
rect 3781 12495 3833 12522
rect 3781 12470 3787 12495
rect 3787 12470 3821 12495
rect 3821 12470 3833 12495
rect 3847 12495 3899 12522
rect 3847 12470 3859 12495
rect 3859 12470 3893 12495
rect 3893 12470 3899 12495
rect 3781 12422 3833 12456
rect 3847 12422 3899 12456
rect 3781 12404 3787 12422
rect 3787 12404 3833 12422
rect 3847 12404 3893 12422
rect 3893 12404 3899 12422
rect 3781 12338 3787 12390
rect 3787 12338 3833 12390
rect 3847 12338 3893 12390
rect 3893 12338 3899 12390
rect 3781 12271 3787 12323
rect 3787 12271 3833 12323
rect 3847 12271 3893 12323
rect 3893 12271 3899 12323
rect 3781 12204 3787 12256
rect 3787 12204 3833 12256
rect 3847 12204 3893 12256
rect 3893 12204 3899 12256
rect 3781 10714 3833 10724
rect 3781 10680 3787 10714
rect 3787 10680 3821 10714
rect 3821 10680 3833 10714
rect 3781 10672 3833 10680
rect 3847 10714 3899 10724
rect 3847 10680 3859 10714
rect 3859 10680 3893 10714
rect 3893 10680 3899 10714
rect 3847 10672 3899 10680
rect 3781 10641 3833 10658
rect 3781 10607 3787 10641
rect 3787 10607 3821 10641
rect 3821 10607 3833 10641
rect 3781 10606 3833 10607
rect 3847 10641 3899 10658
rect 3847 10607 3859 10641
rect 3859 10607 3893 10641
rect 3893 10607 3899 10641
rect 3847 10606 3899 10607
rect 3781 10568 3833 10592
rect 3781 10540 3787 10568
rect 3787 10540 3821 10568
rect 3821 10540 3833 10568
rect 3847 10568 3899 10592
rect 3847 10540 3859 10568
rect 3859 10540 3893 10568
rect 3893 10540 3899 10568
rect 3781 10495 3833 10526
rect 3781 10474 3787 10495
rect 3787 10474 3821 10495
rect 3821 10474 3833 10495
rect 3847 10495 3899 10526
rect 3847 10474 3859 10495
rect 3859 10474 3893 10495
rect 3893 10474 3899 10495
rect 3781 10422 3833 10460
rect 3847 10422 3899 10460
rect 3781 10408 3787 10422
rect 3787 10408 3833 10422
rect 3847 10408 3893 10422
rect 3893 10408 3899 10422
rect 3781 10342 3787 10394
rect 3787 10342 3833 10394
rect 3847 10342 3893 10394
rect 3893 10342 3899 10394
rect 3781 10275 3787 10327
rect 3787 10275 3833 10327
rect 3847 10275 3893 10327
rect 3893 10275 3899 10327
rect 3781 10208 3787 10260
rect 3787 10208 3833 10260
rect 3847 10208 3893 10260
rect 3893 10208 3899 10260
rect 3781 8714 3833 8720
rect 3781 8680 3787 8714
rect 3787 8680 3821 8714
rect 3821 8680 3833 8714
rect 3781 8668 3833 8680
rect 3847 8714 3899 8720
rect 3847 8680 3859 8714
rect 3859 8680 3893 8714
rect 3893 8680 3899 8714
rect 3847 8668 3899 8680
rect 3781 8641 3833 8654
rect 3781 8607 3787 8641
rect 3787 8607 3821 8641
rect 3821 8607 3833 8641
rect 3781 8602 3833 8607
rect 3847 8641 3899 8654
rect 3847 8607 3859 8641
rect 3859 8607 3893 8641
rect 3893 8607 3899 8641
rect 3847 8602 3899 8607
rect 3781 8568 3833 8588
rect 3781 8536 3787 8568
rect 3787 8536 3821 8568
rect 3821 8536 3833 8568
rect 3847 8568 3899 8588
rect 3847 8536 3859 8568
rect 3859 8536 3893 8568
rect 3893 8536 3899 8568
rect 3781 8495 3833 8522
rect 3781 8470 3787 8495
rect 3787 8470 3821 8495
rect 3821 8470 3833 8495
rect 3847 8495 3899 8522
rect 3847 8470 3859 8495
rect 3859 8470 3893 8495
rect 3893 8470 3899 8495
rect 3781 8422 3833 8456
rect 3847 8422 3899 8456
rect 3781 8404 3787 8422
rect 3787 8404 3833 8422
rect 3847 8404 3893 8422
rect 3893 8404 3899 8422
rect 3781 8338 3787 8390
rect 3787 8338 3833 8390
rect 3847 8338 3893 8390
rect 3893 8338 3899 8390
rect 3781 8271 3787 8323
rect 3787 8271 3833 8323
rect 3847 8271 3893 8323
rect 3893 8271 3899 8323
rect 3781 8204 3787 8256
rect 3787 8204 3833 8256
rect 3847 8204 3893 8256
rect 3893 8204 3899 8256
rect 3781 6714 3833 6724
rect 3781 6680 3787 6714
rect 3787 6680 3821 6714
rect 3821 6680 3833 6714
rect 3781 6672 3833 6680
rect 3847 6714 3899 6724
rect 3847 6680 3859 6714
rect 3859 6680 3893 6714
rect 3893 6680 3899 6714
rect 3847 6672 3899 6680
rect 3781 6641 3833 6658
rect 3781 6607 3787 6641
rect 3787 6607 3821 6641
rect 3821 6607 3833 6641
rect 3781 6606 3833 6607
rect 3847 6641 3899 6658
rect 3847 6607 3859 6641
rect 3859 6607 3893 6641
rect 3893 6607 3899 6641
rect 3847 6606 3899 6607
rect 3781 6568 3833 6592
rect 3781 6540 3787 6568
rect 3787 6540 3821 6568
rect 3821 6540 3833 6568
rect 3847 6568 3899 6592
rect 3847 6540 3859 6568
rect 3859 6540 3893 6568
rect 3893 6540 3899 6568
rect 3781 6495 3833 6526
rect 3781 6474 3787 6495
rect 3787 6474 3821 6495
rect 3821 6474 3833 6495
rect 3847 6495 3899 6526
rect 3847 6474 3859 6495
rect 3859 6474 3893 6495
rect 3893 6474 3899 6495
rect 3781 6422 3833 6460
rect 3847 6422 3899 6460
rect 3781 6408 3787 6422
rect 3787 6408 3833 6422
rect 3847 6408 3893 6422
rect 3893 6408 3899 6422
rect 3781 6342 3787 6394
rect 3787 6342 3833 6394
rect 3847 6342 3893 6394
rect 3893 6342 3899 6394
rect 3781 6275 3787 6327
rect 3787 6275 3833 6327
rect 3847 6275 3893 6327
rect 3893 6275 3899 6327
rect 3781 6208 3787 6260
rect 3787 6208 3833 6260
rect 3847 6208 3893 6260
rect 3893 6208 3899 6260
rect 4058 13877 4110 13892
rect 4058 13843 4064 13877
rect 4064 13843 4098 13877
rect 4098 13843 4110 13877
rect 4058 13840 4110 13843
rect 4124 13877 4176 13892
rect 4124 13843 4136 13877
rect 4136 13843 4170 13877
rect 4170 13843 4176 13877
rect 4124 13840 4176 13843
rect 4058 13799 4110 13826
rect 4058 13774 4064 13799
rect 4064 13774 4098 13799
rect 4098 13774 4110 13799
rect 4124 13799 4176 13826
rect 4124 13774 4136 13799
rect 4136 13774 4170 13799
rect 4170 13774 4176 13799
rect 4058 13722 4110 13760
rect 4058 13708 4064 13722
rect 4064 13708 4098 13722
rect 4098 13708 4110 13722
rect 4124 13722 4176 13760
rect 4124 13708 4136 13722
rect 4136 13708 4170 13722
rect 4170 13708 4176 13722
rect 4058 13688 4064 13694
rect 4064 13688 4098 13694
rect 4098 13688 4110 13694
rect 4058 13645 4110 13688
rect 4058 13642 4064 13645
rect 4064 13642 4098 13645
rect 4098 13642 4110 13645
rect 4124 13688 4136 13694
rect 4136 13688 4170 13694
rect 4170 13688 4176 13694
rect 4124 13645 4176 13688
rect 4124 13642 4136 13645
rect 4136 13642 4170 13645
rect 4170 13642 4176 13645
rect 4058 13611 4064 13628
rect 4064 13611 4098 13628
rect 4098 13611 4110 13628
rect 4058 13576 4110 13611
rect 4124 13611 4136 13628
rect 4136 13611 4170 13628
rect 4170 13611 4176 13628
rect 4124 13576 4176 13611
rect 4058 13534 4064 13562
rect 4064 13534 4098 13562
rect 4098 13534 4110 13562
rect 4058 13510 4110 13534
rect 4124 13534 4136 13562
rect 4136 13534 4170 13562
rect 4170 13534 4176 13562
rect 4124 13510 4176 13534
rect 4058 13491 4110 13495
rect 4058 13457 4064 13491
rect 4064 13457 4098 13491
rect 4098 13457 4110 13491
rect 4058 13443 4110 13457
rect 4124 13491 4176 13495
rect 4124 13457 4136 13491
rect 4136 13457 4170 13491
rect 4170 13457 4176 13491
rect 4124 13443 4176 13457
rect 4058 13414 4110 13428
rect 4058 13380 4064 13414
rect 4064 13380 4098 13414
rect 4098 13380 4110 13414
rect 4058 13376 4110 13380
rect 4124 13414 4176 13428
rect 4124 13380 4136 13414
rect 4136 13380 4170 13414
rect 4170 13380 4176 13414
rect 4124 13376 4176 13380
rect 4058 11840 4064 11892
rect 4064 11840 4110 11892
rect 4124 11840 4170 11892
rect 4170 11840 4176 11892
rect 4058 11774 4064 11826
rect 4064 11774 4110 11826
rect 4124 11774 4170 11826
rect 4170 11774 4176 11826
rect 4058 11708 4064 11760
rect 4064 11708 4110 11760
rect 4124 11708 4170 11760
rect 4170 11708 4176 11760
rect 4058 11642 4064 11694
rect 4064 11642 4110 11694
rect 4124 11642 4170 11694
rect 4170 11642 4176 11694
rect 4058 11576 4064 11628
rect 4064 11576 4110 11628
rect 4124 11576 4170 11628
rect 4170 11576 4176 11628
rect 4058 11510 4064 11562
rect 4064 11510 4110 11562
rect 4124 11510 4170 11562
rect 4170 11510 4176 11562
rect 4058 11443 4064 11495
rect 4064 11443 4110 11495
rect 4124 11443 4170 11495
rect 4170 11443 4176 11495
rect 4058 11380 4064 11428
rect 4064 11380 4110 11428
rect 4124 11380 4170 11428
rect 4170 11380 4176 11428
rect 4058 11376 4110 11380
rect 4124 11376 4176 11380
rect 4058 9844 4064 9896
rect 4064 9844 4110 9896
rect 4124 9844 4170 9896
rect 4170 9844 4176 9896
rect 4058 9778 4064 9830
rect 4064 9778 4110 9830
rect 4124 9778 4170 9830
rect 4170 9778 4176 9830
rect 4058 9712 4064 9764
rect 4064 9712 4110 9764
rect 4124 9712 4170 9764
rect 4170 9712 4176 9764
rect 4058 9646 4064 9698
rect 4064 9646 4110 9698
rect 4124 9646 4170 9698
rect 4170 9646 4176 9698
rect 4058 9580 4064 9632
rect 4064 9580 4110 9632
rect 4124 9580 4170 9632
rect 4170 9580 4176 9632
rect 4058 9514 4064 9566
rect 4064 9514 4110 9566
rect 4124 9514 4170 9566
rect 4170 9514 4176 9566
rect 4058 9447 4064 9499
rect 4064 9447 4110 9499
rect 4124 9447 4170 9499
rect 4170 9447 4176 9499
rect 4058 9380 4064 9432
rect 4064 9380 4110 9432
rect 4124 9380 4170 9432
rect 4170 9380 4176 9432
rect 4058 7840 4064 7892
rect 4064 7840 4110 7892
rect 4124 7840 4170 7892
rect 4170 7840 4176 7892
rect 4058 7774 4064 7826
rect 4064 7774 4110 7826
rect 4124 7774 4170 7826
rect 4170 7774 4176 7826
rect 4058 7708 4064 7760
rect 4064 7708 4110 7760
rect 4124 7708 4170 7760
rect 4170 7708 4176 7760
rect 4058 7642 4064 7694
rect 4064 7642 4110 7694
rect 4124 7642 4170 7694
rect 4170 7642 4176 7694
rect 4058 7576 4064 7628
rect 4064 7576 4110 7628
rect 4124 7576 4170 7628
rect 4170 7576 4176 7628
rect 4058 7510 4064 7562
rect 4064 7510 4110 7562
rect 4124 7510 4170 7562
rect 4170 7510 4176 7562
rect 4058 7443 4064 7495
rect 4064 7443 4110 7495
rect 4124 7443 4170 7495
rect 4170 7443 4176 7495
rect 4058 7380 4064 7428
rect 4064 7380 4110 7428
rect 4124 7380 4170 7428
rect 4170 7380 4176 7428
rect 4058 7376 4110 7380
rect 4124 7376 4176 7380
rect 4058 5844 4064 5896
rect 4064 5844 4110 5896
rect 4124 5844 4170 5896
rect 4170 5844 4176 5896
rect 4058 5778 4064 5830
rect 4064 5778 4110 5830
rect 4124 5778 4170 5830
rect 4170 5778 4176 5830
rect 4058 5712 4064 5764
rect 4064 5712 4110 5764
rect 4124 5712 4170 5764
rect 4170 5712 4176 5764
rect 4058 5646 4064 5698
rect 4064 5646 4110 5698
rect 4124 5646 4170 5698
rect 4170 5646 4176 5698
rect 4058 5580 4064 5632
rect 4064 5580 4110 5632
rect 4124 5580 4170 5632
rect 4170 5580 4176 5632
rect 4058 5514 4064 5566
rect 4064 5514 4110 5566
rect 4124 5514 4170 5566
rect 4170 5514 4176 5566
rect 4058 5447 4064 5499
rect 4064 5447 4110 5499
rect 4124 5447 4170 5499
rect 4170 5447 4176 5499
rect 4058 5380 4064 5432
rect 4064 5380 4110 5432
rect 4124 5380 4170 5432
rect 4170 5380 4176 5432
rect 4335 14345 4387 14390
rect 4335 14338 4341 14345
rect 4341 14338 4375 14345
rect 4375 14338 4387 14345
rect 4401 14345 4453 14390
rect 4889 14668 4941 14720
rect 4955 14668 5007 14720
rect 4889 14602 4941 14654
rect 4955 14602 5007 14654
rect 4889 14536 4941 14588
rect 4955 14536 5007 14588
rect 4889 14470 4941 14522
rect 4955 14470 5007 14522
rect 4889 14404 4941 14456
rect 4955 14404 5007 14456
rect 4401 14338 4413 14345
rect 4413 14338 4447 14345
rect 4447 14338 4453 14345
rect 4335 14311 4341 14323
rect 4341 14311 4375 14323
rect 4375 14311 4387 14323
rect 4335 14271 4387 14311
rect 4401 14311 4413 14323
rect 4413 14311 4447 14323
rect 4447 14311 4453 14323
rect 4401 14271 4453 14311
rect 4335 14233 4341 14256
rect 4341 14233 4375 14256
rect 4375 14233 4387 14256
rect 4335 14204 4387 14233
rect 4401 14233 4413 14256
rect 4413 14233 4447 14256
rect 4447 14233 4453 14256
rect 4401 14204 4453 14233
rect 4335 12714 4387 12720
rect 4335 12680 4341 12714
rect 4341 12680 4375 12714
rect 4375 12680 4387 12714
rect 4335 12668 4387 12680
rect 4401 12714 4453 12720
rect 4401 12680 4413 12714
rect 4413 12680 4447 12714
rect 4447 12680 4453 12714
rect 4401 12668 4453 12680
rect 4335 12641 4387 12654
rect 4335 12607 4341 12641
rect 4341 12607 4375 12641
rect 4375 12607 4387 12641
rect 4335 12602 4387 12607
rect 4401 12641 4453 12654
rect 4401 12607 4413 12641
rect 4413 12607 4447 12641
rect 4447 12607 4453 12641
rect 4401 12602 4453 12607
rect 4335 12568 4387 12588
rect 4335 12536 4341 12568
rect 4341 12536 4375 12568
rect 4375 12536 4387 12568
rect 4401 12568 4453 12588
rect 4401 12536 4413 12568
rect 4413 12536 4447 12568
rect 4447 12536 4453 12568
rect 4335 12495 4387 12522
rect 4335 12470 4341 12495
rect 4341 12470 4375 12495
rect 4375 12470 4387 12495
rect 4401 12495 4453 12522
rect 4401 12470 4413 12495
rect 4413 12470 4447 12495
rect 4447 12470 4453 12495
rect 4335 12422 4387 12456
rect 4401 12422 4453 12456
rect 4335 12404 4341 12422
rect 4341 12404 4387 12422
rect 4401 12404 4447 12422
rect 4447 12404 4453 12422
rect 4335 12338 4341 12390
rect 4341 12338 4387 12390
rect 4401 12338 4447 12390
rect 4447 12338 4453 12390
rect 4335 12271 4341 12323
rect 4341 12271 4387 12323
rect 4401 12271 4447 12323
rect 4447 12271 4453 12323
rect 4335 12204 4341 12256
rect 4341 12204 4387 12256
rect 4401 12204 4447 12256
rect 4447 12204 4453 12256
rect 4335 10714 4387 10724
rect 4335 10680 4341 10714
rect 4341 10680 4375 10714
rect 4375 10680 4387 10714
rect 4335 10672 4387 10680
rect 4401 10714 4453 10724
rect 4401 10680 4413 10714
rect 4413 10680 4447 10714
rect 4447 10680 4453 10714
rect 4401 10672 4453 10680
rect 4335 10641 4387 10658
rect 4335 10607 4341 10641
rect 4341 10607 4375 10641
rect 4375 10607 4387 10641
rect 4335 10606 4387 10607
rect 4401 10641 4453 10658
rect 4401 10607 4413 10641
rect 4413 10607 4447 10641
rect 4447 10607 4453 10641
rect 4401 10606 4453 10607
rect 4335 10568 4387 10592
rect 4335 10540 4341 10568
rect 4341 10540 4375 10568
rect 4375 10540 4387 10568
rect 4401 10568 4453 10592
rect 4401 10540 4413 10568
rect 4413 10540 4447 10568
rect 4447 10540 4453 10568
rect 4335 10495 4387 10526
rect 4335 10474 4341 10495
rect 4341 10474 4375 10495
rect 4375 10474 4387 10495
rect 4401 10495 4453 10526
rect 4401 10474 4413 10495
rect 4413 10474 4447 10495
rect 4447 10474 4453 10495
rect 4335 10422 4387 10460
rect 4401 10422 4453 10460
rect 4335 10408 4341 10422
rect 4341 10408 4387 10422
rect 4401 10408 4447 10422
rect 4447 10408 4453 10422
rect 4335 10342 4341 10394
rect 4341 10342 4387 10394
rect 4401 10342 4447 10394
rect 4447 10342 4453 10394
rect 4335 10275 4341 10327
rect 4341 10275 4387 10327
rect 4401 10275 4447 10327
rect 4447 10275 4453 10327
rect 4335 10208 4341 10260
rect 4341 10208 4387 10260
rect 4401 10208 4447 10260
rect 4447 10208 4453 10260
rect 4335 8714 4387 8720
rect 4335 8680 4341 8714
rect 4341 8680 4375 8714
rect 4375 8680 4387 8714
rect 4335 8668 4387 8680
rect 4401 8714 4453 8720
rect 4401 8680 4413 8714
rect 4413 8680 4447 8714
rect 4447 8680 4453 8714
rect 4401 8668 4453 8680
rect 4335 8641 4387 8654
rect 4335 8607 4341 8641
rect 4341 8607 4375 8641
rect 4375 8607 4387 8641
rect 4335 8602 4387 8607
rect 4401 8641 4453 8654
rect 4401 8607 4413 8641
rect 4413 8607 4447 8641
rect 4447 8607 4453 8641
rect 4401 8602 4453 8607
rect 4335 8568 4387 8588
rect 4335 8536 4341 8568
rect 4341 8536 4375 8568
rect 4375 8536 4387 8568
rect 4401 8568 4453 8588
rect 4401 8536 4413 8568
rect 4413 8536 4447 8568
rect 4447 8536 4453 8568
rect 4335 8495 4387 8522
rect 4335 8470 4341 8495
rect 4341 8470 4375 8495
rect 4375 8470 4387 8495
rect 4401 8495 4453 8522
rect 4401 8470 4413 8495
rect 4413 8470 4447 8495
rect 4447 8470 4453 8495
rect 4335 8422 4387 8456
rect 4401 8422 4453 8456
rect 4335 8404 4341 8422
rect 4341 8404 4387 8422
rect 4401 8404 4447 8422
rect 4447 8404 4453 8422
rect 4335 8338 4341 8390
rect 4341 8338 4387 8390
rect 4401 8338 4447 8390
rect 4447 8338 4453 8390
rect 4335 8271 4341 8323
rect 4341 8271 4387 8323
rect 4401 8271 4447 8323
rect 4447 8271 4453 8323
rect 4335 8204 4341 8256
rect 4341 8204 4387 8256
rect 4401 8204 4447 8256
rect 4447 8204 4453 8256
rect 4335 6714 4387 6724
rect 4335 6680 4341 6714
rect 4341 6680 4375 6714
rect 4375 6680 4387 6714
rect 4335 6672 4387 6680
rect 4401 6714 4453 6724
rect 4401 6680 4413 6714
rect 4413 6680 4447 6714
rect 4447 6680 4453 6714
rect 4401 6672 4453 6680
rect 4335 6641 4387 6658
rect 4335 6607 4341 6641
rect 4341 6607 4375 6641
rect 4375 6607 4387 6641
rect 4335 6606 4387 6607
rect 4401 6641 4453 6658
rect 4401 6607 4413 6641
rect 4413 6607 4447 6641
rect 4447 6607 4453 6641
rect 4401 6606 4453 6607
rect 4335 6568 4387 6592
rect 4335 6540 4341 6568
rect 4341 6540 4375 6568
rect 4375 6540 4387 6568
rect 4401 6568 4453 6592
rect 4401 6540 4413 6568
rect 4413 6540 4447 6568
rect 4447 6540 4453 6568
rect 4335 6495 4387 6526
rect 4335 6474 4341 6495
rect 4341 6474 4375 6495
rect 4375 6474 4387 6495
rect 4401 6495 4453 6526
rect 4401 6474 4413 6495
rect 4413 6474 4447 6495
rect 4447 6474 4453 6495
rect 4335 6422 4387 6460
rect 4401 6422 4453 6460
rect 4335 6408 4341 6422
rect 4341 6408 4387 6422
rect 4401 6408 4447 6422
rect 4447 6408 4453 6422
rect 4335 6342 4341 6394
rect 4341 6342 4387 6394
rect 4401 6342 4447 6394
rect 4447 6342 4453 6394
rect 4335 6275 4341 6327
rect 4341 6275 4387 6327
rect 4401 6275 4447 6327
rect 4447 6275 4453 6327
rect 4335 6208 4341 6260
rect 4341 6208 4387 6260
rect 4401 6208 4447 6260
rect 4447 6208 4453 6260
rect 4612 13877 4664 13892
rect 4612 13843 4618 13877
rect 4618 13843 4652 13877
rect 4652 13843 4664 13877
rect 4612 13840 4664 13843
rect 4678 13877 4730 13892
rect 4678 13843 4690 13877
rect 4690 13843 4724 13877
rect 4724 13843 4730 13877
rect 4678 13840 4730 13843
rect 4612 13799 4664 13826
rect 4612 13774 4618 13799
rect 4618 13774 4652 13799
rect 4652 13774 4664 13799
rect 4678 13799 4730 13826
rect 4678 13774 4690 13799
rect 4690 13774 4724 13799
rect 4724 13774 4730 13799
rect 4612 13722 4664 13760
rect 4612 13708 4618 13722
rect 4618 13708 4652 13722
rect 4652 13708 4664 13722
rect 4678 13722 4730 13760
rect 4678 13708 4690 13722
rect 4690 13708 4724 13722
rect 4724 13708 4730 13722
rect 4612 13688 4618 13694
rect 4618 13688 4652 13694
rect 4652 13688 4664 13694
rect 4612 13645 4664 13688
rect 4612 13642 4618 13645
rect 4618 13642 4652 13645
rect 4652 13642 4664 13645
rect 4678 13688 4690 13694
rect 4690 13688 4724 13694
rect 4724 13688 4730 13694
rect 4678 13645 4730 13688
rect 4678 13642 4690 13645
rect 4690 13642 4724 13645
rect 4724 13642 4730 13645
rect 4612 13611 4618 13628
rect 4618 13611 4652 13628
rect 4652 13611 4664 13628
rect 4612 13576 4664 13611
rect 4678 13611 4690 13628
rect 4690 13611 4724 13628
rect 4724 13611 4730 13628
rect 4678 13576 4730 13611
rect 4612 13534 4618 13562
rect 4618 13534 4652 13562
rect 4652 13534 4664 13562
rect 4612 13510 4664 13534
rect 4678 13534 4690 13562
rect 4690 13534 4724 13562
rect 4724 13534 4730 13562
rect 4678 13510 4730 13534
rect 4612 13491 4664 13495
rect 4612 13457 4618 13491
rect 4618 13457 4652 13491
rect 4652 13457 4664 13491
rect 4612 13443 4664 13457
rect 4678 13491 4730 13495
rect 4678 13457 4690 13491
rect 4690 13457 4724 13491
rect 4724 13457 4730 13491
rect 4678 13443 4730 13457
rect 4612 13414 4664 13428
rect 4612 13380 4618 13414
rect 4618 13380 4652 13414
rect 4652 13380 4664 13414
rect 4612 13376 4664 13380
rect 4678 13414 4730 13428
rect 4678 13380 4690 13414
rect 4690 13380 4724 13414
rect 4724 13380 4730 13414
rect 4678 13376 4730 13380
rect 4612 11840 4618 11892
rect 4618 11840 4664 11892
rect 4678 11840 4724 11892
rect 4724 11840 4730 11892
rect 4612 11774 4618 11826
rect 4618 11774 4664 11826
rect 4678 11774 4724 11826
rect 4724 11774 4730 11826
rect 4612 11708 4618 11760
rect 4618 11708 4664 11760
rect 4678 11708 4724 11760
rect 4724 11708 4730 11760
rect 4612 11642 4618 11694
rect 4618 11642 4664 11694
rect 4678 11642 4724 11694
rect 4724 11642 4730 11694
rect 4612 11576 4618 11628
rect 4618 11576 4664 11628
rect 4678 11576 4724 11628
rect 4724 11576 4730 11628
rect 4612 11510 4618 11562
rect 4618 11510 4664 11562
rect 4678 11510 4724 11562
rect 4724 11510 4730 11562
rect 4612 11443 4618 11495
rect 4618 11443 4664 11495
rect 4678 11443 4724 11495
rect 4724 11443 4730 11495
rect 4612 11380 4618 11428
rect 4618 11380 4664 11428
rect 4678 11380 4724 11428
rect 4724 11380 4730 11428
rect 4612 11376 4664 11380
rect 4678 11376 4730 11380
rect 4612 9844 4618 9896
rect 4618 9844 4664 9896
rect 4678 9844 4724 9896
rect 4724 9844 4730 9896
rect 4612 9778 4618 9830
rect 4618 9778 4664 9830
rect 4678 9778 4724 9830
rect 4724 9778 4730 9830
rect 4612 9712 4618 9764
rect 4618 9712 4664 9764
rect 4678 9712 4724 9764
rect 4724 9712 4730 9764
rect 4612 9646 4618 9698
rect 4618 9646 4664 9698
rect 4678 9646 4724 9698
rect 4724 9646 4730 9698
rect 4612 9580 4618 9632
rect 4618 9580 4664 9632
rect 4678 9580 4724 9632
rect 4724 9580 4730 9632
rect 4612 9514 4618 9566
rect 4618 9514 4664 9566
rect 4678 9514 4724 9566
rect 4724 9514 4730 9566
rect 4612 9447 4618 9499
rect 4618 9447 4664 9499
rect 4678 9447 4724 9499
rect 4724 9447 4730 9499
rect 4612 9380 4618 9432
rect 4618 9380 4664 9432
rect 4678 9380 4724 9432
rect 4724 9380 4730 9432
rect 4612 7840 4618 7892
rect 4618 7840 4664 7892
rect 4678 7840 4724 7892
rect 4724 7840 4730 7892
rect 4612 7774 4618 7826
rect 4618 7774 4664 7826
rect 4678 7774 4724 7826
rect 4724 7774 4730 7826
rect 4612 7708 4618 7760
rect 4618 7708 4664 7760
rect 4678 7708 4724 7760
rect 4724 7708 4730 7760
rect 4612 7642 4618 7694
rect 4618 7642 4664 7694
rect 4678 7642 4724 7694
rect 4724 7642 4730 7694
rect 4612 7576 4618 7628
rect 4618 7576 4664 7628
rect 4678 7576 4724 7628
rect 4724 7576 4730 7628
rect 4612 7510 4618 7562
rect 4618 7510 4664 7562
rect 4678 7510 4724 7562
rect 4724 7510 4730 7562
rect 4612 7443 4618 7495
rect 4618 7443 4664 7495
rect 4678 7443 4724 7495
rect 4724 7443 4730 7495
rect 4612 7380 4618 7428
rect 4618 7380 4664 7428
rect 4678 7380 4724 7428
rect 4724 7380 4730 7428
rect 4612 7376 4664 7380
rect 4678 7376 4730 7380
rect 4612 5844 4618 5896
rect 4618 5844 4664 5896
rect 4678 5844 4724 5896
rect 4724 5844 4730 5896
rect 4612 5778 4618 5830
rect 4618 5778 4664 5830
rect 4678 5778 4724 5830
rect 4724 5778 4730 5830
rect 4612 5712 4618 5764
rect 4618 5712 4664 5764
rect 4678 5712 4724 5764
rect 4724 5712 4730 5764
rect 4612 5646 4618 5698
rect 4618 5646 4664 5698
rect 4678 5646 4724 5698
rect 4724 5646 4730 5698
rect 4612 5580 4618 5632
rect 4618 5580 4664 5632
rect 4678 5580 4724 5632
rect 4724 5580 4730 5632
rect 4612 5514 4618 5566
rect 4618 5514 4664 5566
rect 4678 5514 4724 5566
rect 4724 5514 4730 5566
rect 4612 5447 4618 5499
rect 4618 5447 4664 5499
rect 4678 5447 4724 5499
rect 4724 5447 4730 5499
rect 4612 5380 4618 5432
rect 4618 5380 4664 5432
rect 4678 5380 4724 5432
rect 4724 5380 4730 5432
rect 4889 14345 4941 14390
rect 4889 14338 4895 14345
rect 4895 14338 4929 14345
rect 4929 14338 4941 14345
rect 4955 14345 5007 14390
rect 5443 14668 5495 14720
rect 5509 14668 5561 14720
rect 5443 14602 5495 14654
rect 5509 14602 5561 14654
rect 5443 14536 5495 14588
rect 5509 14536 5561 14588
rect 5443 14470 5495 14522
rect 5509 14470 5561 14522
rect 5443 14404 5495 14456
rect 5509 14404 5561 14456
rect 4955 14338 4967 14345
rect 4967 14338 5001 14345
rect 5001 14338 5007 14345
rect 4889 14311 4895 14323
rect 4895 14311 4929 14323
rect 4929 14311 4941 14323
rect 4889 14271 4941 14311
rect 4955 14311 4967 14323
rect 4967 14311 5001 14323
rect 5001 14311 5007 14323
rect 4955 14271 5007 14311
rect 4889 14233 4895 14256
rect 4895 14233 4929 14256
rect 4929 14233 4941 14256
rect 4889 14204 4941 14233
rect 4955 14233 4967 14256
rect 4967 14233 5001 14256
rect 5001 14233 5007 14256
rect 4955 14204 5007 14233
rect 4889 12714 4941 12720
rect 4889 12680 4895 12714
rect 4895 12680 4929 12714
rect 4929 12680 4941 12714
rect 4889 12668 4941 12680
rect 4955 12714 5007 12720
rect 4955 12680 4967 12714
rect 4967 12680 5001 12714
rect 5001 12680 5007 12714
rect 4955 12668 5007 12680
rect 4889 12641 4941 12654
rect 4889 12607 4895 12641
rect 4895 12607 4929 12641
rect 4929 12607 4941 12641
rect 4889 12602 4941 12607
rect 4955 12641 5007 12654
rect 4955 12607 4967 12641
rect 4967 12607 5001 12641
rect 5001 12607 5007 12641
rect 4955 12602 5007 12607
rect 4889 12568 4941 12588
rect 4889 12536 4895 12568
rect 4895 12536 4929 12568
rect 4929 12536 4941 12568
rect 4955 12568 5007 12588
rect 4955 12536 4967 12568
rect 4967 12536 5001 12568
rect 5001 12536 5007 12568
rect 4889 12495 4941 12522
rect 4889 12470 4895 12495
rect 4895 12470 4929 12495
rect 4929 12470 4941 12495
rect 4955 12495 5007 12522
rect 4955 12470 4967 12495
rect 4967 12470 5001 12495
rect 5001 12470 5007 12495
rect 4889 12422 4941 12456
rect 4955 12422 5007 12456
rect 4889 12404 4895 12422
rect 4895 12404 4941 12422
rect 4955 12404 5001 12422
rect 5001 12404 5007 12422
rect 4889 12338 4895 12390
rect 4895 12338 4941 12390
rect 4955 12338 5001 12390
rect 5001 12338 5007 12390
rect 4889 12271 4895 12323
rect 4895 12271 4941 12323
rect 4955 12271 5001 12323
rect 5001 12271 5007 12323
rect 4889 12204 4895 12256
rect 4895 12204 4941 12256
rect 4955 12204 5001 12256
rect 5001 12204 5007 12256
rect 4889 10714 4941 10724
rect 4889 10680 4895 10714
rect 4895 10680 4929 10714
rect 4929 10680 4941 10714
rect 4889 10672 4941 10680
rect 4955 10714 5007 10724
rect 4955 10680 4967 10714
rect 4967 10680 5001 10714
rect 5001 10680 5007 10714
rect 4955 10672 5007 10680
rect 4889 10641 4941 10658
rect 4889 10607 4895 10641
rect 4895 10607 4929 10641
rect 4929 10607 4941 10641
rect 4889 10606 4941 10607
rect 4955 10641 5007 10658
rect 4955 10607 4967 10641
rect 4967 10607 5001 10641
rect 5001 10607 5007 10641
rect 4955 10606 5007 10607
rect 4889 10568 4941 10592
rect 4889 10540 4895 10568
rect 4895 10540 4929 10568
rect 4929 10540 4941 10568
rect 4955 10568 5007 10592
rect 4955 10540 4967 10568
rect 4967 10540 5001 10568
rect 5001 10540 5007 10568
rect 4889 10495 4941 10526
rect 4889 10474 4895 10495
rect 4895 10474 4929 10495
rect 4929 10474 4941 10495
rect 4955 10495 5007 10526
rect 4955 10474 4967 10495
rect 4967 10474 5001 10495
rect 5001 10474 5007 10495
rect 4889 10422 4941 10460
rect 4955 10422 5007 10460
rect 4889 10408 4895 10422
rect 4895 10408 4941 10422
rect 4955 10408 5001 10422
rect 5001 10408 5007 10422
rect 4889 10342 4895 10394
rect 4895 10342 4941 10394
rect 4955 10342 5001 10394
rect 5001 10342 5007 10394
rect 4889 10275 4895 10327
rect 4895 10275 4941 10327
rect 4955 10275 5001 10327
rect 5001 10275 5007 10327
rect 4889 10208 4895 10260
rect 4895 10208 4941 10260
rect 4955 10208 5001 10260
rect 5001 10208 5007 10260
rect 4889 8714 4941 8720
rect 4889 8680 4895 8714
rect 4895 8680 4929 8714
rect 4929 8680 4941 8714
rect 4889 8668 4941 8680
rect 4955 8714 5007 8720
rect 4955 8680 4967 8714
rect 4967 8680 5001 8714
rect 5001 8680 5007 8714
rect 4955 8668 5007 8680
rect 4889 8641 4941 8654
rect 4889 8607 4895 8641
rect 4895 8607 4929 8641
rect 4929 8607 4941 8641
rect 4889 8602 4941 8607
rect 4955 8641 5007 8654
rect 4955 8607 4967 8641
rect 4967 8607 5001 8641
rect 5001 8607 5007 8641
rect 4955 8602 5007 8607
rect 4889 8568 4941 8588
rect 4889 8536 4895 8568
rect 4895 8536 4929 8568
rect 4929 8536 4941 8568
rect 4955 8568 5007 8588
rect 4955 8536 4967 8568
rect 4967 8536 5001 8568
rect 5001 8536 5007 8568
rect 4889 8495 4941 8522
rect 4889 8470 4895 8495
rect 4895 8470 4929 8495
rect 4929 8470 4941 8495
rect 4955 8495 5007 8522
rect 4955 8470 4967 8495
rect 4967 8470 5001 8495
rect 5001 8470 5007 8495
rect 4889 8422 4941 8456
rect 4955 8422 5007 8456
rect 4889 8404 4895 8422
rect 4895 8404 4941 8422
rect 4955 8404 5001 8422
rect 5001 8404 5007 8422
rect 4889 8338 4895 8390
rect 4895 8338 4941 8390
rect 4955 8338 5001 8390
rect 5001 8338 5007 8390
rect 4889 8271 4895 8323
rect 4895 8271 4941 8323
rect 4955 8271 5001 8323
rect 5001 8271 5007 8323
rect 4889 8204 4895 8256
rect 4895 8204 4941 8256
rect 4955 8204 5001 8256
rect 5001 8204 5007 8256
rect 4889 6714 4941 6724
rect 4889 6680 4895 6714
rect 4895 6680 4929 6714
rect 4929 6680 4941 6714
rect 4889 6672 4941 6680
rect 4955 6714 5007 6724
rect 4955 6680 4967 6714
rect 4967 6680 5001 6714
rect 5001 6680 5007 6714
rect 4955 6672 5007 6680
rect 4889 6641 4941 6658
rect 4889 6607 4895 6641
rect 4895 6607 4929 6641
rect 4929 6607 4941 6641
rect 4889 6606 4941 6607
rect 4955 6641 5007 6658
rect 4955 6607 4967 6641
rect 4967 6607 5001 6641
rect 5001 6607 5007 6641
rect 4955 6606 5007 6607
rect 4889 6568 4941 6592
rect 4889 6540 4895 6568
rect 4895 6540 4929 6568
rect 4929 6540 4941 6568
rect 4955 6568 5007 6592
rect 4955 6540 4967 6568
rect 4967 6540 5001 6568
rect 5001 6540 5007 6568
rect 4889 6495 4941 6526
rect 4889 6474 4895 6495
rect 4895 6474 4929 6495
rect 4929 6474 4941 6495
rect 4955 6495 5007 6526
rect 4955 6474 4967 6495
rect 4967 6474 5001 6495
rect 5001 6474 5007 6495
rect 4889 6422 4941 6460
rect 4955 6422 5007 6460
rect 4889 6408 4895 6422
rect 4895 6408 4941 6422
rect 4955 6408 5001 6422
rect 5001 6408 5007 6422
rect 4889 6342 4895 6394
rect 4895 6342 4941 6394
rect 4955 6342 5001 6394
rect 5001 6342 5007 6394
rect 4889 6275 4895 6327
rect 4895 6275 4941 6327
rect 4955 6275 5001 6327
rect 5001 6275 5007 6327
rect 4889 6208 4895 6260
rect 4895 6208 4941 6260
rect 4955 6208 5001 6260
rect 5001 6208 5007 6260
rect 5166 13877 5218 13892
rect 5166 13843 5172 13877
rect 5172 13843 5206 13877
rect 5206 13843 5218 13877
rect 5166 13840 5218 13843
rect 5232 13877 5284 13892
rect 5232 13843 5244 13877
rect 5244 13843 5278 13877
rect 5278 13843 5284 13877
rect 5232 13840 5284 13843
rect 5166 13799 5218 13826
rect 5166 13774 5172 13799
rect 5172 13774 5206 13799
rect 5206 13774 5218 13799
rect 5232 13799 5284 13826
rect 5232 13774 5244 13799
rect 5244 13774 5278 13799
rect 5278 13774 5284 13799
rect 5166 13722 5218 13760
rect 5166 13708 5172 13722
rect 5172 13708 5206 13722
rect 5206 13708 5218 13722
rect 5232 13722 5284 13760
rect 5232 13708 5244 13722
rect 5244 13708 5278 13722
rect 5278 13708 5284 13722
rect 5166 13688 5172 13694
rect 5172 13688 5206 13694
rect 5206 13688 5218 13694
rect 5166 13645 5218 13688
rect 5166 13642 5172 13645
rect 5172 13642 5206 13645
rect 5206 13642 5218 13645
rect 5232 13688 5244 13694
rect 5244 13688 5278 13694
rect 5278 13688 5284 13694
rect 5232 13645 5284 13688
rect 5232 13642 5244 13645
rect 5244 13642 5278 13645
rect 5278 13642 5284 13645
rect 5166 13611 5172 13628
rect 5172 13611 5206 13628
rect 5206 13611 5218 13628
rect 5166 13576 5218 13611
rect 5232 13611 5244 13628
rect 5244 13611 5278 13628
rect 5278 13611 5284 13628
rect 5232 13576 5284 13611
rect 5166 13534 5172 13562
rect 5172 13534 5206 13562
rect 5206 13534 5218 13562
rect 5166 13510 5218 13534
rect 5232 13534 5244 13562
rect 5244 13534 5278 13562
rect 5278 13534 5284 13562
rect 5232 13510 5284 13534
rect 5166 13491 5218 13495
rect 5166 13457 5172 13491
rect 5172 13457 5206 13491
rect 5206 13457 5218 13491
rect 5166 13443 5218 13457
rect 5232 13491 5284 13495
rect 5232 13457 5244 13491
rect 5244 13457 5278 13491
rect 5278 13457 5284 13491
rect 5232 13443 5284 13457
rect 5166 13414 5218 13428
rect 5166 13380 5172 13414
rect 5172 13380 5206 13414
rect 5206 13380 5218 13414
rect 5166 13376 5218 13380
rect 5232 13414 5284 13428
rect 5232 13380 5244 13414
rect 5244 13380 5278 13414
rect 5278 13380 5284 13414
rect 5232 13376 5284 13380
rect 5166 11840 5172 11892
rect 5172 11840 5218 11892
rect 5232 11840 5278 11892
rect 5278 11840 5284 11892
rect 5166 11774 5172 11826
rect 5172 11774 5218 11826
rect 5232 11774 5278 11826
rect 5278 11774 5284 11826
rect 5166 11708 5172 11760
rect 5172 11708 5218 11760
rect 5232 11708 5278 11760
rect 5278 11708 5284 11760
rect 5166 11642 5172 11694
rect 5172 11642 5218 11694
rect 5232 11642 5278 11694
rect 5278 11642 5284 11694
rect 5166 11576 5172 11628
rect 5172 11576 5218 11628
rect 5232 11576 5278 11628
rect 5278 11576 5284 11628
rect 5166 11510 5172 11562
rect 5172 11510 5218 11562
rect 5232 11510 5278 11562
rect 5278 11510 5284 11562
rect 5166 11443 5172 11495
rect 5172 11443 5218 11495
rect 5232 11443 5278 11495
rect 5278 11443 5284 11495
rect 5166 11380 5172 11428
rect 5172 11380 5218 11428
rect 5232 11380 5278 11428
rect 5278 11380 5284 11428
rect 5166 11376 5218 11380
rect 5232 11376 5284 11380
rect 5166 9844 5172 9896
rect 5172 9844 5218 9896
rect 5232 9844 5278 9896
rect 5278 9844 5284 9896
rect 5166 9778 5172 9830
rect 5172 9778 5218 9830
rect 5232 9778 5278 9830
rect 5278 9778 5284 9830
rect 5166 9712 5172 9764
rect 5172 9712 5218 9764
rect 5232 9712 5278 9764
rect 5278 9712 5284 9764
rect 5166 9646 5172 9698
rect 5172 9646 5218 9698
rect 5232 9646 5278 9698
rect 5278 9646 5284 9698
rect 5166 9580 5172 9632
rect 5172 9580 5218 9632
rect 5232 9580 5278 9632
rect 5278 9580 5284 9632
rect 5166 9514 5172 9566
rect 5172 9514 5218 9566
rect 5232 9514 5278 9566
rect 5278 9514 5284 9566
rect 5166 9447 5172 9499
rect 5172 9447 5218 9499
rect 5232 9447 5278 9499
rect 5278 9447 5284 9499
rect 5166 9380 5172 9432
rect 5172 9380 5218 9432
rect 5232 9380 5278 9432
rect 5278 9380 5284 9432
rect 5166 7840 5172 7892
rect 5172 7840 5218 7892
rect 5232 7840 5278 7892
rect 5278 7840 5284 7892
rect 5166 7774 5172 7826
rect 5172 7774 5218 7826
rect 5232 7774 5278 7826
rect 5278 7774 5284 7826
rect 5166 7708 5172 7760
rect 5172 7708 5218 7760
rect 5232 7708 5278 7760
rect 5278 7708 5284 7760
rect 5166 7642 5172 7694
rect 5172 7642 5218 7694
rect 5232 7642 5278 7694
rect 5278 7642 5284 7694
rect 5166 7576 5172 7628
rect 5172 7576 5218 7628
rect 5232 7576 5278 7628
rect 5278 7576 5284 7628
rect 5166 7510 5172 7562
rect 5172 7510 5218 7562
rect 5232 7510 5278 7562
rect 5278 7510 5284 7562
rect 5166 7443 5172 7495
rect 5172 7443 5218 7495
rect 5232 7443 5278 7495
rect 5278 7443 5284 7495
rect 5166 7380 5172 7428
rect 5172 7380 5218 7428
rect 5232 7380 5278 7428
rect 5278 7380 5284 7428
rect 5166 7376 5218 7380
rect 5232 7376 5284 7380
rect 5166 5844 5172 5896
rect 5172 5844 5218 5896
rect 5232 5844 5278 5896
rect 5278 5844 5284 5896
rect 5166 5778 5172 5830
rect 5172 5778 5218 5830
rect 5232 5778 5278 5830
rect 5278 5778 5284 5830
rect 5166 5712 5172 5764
rect 5172 5712 5218 5764
rect 5232 5712 5278 5764
rect 5278 5712 5284 5764
rect 5166 5646 5172 5698
rect 5172 5646 5218 5698
rect 5232 5646 5278 5698
rect 5278 5646 5284 5698
rect 5166 5580 5172 5632
rect 5172 5580 5218 5632
rect 5232 5580 5278 5632
rect 5278 5580 5284 5632
rect 5166 5514 5172 5566
rect 5172 5514 5218 5566
rect 5232 5514 5278 5566
rect 5278 5514 5284 5566
rect 5166 5447 5172 5499
rect 5172 5447 5218 5499
rect 5232 5447 5278 5499
rect 5278 5447 5284 5499
rect 5166 5380 5172 5432
rect 5172 5380 5218 5432
rect 5232 5380 5278 5432
rect 5278 5380 5284 5432
rect 5443 14345 5495 14390
rect 5443 14338 5449 14345
rect 5449 14338 5483 14345
rect 5483 14338 5495 14345
rect 5509 14345 5561 14390
rect 5997 14668 6049 14720
rect 6063 14668 6115 14720
rect 5997 14602 6049 14654
rect 6063 14602 6115 14654
rect 5997 14536 6049 14588
rect 6063 14536 6115 14588
rect 5997 14470 6049 14522
rect 6063 14470 6115 14522
rect 5997 14404 6049 14456
rect 6063 14404 6115 14456
rect 5509 14338 5521 14345
rect 5521 14338 5555 14345
rect 5555 14338 5561 14345
rect 5443 14311 5449 14323
rect 5449 14311 5483 14323
rect 5483 14311 5495 14323
rect 5443 14271 5495 14311
rect 5509 14311 5521 14323
rect 5521 14311 5555 14323
rect 5555 14311 5561 14323
rect 5509 14271 5561 14311
rect 5443 14233 5449 14256
rect 5449 14233 5483 14256
rect 5483 14233 5495 14256
rect 5443 14204 5495 14233
rect 5509 14233 5521 14256
rect 5521 14233 5555 14256
rect 5555 14233 5561 14256
rect 5509 14204 5561 14233
rect 5443 12714 5495 12720
rect 5443 12680 5449 12714
rect 5449 12680 5483 12714
rect 5483 12680 5495 12714
rect 5443 12668 5495 12680
rect 5509 12714 5561 12720
rect 5509 12680 5521 12714
rect 5521 12680 5555 12714
rect 5555 12680 5561 12714
rect 5509 12668 5561 12680
rect 5443 12641 5495 12654
rect 5443 12607 5449 12641
rect 5449 12607 5483 12641
rect 5483 12607 5495 12641
rect 5443 12602 5495 12607
rect 5509 12641 5561 12654
rect 5509 12607 5521 12641
rect 5521 12607 5555 12641
rect 5555 12607 5561 12641
rect 5509 12602 5561 12607
rect 5443 12568 5495 12588
rect 5443 12536 5449 12568
rect 5449 12536 5483 12568
rect 5483 12536 5495 12568
rect 5509 12568 5561 12588
rect 5509 12536 5521 12568
rect 5521 12536 5555 12568
rect 5555 12536 5561 12568
rect 5443 12495 5495 12522
rect 5443 12470 5449 12495
rect 5449 12470 5483 12495
rect 5483 12470 5495 12495
rect 5509 12495 5561 12522
rect 5509 12470 5521 12495
rect 5521 12470 5555 12495
rect 5555 12470 5561 12495
rect 5443 12422 5495 12456
rect 5509 12422 5561 12456
rect 5443 12404 5449 12422
rect 5449 12404 5495 12422
rect 5509 12404 5555 12422
rect 5555 12404 5561 12422
rect 5443 12338 5449 12390
rect 5449 12338 5495 12390
rect 5509 12338 5555 12390
rect 5555 12338 5561 12390
rect 5443 12271 5449 12323
rect 5449 12271 5495 12323
rect 5509 12271 5555 12323
rect 5555 12271 5561 12323
rect 5443 12204 5449 12256
rect 5449 12204 5495 12256
rect 5509 12204 5555 12256
rect 5555 12204 5561 12256
rect 5443 10714 5495 10724
rect 5443 10680 5449 10714
rect 5449 10680 5483 10714
rect 5483 10680 5495 10714
rect 5443 10672 5495 10680
rect 5509 10714 5561 10724
rect 5509 10680 5521 10714
rect 5521 10680 5555 10714
rect 5555 10680 5561 10714
rect 5509 10672 5561 10680
rect 5443 10641 5495 10658
rect 5443 10607 5449 10641
rect 5449 10607 5483 10641
rect 5483 10607 5495 10641
rect 5443 10606 5495 10607
rect 5509 10641 5561 10658
rect 5509 10607 5521 10641
rect 5521 10607 5555 10641
rect 5555 10607 5561 10641
rect 5509 10606 5561 10607
rect 5443 10568 5495 10592
rect 5443 10540 5449 10568
rect 5449 10540 5483 10568
rect 5483 10540 5495 10568
rect 5509 10568 5561 10592
rect 5509 10540 5521 10568
rect 5521 10540 5555 10568
rect 5555 10540 5561 10568
rect 5443 10495 5495 10526
rect 5443 10474 5449 10495
rect 5449 10474 5483 10495
rect 5483 10474 5495 10495
rect 5509 10495 5561 10526
rect 5509 10474 5521 10495
rect 5521 10474 5555 10495
rect 5555 10474 5561 10495
rect 5443 10422 5495 10460
rect 5509 10422 5561 10460
rect 5443 10408 5449 10422
rect 5449 10408 5495 10422
rect 5509 10408 5555 10422
rect 5555 10408 5561 10422
rect 5443 10342 5449 10394
rect 5449 10342 5495 10394
rect 5509 10342 5555 10394
rect 5555 10342 5561 10394
rect 5443 10275 5449 10327
rect 5449 10275 5495 10327
rect 5509 10275 5555 10327
rect 5555 10275 5561 10327
rect 5443 10208 5449 10260
rect 5449 10208 5495 10260
rect 5509 10208 5555 10260
rect 5555 10208 5561 10260
rect 5443 8714 5495 8720
rect 5443 8680 5449 8714
rect 5449 8680 5483 8714
rect 5483 8680 5495 8714
rect 5443 8668 5495 8680
rect 5509 8714 5561 8720
rect 5509 8680 5521 8714
rect 5521 8680 5555 8714
rect 5555 8680 5561 8714
rect 5509 8668 5561 8680
rect 5443 8641 5495 8654
rect 5443 8607 5449 8641
rect 5449 8607 5483 8641
rect 5483 8607 5495 8641
rect 5443 8602 5495 8607
rect 5509 8641 5561 8654
rect 5509 8607 5521 8641
rect 5521 8607 5555 8641
rect 5555 8607 5561 8641
rect 5509 8602 5561 8607
rect 5443 8568 5495 8588
rect 5443 8536 5449 8568
rect 5449 8536 5483 8568
rect 5483 8536 5495 8568
rect 5509 8568 5561 8588
rect 5509 8536 5521 8568
rect 5521 8536 5555 8568
rect 5555 8536 5561 8568
rect 5443 8495 5495 8522
rect 5443 8470 5449 8495
rect 5449 8470 5483 8495
rect 5483 8470 5495 8495
rect 5509 8495 5561 8522
rect 5509 8470 5521 8495
rect 5521 8470 5555 8495
rect 5555 8470 5561 8495
rect 5443 8422 5495 8456
rect 5509 8422 5561 8456
rect 5443 8404 5449 8422
rect 5449 8404 5495 8422
rect 5509 8404 5555 8422
rect 5555 8404 5561 8422
rect 5443 8338 5449 8390
rect 5449 8338 5495 8390
rect 5509 8338 5555 8390
rect 5555 8338 5561 8390
rect 5443 8271 5449 8323
rect 5449 8271 5495 8323
rect 5509 8271 5555 8323
rect 5555 8271 5561 8323
rect 5443 8204 5449 8256
rect 5449 8204 5495 8256
rect 5509 8204 5555 8256
rect 5555 8204 5561 8256
rect 5443 6714 5495 6724
rect 5443 6680 5449 6714
rect 5449 6680 5483 6714
rect 5483 6680 5495 6714
rect 5443 6672 5495 6680
rect 5509 6714 5561 6724
rect 5509 6680 5521 6714
rect 5521 6680 5555 6714
rect 5555 6680 5561 6714
rect 5509 6672 5561 6680
rect 5443 6641 5495 6658
rect 5443 6607 5449 6641
rect 5449 6607 5483 6641
rect 5483 6607 5495 6641
rect 5443 6606 5495 6607
rect 5509 6641 5561 6658
rect 5509 6607 5521 6641
rect 5521 6607 5555 6641
rect 5555 6607 5561 6641
rect 5509 6606 5561 6607
rect 5443 6568 5495 6592
rect 5443 6540 5449 6568
rect 5449 6540 5483 6568
rect 5483 6540 5495 6568
rect 5509 6568 5561 6592
rect 5509 6540 5521 6568
rect 5521 6540 5555 6568
rect 5555 6540 5561 6568
rect 5443 6495 5495 6526
rect 5443 6474 5449 6495
rect 5449 6474 5483 6495
rect 5483 6474 5495 6495
rect 5509 6495 5561 6526
rect 5509 6474 5521 6495
rect 5521 6474 5555 6495
rect 5555 6474 5561 6495
rect 5443 6422 5495 6460
rect 5509 6422 5561 6460
rect 5443 6408 5449 6422
rect 5449 6408 5495 6422
rect 5509 6408 5555 6422
rect 5555 6408 5561 6422
rect 5443 6342 5449 6394
rect 5449 6342 5495 6394
rect 5509 6342 5555 6394
rect 5555 6342 5561 6394
rect 5443 6275 5449 6327
rect 5449 6275 5495 6327
rect 5509 6275 5555 6327
rect 5555 6275 5561 6327
rect 5443 6208 5449 6260
rect 5449 6208 5495 6260
rect 5509 6208 5555 6260
rect 5555 6208 5561 6260
rect 5720 13877 5772 13892
rect 5720 13843 5726 13877
rect 5726 13843 5760 13877
rect 5760 13843 5772 13877
rect 5720 13840 5772 13843
rect 5786 13877 5838 13892
rect 5786 13843 5798 13877
rect 5798 13843 5832 13877
rect 5832 13843 5838 13877
rect 5786 13840 5838 13843
rect 5720 13799 5772 13826
rect 5720 13774 5726 13799
rect 5726 13774 5760 13799
rect 5760 13774 5772 13799
rect 5786 13799 5838 13826
rect 5786 13774 5798 13799
rect 5798 13774 5832 13799
rect 5832 13774 5838 13799
rect 5720 13722 5772 13760
rect 5720 13708 5726 13722
rect 5726 13708 5760 13722
rect 5760 13708 5772 13722
rect 5786 13722 5838 13760
rect 5786 13708 5798 13722
rect 5798 13708 5832 13722
rect 5832 13708 5838 13722
rect 5720 13688 5726 13694
rect 5726 13688 5760 13694
rect 5760 13688 5772 13694
rect 5720 13645 5772 13688
rect 5720 13642 5726 13645
rect 5726 13642 5760 13645
rect 5760 13642 5772 13645
rect 5786 13688 5798 13694
rect 5798 13688 5832 13694
rect 5832 13688 5838 13694
rect 5786 13645 5838 13688
rect 5786 13642 5798 13645
rect 5798 13642 5832 13645
rect 5832 13642 5838 13645
rect 5720 13611 5726 13628
rect 5726 13611 5760 13628
rect 5760 13611 5772 13628
rect 5720 13576 5772 13611
rect 5786 13611 5798 13628
rect 5798 13611 5832 13628
rect 5832 13611 5838 13628
rect 5786 13576 5838 13611
rect 5720 13534 5726 13562
rect 5726 13534 5760 13562
rect 5760 13534 5772 13562
rect 5720 13510 5772 13534
rect 5786 13534 5798 13562
rect 5798 13534 5832 13562
rect 5832 13534 5838 13562
rect 5786 13510 5838 13534
rect 5720 13491 5772 13495
rect 5720 13457 5726 13491
rect 5726 13457 5760 13491
rect 5760 13457 5772 13491
rect 5720 13443 5772 13457
rect 5786 13491 5838 13495
rect 5786 13457 5798 13491
rect 5798 13457 5832 13491
rect 5832 13457 5838 13491
rect 5786 13443 5838 13457
rect 5720 13414 5772 13428
rect 5720 13380 5726 13414
rect 5726 13380 5760 13414
rect 5760 13380 5772 13414
rect 5720 13376 5772 13380
rect 5786 13414 5838 13428
rect 5786 13380 5798 13414
rect 5798 13380 5832 13414
rect 5832 13380 5838 13414
rect 5786 13376 5838 13380
rect 5720 11840 5726 11892
rect 5726 11840 5772 11892
rect 5786 11840 5832 11892
rect 5832 11840 5838 11892
rect 5720 11774 5726 11826
rect 5726 11774 5772 11826
rect 5786 11774 5832 11826
rect 5832 11774 5838 11826
rect 5720 11708 5726 11760
rect 5726 11708 5772 11760
rect 5786 11708 5832 11760
rect 5832 11708 5838 11760
rect 5720 11642 5726 11694
rect 5726 11642 5772 11694
rect 5786 11642 5832 11694
rect 5832 11642 5838 11694
rect 5720 11576 5726 11628
rect 5726 11576 5772 11628
rect 5786 11576 5832 11628
rect 5832 11576 5838 11628
rect 5720 11510 5726 11562
rect 5726 11510 5772 11562
rect 5786 11510 5832 11562
rect 5832 11510 5838 11562
rect 5720 11443 5726 11495
rect 5726 11443 5772 11495
rect 5786 11443 5832 11495
rect 5832 11443 5838 11495
rect 5720 11380 5726 11428
rect 5726 11380 5772 11428
rect 5786 11380 5832 11428
rect 5832 11380 5838 11428
rect 5720 11376 5772 11380
rect 5786 11376 5838 11380
rect 5720 9844 5726 9896
rect 5726 9844 5772 9896
rect 5786 9844 5832 9896
rect 5832 9844 5838 9896
rect 5720 9778 5726 9830
rect 5726 9778 5772 9830
rect 5786 9778 5832 9830
rect 5832 9778 5838 9830
rect 5720 9712 5726 9764
rect 5726 9712 5772 9764
rect 5786 9712 5832 9764
rect 5832 9712 5838 9764
rect 5720 9646 5726 9698
rect 5726 9646 5772 9698
rect 5786 9646 5832 9698
rect 5832 9646 5838 9698
rect 5720 9580 5726 9632
rect 5726 9580 5772 9632
rect 5786 9580 5832 9632
rect 5832 9580 5838 9632
rect 5720 9514 5726 9566
rect 5726 9514 5772 9566
rect 5786 9514 5832 9566
rect 5832 9514 5838 9566
rect 5720 9447 5726 9499
rect 5726 9447 5772 9499
rect 5786 9447 5832 9499
rect 5832 9447 5838 9499
rect 5720 9380 5726 9432
rect 5726 9380 5772 9432
rect 5786 9380 5832 9432
rect 5832 9380 5838 9432
rect 5720 7840 5726 7892
rect 5726 7840 5772 7892
rect 5786 7840 5832 7892
rect 5832 7840 5838 7892
rect 5720 7774 5726 7826
rect 5726 7774 5772 7826
rect 5786 7774 5832 7826
rect 5832 7774 5838 7826
rect 5720 7708 5726 7760
rect 5726 7708 5772 7760
rect 5786 7708 5832 7760
rect 5832 7708 5838 7760
rect 5720 7642 5726 7694
rect 5726 7642 5772 7694
rect 5786 7642 5832 7694
rect 5832 7642 5838 7694
rect 5720 7576 5726 7628
rect 5726 7576 5772 7628
rect 5786 7576 5832 7628
rect 5832 7576 5838 7628
rect 5720 7510 5726 7562
rect 5726 7510 5772 7562
rect 5786 7510 5832 7562
rect 5832 7510 5838 7562
rect 5720 7443 5726 7495
rect 5726 7443 5772 7495
rect 5786 7443 5832 7495
rect 5832 7443 5838 7495
rect 5720 7380 5726 7428
rect 5726 7380 5772 7428
rect 5786 7380 5832 7428
rect 5832 7380 5838 7428
rect 5720 7376 5772 7380
rect 5786 7376 5838 7380
rect 5720 5844 5726 5896
rect 5726 5844 5772 5896
rect 5786 5844 5832 5896
rect 5832 5844 5838 5896
rect 5720 5778 5726 5830
rect 5726 5778 5772 5830
rect 5786 5778 5832 5830
rect 5832 5778 5838 5830
rect 5720 5712 5726 5764
rect 5726 5712 5772 5764
rect 5786 5712 5832 5764
rect 5832 5712 5838 5764
rect 5720 5646 5726 5698
rect 5726 5646 5772 5698
rect 5786 5646 5832 5698
rect 5832 5646 5838 5698
rect 5720 5580 5726 5632
rect 5726 5580 5772 5632
rect 5786 5580 5832 5632
rect 5832 5580 5838 5632
rect 5720 5514 5726 5566
rect 5726 5514 5772 5566
rect 5786 5514 5832 5566
rect 5832 5514 5838 5566
rect 5720 5447 5726 5499
rect 5726 5447 5772 5499
rect 5786 5447 5832 5499
rect 5832 5447 5838 5499
rect 5720 5380 5726 5432
rect 5726 5380 5772 5432
rect 5786 5380 5832 5432
rect 5832 5380 5838 5432
rect 5997 14345 6049 14390
rect 5997 14338 6003 14345
rect 6003 14338 6037 14345
rect 6037 14338 6049 14345
rect 6063 14345 6115 14390
rect 6551 14668 6603 14720
rect 6617 14668 6669 14720
rect 6551 14602 6603 14654
rect 6617 14602 6669 14654
rect 6551 14536 6603 14588
rect 6617 14536 6669 14588
rect 6551 14470 6603 14522
rect 6617 14470 6669 14522
rect 6551 14404 6603 14456
rect 6617 14404 6669 14456
rect 6063 14338 6075 14345
rect 6075 14338 6109 14345
rect 6109 14338 6115 14345
rect 5997 14311 6003 14323
rect 6003 14311 6037 14323
rect 6037 14311 6049 14323
rect 5997 14271 6049 14311
rect 6063 14311 6075 14323
rect 6075 14311 6109 14323
rect 6109 14311 6115 14323
rect 6063 14271 6115 14311
rect 5997 14233 6003 14256
rect 6003 14233 6037 14256
rect 6037 14233 6049 14256
rect 5997 14204 6049 14233
rect 6063 14233 6075 14256
rect 6075 14233 6109 14256
rect 6109 14233 6115 14256
rect 6063 14204 6115 14233
rect 5997 12714 6049 12720
rect 5997 12680 6003 12714
rect 6003 12680 6037 12714
rect 6037 12680 6049 12714
rect 5997 12668 6049 12680
rect 6063 12714 6115 12720
rect 6063 12680 6075 12714
rect 6075 12680 6109 12714
rect 6109 12680 6115 12714
rect 6063 12668 6115 12680
rect 5997 12641 6049 12654
rect 5997 12607 6003 12641
rect 6003 12607 6037 12641
rect 6037 12607 6049 12641
rect 5997 12602 6049 12607
rect 6063 12641 6115 12654
rect 6063 12607 6075 12641
rect 6075 12607 6109 12641
rect 6109 12607 6115 12641
rect 6063 12602 6115 12607
rect 5997 12568 6049 12588
rect 5997 12536 6003 12568
rect 6003 12536 6037 12568
rect 6037 12536 6049 12568
rect 6063 12568 6115 12588
rect 6063 12536 6075 12568
rect 6075 12536 6109 12568
rect 6109 12536 6115 12568
rect 5997 12495 6049 12522
rect 5997 12470 6003 12495
rect 6003 12470 6037 12495
rect 6037 12470 6049 12495
rect 6063 12495 6115 12522
rect 6063 12470 6075 12495
rect 6075 12470 6109 12495
rect 6109 12470 6115 12495
rect 5997 12422 6049 12456
rect 6063 12422 6115 12456
rect 5997 12404 6003 12422
rect 6003 12404 6049 12422
rect 6063 12404 6109 12422
rect 6109 12404 6115 12422
rect 5997 12338 6003 12390
rect 6003 12338 6049 12390
rect 6063 12338 6109 12390
rect 6109 12338 6115 12390
rect 5997 12271 6003 12323
rect 6003 12271 6049 12323
rect 6063 12271 6109 12323
rect 6109 12271 6115 12323
rect 5997 12204 6003 12256
rect 6003 12204 6049 12256
rect 6063 12204 6109 12256
rect 6109 12204 6115 12256
rect 5997 10714 6049 10724
rect 5997 10680 6003 10714
rect 6003 10680 6037 10714
rect 6037 10680 6049 10714
rect 5997 10672 6049 10680
rect 6063 10714 6115 10724
rect 6063 10680 6075 10714
rect 6075 10680 6109 10714
rect 6109 10680 6115 10714
rect 6063 10672 6115 10680
rect 5997 10641 6049 10658
rect 5997 10607 6003 10641
rect 6003 10607 6037 10641
rect 6037 10607 6049 10641
rect 5997 10606 6049 10607
rect 6063 10641 6115 10658
rect 6063 10607 6075 10641
rect 6075 10607 6109 10641
rect 6109 10607 6115 10641
rect 6063 10606 6115 10607
rect 5997 10568 6049 10592
rect 5997 10540 6003 10568
rect 6003 10540 6037 10568
rect 6037 10540 6049 10568
rect 6063 10568 6115 10592
rect 6063 10540 6075 10568
rect 6075 10540 6109 10568
rect 6109 10540 6115 10568
rect 5997 10495 6049 10526
rect 5997 10474 6003 10495
rect 6003 10474 6037 10495
rect 6037 10474 6049 10495
rect 6063 10495 6115 10526
rect 6063 10474 6075 10495
rect 6075 10474 6109 10495
rect 6109 10474 6115 10495
rect 5997 10422 6049 10460
rect 6063 10422 6115 10460
rect 5997 10408 6003 10422
rect 6003 10408 6049 10422
rect 6063 10408 6109 10422
rect 6109 10408 6115 10422
rect 5997 10342 6003 10394
rect 6003 10342 6049 10394
rect 6063 10342 6109 10394
rect 6109 10342 6115 10394
rect 5997 10275 6003 10327
rect 6003 10275 6049 10327
rect 6063 10275 6109 10327
rect 6109 10275 6115 10327
rect 5997 10208 6003 10260
rect 6003 10208 6049 10260
rect 6063 10208 6109 10260
rect 6109 10208 6115 10260
rect 5997 8714 6049 8720
rect 5997 8680 6003 8714
rect 6003 8680 6037 8714
rect 6037 8680 6049 8714
rect 5997 8668 6049 8680
rect 6063 8714 6115 8720
rect 6063 8680 6075 8714
rect 6075 8680 6109 8714
rect 6109 8680 6115 8714
rect 6063 8668 6115 8680
rect 5997 8641 6049 8654
rect 5997 8607 6003 8641
rect 6003 8607 6037 8641
rect 6037 8607 6049 8641
rect 5997 8602 6049 8607
rect 6063 8641 6115 8654
rect 6063 8607 6075 8641
rect 6075 8607 6109 8641
rect 6109 8607 6115 8641
rect 6063 8602 6115 8607
rect 5997 8568 6049 8588
rect 5997 8536 6003 8568
rect 6003 8536 6037 8568
rect 6037 8536 6049 8568
rect 6063 8568 6115 8588
rect 6063 8536 6075 8568
rect 6075 8536 6109 8568
rect 6109 8536 6115 8568
rect 5997 8495 6049 8522
rect 5997 8470 6003 8495
rect 6003 8470 6037 8495
rect 6037 8470 6049 8495
rect 6063 8495 6115 8522
rect 6063 8470 6075 8495
rect 6075 8470 6109 8495
rect 6109 8470 6115 8495
rect 5997 8422 6049 8456
rect 6063 8422 6115 8456
rect 5997 8404 6003 8422
rect 6003 8404 6049 8422
rect 6063 8404 6109 8422
rect 6109 8404 6115 8422
rect 5997 8338 6003 8390
rect 6003 8338 6049 8390
rect 6063 8338 6109 8390
rect 6109 8338 6115 8390
rect 5997 8271 6003 8323
rect 6003 8271 6049 8323
rect 6063 8271 6109 8323
rect 6109 8271 6115 8323
rect 5997 8204 6003 8256
rect 6003 8204 6049 8256
rect 6063 8204 6109 8256
rect 6109 8204 6115 8256
rect 5997 6714 6049 6724
rect 5997 6680 6003 6714
rect 6003 6680 6037 6714
rect 6037 6680 6049 6714
rect 5997 6672 6049 6680
rect 6063 6714 6115 6724
rect 6063 6680 6075 6714
rect 6075 6680 6109 6714
rect 6109 6680 6115 6714
rect 6063 6672 6115 6680
rect 5997 6641 6049 6658
rect 5997 6607 6003 6641
rect 6003 6607 6037 6641
rect 6037 6607 6049 6641
rect 5997 6606 6049 6607
rect 6063 6641 6115 6658
rect 6063 6607 6075 6641
rect 6075 6607 6109 6641
rect 6109 6607 6115 6641
rect 6063 6606 6115 6607
rect 5997 6568 6049 6592
rect 5997 6540 6003 6568
rect 6003 6540 6037 6568
rect 6037 6540 6049 6568
rect 6063 6568 6115 6592
rect 6063 6540 6075 6568
rect 6075 6540 6109 6568
rect 6109 6540 6115 6568
rect 5997 6495 6049 6526
rect 5997 6474 6003 6495
rect 6003 6474 6037 6495
rect 6037 6474 6049 6495
rect 6063 6495 6115 6526
rect 6063 6474 6075 6495
rect 6075 6474 6109 6495
rect 6109 6474 6115 6495
rect 5997 6422 6049 6460
rect 6063 6422 6115 6460
rect 5997 6408 6003 6422
rect 6003 6408 6049 6422
rect 6063 6408 6109 6422
rect 6109 6408 6115 6422
rect 5997 6342 6003 6394
rect 6003 6342 6049 6394
rect 6063 6342 6109 6394
rect 6109 6342 6115 6394
rect 5997 6275 6003 6327
rect 6003 6275 6049 6327
rect 6063 6275 6109 6327
rect 6109 6275 6115 6327
rect 5997 6208 6003 6260
rect 6003 6208 6049 6260
rect 6063 6208 6109 6260
rect 6109 6208 6115 6260
rect 6274 13877 6326 13892
rect 6274 13843 6280 13877
rect 6280 13843 6314 13877
rect 6314 13843 6326 13877
rect 6274 13840 6326 13843
rect 6340 13877 6392 13892
rect 6340 13843 6352 13877
rect 6352 13843 6386 13877
rect 6386 13843 6392 13877
rect 6340 13840 6392 13843
rect 6274 13799 6326 13826
rect 6274 13774 6280 13799
rect 6280 13774 6314 13799
rect 6314 13774 6326 13799
rect 6340 13799 6392 13826
rect 6340 13774 6352 13799
rect 6352 13774 6386 13799
rect 6386 13774 6392 13799
rect 6274 13722 6326 13760
rect 6274 13708 6280 13722
rect 6280 13708 6314 13722
rect 6314 13708 6326 13722
rect 6340 13722 6392 13760
rect 6340 13708 6352 13722
rect 6352 13708 6386 13722
rect 6386 13708 6392 13722
rect 6274 13688 6280 13694
rect 6280 13688 6314 13694
rect 6314 13688 6326 13694
rect 6274 13645 6326 13688
rect 6274 13642 6280 13645
rect 6280 13642 6314 13645
rect 6314 13642 6326 13645
rect 6340 13688 6352 13694
rect 6352 13688 6386 13694
rect 6386 13688 6392 13694
rect 6340 13645 6392 13688
rect 6340 13642 6352 13645
rect 6352 13642 6386 13645
rect 6386 13642 6392 13645
rect 6274 13611 6280 13628
rect 6280 13611 6314 13628
rect 6314 13611 6326 13628
rect 6274 13576 6326 13611
rect 6340 13611 6352 13628
rect 6352 13611 6386 13628
rect 6386 13611 6392 13628
rect 6340 13576 6392 13611
rect 6274 13534 6280 13562
rect 6280 13534 6314 13562
rect 6314 13534 6326 13562
rect 6274 13510 6326 13534
rect 6340 13534 6352 13562
rect 6352 13534 6386 13562
rect 6386 13534 6392 13562
rect 6340 13510 6392 13534
rect 6274 13491 6326 13495
rect 6274 13457 6280 13491
rect 6280 13457 6314 13491
rect 6314 13457 6326 13491
rect 6274 13443 6326 13457
rect 6340 13491 6392 13495
rect 6340 13457 6352 13491
rect 6352 13457 6386 13491
rect 6386 13457 6392 13491
rect 6340 13443 6392 13457
rect 6274 13414 6326 13428
rect 6274 13380 6280 13414
rect 6280 13380 6314 13414
rect 6314 13380 6326 13414
rect 6274 13376 6326 13380
rect 6340 13414 6392 13428
rect 6340 13380 6352 13414
rect 6352 13380 6386 13414
rect 6386 13380 6392 13414
rect 6340 13376 6392 13380
rect 6274 11840 6280 11892
rect 6280 11840 6326 11892
rect 6340 11840 6386 11892
rect 6386 11840 6392 11892
rect 6274 11774 6280 11826
rect 6280 11774 6326 11826
rect 6340 11774 6386 11826
rect 6386 11774 6392 11826
rect 6274 11708 6280 11760
rect 6280 11708 6326 11760
rect 6340 11708 6386 11760
rect 6386 11708 6392 11760
rect 6274 11642 6280 11694
rect 6280 11642 6326 11694
rect 6340 11642 6386 11694
rect 6386 11642 6392 11694
rect 6274 11576 6280 11628
rect 6280 11576 6326 11628
rect 6340 11576 6386 11628
rect 6386 11576 6392 11628
rect 6274 11510 6280 11562
rect 6280 11510 6326 11562
rect 6340 11510 6386 11562
rect 6386 11510 6392 11562
rect 6274 11443 6280 11495
rect 6280 11443 6326 11495
rect 6340 11443 6386 11495
rect 6386 11443 6392 11495
rect 6274 11380 6280 11428
rect 6280 11380 6326 11428
rect 6340 11380 6386 11428
rect 6386 11380 6392 11428
rect 6274 11376 6326 11380
rect 6340 11376 6392 11380
rect 6274 9844 6280 9896
rect 6280 9844 6326 9896
rect 6340 9844 6386 9896
rect 6386 9844 6392 9896
rect 6274 9778 6280 9830
rect 6280 9778 6326 9830
rect 6340 9778 6386 9830
rect 6386 9778 6392 9830
rect 6274 9712 6280 9764
rect 6280 9712 6326 9764
rect 6340 9712 6386 9764
rect 6386 9712 6392 9764
rect 6274 9646 6280 9698
rect 6280 9646 6326 9698
rect 6340 9646 6386 9698
rect 6386 9646 6392 9698
rect 6274 9580 6280 9632
rect 6280 9580 6326 9632
rect 6340 9580 6386 9632
rect 6386 9580 6392 9632
rect 6274 9514 6280 9566
rect 6280 9514 6326 9566
rect 6340 9514 6386 9566
rect 6386 9514 6392 9566
rect 6274 9447 6280 9499
rect 6280 9447 6326 9499
rect 6340 9447 6386 9499
rect 6386 9447 6392 9499
rect 6274 9380 6280 9432
rect 6280 9380 6326 9432
rect 6340 9380 6386 9432
rect 6386 9380 6392 9432
rect 6274 7840 6280 7892
rect 6280 7840 6326 7892
rect 6340 7840 6386 7892
rect 6386 7840 6392 7892
rect 6274 7774 6280 7826
rect 6280 7774 6326 7826
rect 6340 7774 6386 7826
rect 6386 7774 6392 7826
rect 6274 7708 6280 7760
rect 6280 7708 6326 7760
rect 6340 7708 6386 7760
rect 6386 7708 6392 7760
rect 6274 7642 6280 7694
rect 6280 7642 6326 7694
rect 6340 7642 6386 7694
rect 6386 7642 6392 7694
rect 6274 7576 6280 7628
rect 6280 7576 6326 7628
rect 6340 7576 6386 7628
rect 6386 7576 6392 7628
rect 6274 7510 6280 7562
rect 6280 7510 6326 7562
rect 6340 7510 6386 7562
rect 6386 7510 6392 7562
rect 6274 7443 6280 7495
rect 6280 7443 6326 7495
rect 6340 7443 6386 7495
rect 6386 7443 6392 7495
rect 6274 7380 6280 7428
rect 6280 7380 6326 7428
rect 6340 7380 6386 7428
rect 6386 7380 6392 7428
rect 6274 7376 6326 7380
rect 6340 7376 6392 7380
rect 6274 5844 6280 5896
rect 6280 5844 6326 5896
rect 6340 5844 6386 5896
rect 6386 5844 6392 5896
rect 6274 5778 6280 5830
rect 6280 5778 6326 5830
rect 6340 5778 6386 5830
rect 6386 5778 6392 5830
rect 6274 5712 6280 5764
rect 6280 5712 6326 5764
rect 6340 5712 6386 5764
rect 6386 5712 6392 5764
rect 6274 5646 6280 5698
rect 6280 5646 6326 5698
rect 6340 5646 6386 5698
rect 6386 5646 6392 5698
rect 6274 5580 6280 5632
rect 6280 5580 6326 5632
rect 6340 5580 6386 5632
rect 6386 5580 6392 5632
rect 6274 5514 6280 5566
rect 6280 5514 6326 5566
rect 6340 5514 6386 5566
rect 6386 5514 6392 5566
rect 6274 5447 6280 5499
rect 6280 5447 6326 5499
rect 6340 5447 6386 5499
rect 6386 5447 6392 5499
rect 6274 5380 6280 5432
rect 6280 5380 6326 5432
rect 6340 5380 6386 5432
rect 6386 5380 6392 5432
rect 6551 14345 6603 14390
rect 6551 14338 6557 14345
rect 6557 14338 6591 14345
rect 6591 14338 6603 14345
rect 6617 14345 6669 14390
rect 7105 14668 7157 14720
rect 7171 14668 7223 14720
rect 7105 14602 7157 14654
rect 7171 14602 7223 14654
rect 7105 14536 7157 14588
rect 7171 14536 7223 14588
rect 7105 14470 7157 14522
rect 7171 14470 7223 14522
rect 7105 14404 7157 14456
rect 7171 14404 7223 14456
rect 6617 14338 6629 14345
rect 6629 14338 6663 14345
rect 6663 14338 6669 14345
rect 6551 14311 6557 14323
rect 6557 14311 6591 14323
rect 6591 14311 6603 14323
rect 6551 14271 6603 14311
rect 6617 14311 6629 14323
rect 6629 14311 6663 14323
rect 6663 14311 6669 14323
rect 6617 14271 6669 14311
rect 6551 14233 6557 14256
rect 6557 14233 6591 14256
rect 6591 14233 6603 14256
rect 6551 14204 6603 14233
rect 6617 14233 6629 14256
rect 6629 14233 6663 14256
rect 6663 14233 6669 14256
rect 6617 14204 6669 14233
rect 6551 12714 6603 12720
rect 6551 12680 6557 12714
rect 6557 12680 6591 12714
rect 6591 12680 6603 12714
rect 6551 12668 6603 12680
rect 6617 12714 6669 12720
rect 6617 12680 6629 12714
rect 6629 12680 6663 12714
rect 6663 12680 6669 12714
rect 6617 12668 6669 12680
rect 6551 12641 6603 12654
rect 6551 12607 6557 12641
rect 6557 12607 6591 12641
rect 6591 12607 6603 12641
rect 6551 12602 6603 12607
rect 6617 12641 6669 12654
rect 6617 12607 6629 12641
rect 6629 12607 6663 12641
rect 6663 12607 6669 12641
rect 6617 12602 6669 12607
rect 6551 12568 6603 12588
rect 6551 12536 6557 12568
rect 6557 12536 6591 12568
rect 6591 12536 6603 12568
rect 6617 12568 6669 12588
rect 6617 12536 6629 12568
rect 6629 12536 6663 12568
rect 6663 12536 6669 12568
rect 6551 12495 6603 12522
rect 6551 12470 6557 12495
rect 6557 12470 6591 12495
rect 6591 12470 6603 12495
rect 6617 12495 6669 12522
rect 6617 12470 6629 12495
rect 6629 12470 6663 12495
rect 6663 12470 6669 12495
rect 6551 12422 6603 12456
rect 6617 12422 6669 12456
rect 6551 12404 6557 12422
rect 6557 12404 6603 12422
rect 6617 12404 6663 12422
rect 6663 12404 6669 12422
rect 6551 12338 6557 12390
rect 6557 12338 6603 12390
rect 6617 12338 6663 12390
rect 6663 12338 6669 12390
rect 6551 12271 6557 12323
rect 6557 12271 6603 12323
rect 6617 12271 6663 12323
rect 6663 12271 6669 12323
rect 6551 12204 6557 12256
rect 6557 12204 6603 12256
rect 6617 12204 6663 12256
rect 6663 12204 6669 12256
rect 6551 10714 6603 10724
rect 6551 10680 6557 10714
rect 6557 10680 6591 10714
rect 6591 10680 6603 10714
rect 6551 10672 6603 10680
rect 6617 10714 6669 10724
rect 6617 10680 6629 10714
rect 6629 10680 6663 10714
rect 6663 10680 6669 10714
rect 6617 10672 6669 10680
rect 6551 10641 6603 10658
rect 6551 10607 6557 10641
rect 6557 10607 6591 10641
rect 6591 10607 6603 10641
rect 6551 10606 6603 10607
rect 6617 10641 6669 10658
rect 6617 10607 6629 10641
rect 6629 10607 6663 10641
rect 6663 10607 6669 10641
rect 6617 10606 6669 10607
rect 6551 10568 6603 10592
rect 6551 10540 6557 10568
rect 6557 10540 6591 10568
rect 6591 10540 6603 10568
rect 6617 10568 6669 10592
rect 6617 10540 6629 10568
rect 6629 10540 6663 10568
rect 6663 10540 6669 10568
rect 6551 10495 6603 10526
rect 6551 10474 6557 10495
rect 6557 10474 6591 10495
rect 6591 10474 6603 10495
rect 6617 10495 6669 10526
rect 6617 10474 6629 10495
rect 6629 10474 6663 10495
rect 6663 10474 6669 10495
rect 6551 10422 6603 10460
rect 6617 10422 6669 10460
rect 6551 10408 6557 10422
rect 6557 10408 6603 10422
rect 6617 10408 6663 10422
rect 6663 10408 6669 10422
rect 6551 10342 6557 10394
rect 6557 10342 6603 10394
rect 6617 10342 6663 10394
rect 6663 10342 6669 10394
rect 6551 10275 6557 10327
rect 6557 10275 6603 10327
rect 6617 10275 6663 10327
rect 6663 10275 6669 10327
rect 6551 10208 6557 10260
rect 6557 10208 6603 10260
rect 6617 10208 6663 10260
rect 6663 10208 6669 10260
rect 6551 8714 6603 8720
rect 6551 8680 6557 8714
rect 6557 8680 6591 8714
rect 6591 8680 6603 8714
rect 6551 8668 6603 8680
rect 6617 8714 6669 8720
rect 6617 8680 6629 8714
rect 6629 8680 6663 8714
rect 6663 8680 6669 8714
rect 6617 8668 6669 8680
rect 6551 8641 6603 8654
rect 6551 8607 6557 8641
rect 6557 8607 6591 8641
rect 6591 8607 6603 8641
rect 6551 8602 6603 8607
rect 6617 8641 6669 8654
rect 6617 8607 6629 8641
rect 6629 8607 6663 8641
rect 6663 8607 6669 8641
rect 6617 8602 6669 8607
rect 6551 8568 6603 8588
rect 6551 8536 6557 8568
rect 6557 8536 6591 8568
rect 6591 8536 6603 8568
rect 6617 8568 6669 8588
rect 6617 8536 6629 8568
rect 6629 8536 6663 8568
rect 6663 8536 6669 8568
rect 6551 8495 6603 8522
rect 6551 8470 6557 8495
rect 6557 8470 6591 8495
rect 6591 8470 6603 8495
rect 6617 8495 6669 8522
rect 6617 8470 6629 8495
rect 6629 8470 6663 8495
rect 6663 8470 6669 8495
rect 6551 8422 6603 8456
rect 6617 8422 6669 8456
rect 6551 8404 6557 8422
rect 6557 8404 6603 8422
rect 6617 8404 6663 8422
rect 6663 8404 6669 8422
rect 6551 8338 6557 8390
rect 6557 8338 6603 8390
rect 6617 8338 6663 8390
rect 6663 8338 6669 8390
rect 6551 8271 6557 8323
rect 6557 8271 6603 8323
rect 6617 8271 6663 8323
rect 6663 8271 6669 8323
rect 6551 8204 6557 8256
rect 6557 8204 6603 8256
rect 6617 8204 6663 8256
rect 6663 8204 6669 8256
rect 6551 6714 6603 6724
rect 6551 6680 6557 6714
rect 6557 6680 6591 6714
rect 6591 6680 6603 6714
rect 6551 6672 6603 6680
rect 6617 6714 6669 6724
rect 6617 6680 6629 6714
rect 6629 6680 6663 6714
rect 6663 6680 6669 6714
rect 6617 6672 6669 6680
rect 6551 6641 6603 6658
rect 6551 6607 6557 6641
rect 6557 6607 6591 6641
rect 6591 6607 6603 6641
rect 6551 6606 6603 6607
rect 6617 6641 6669 6658
rect 6617 6607 6629 6641
rect 6629 6607 6663 6641
rect 6663 6607 6669 6641
rect 6617 6606 6669 6607
rect 6551 6568 6603 6592
rect 6551 6540 6557 6568
rect 6557 6540 6591 6568
rect 6591 6540 6603 6568
rect 6617 6568 6669 6592
rect 6617 6540 6629 6568
rect 6629 6540 6663 6568
rect 6663 6540 6669 6568
rect 6551 6495 6603 6526
rect 6551 6474 6557 6495
rect 6557 6474 6591 6495
rect 6591 6474 6603 6495
rect 6617 6495 6669 6526
rect 6617 6474 6629 6495
rect 6629 6474 6663 6495
rect 6663 6474 6669 6495
rect 6551 6422 6603 6460
rect 6617 6422 6669 6460
rect 6551 6408 6557 6422
rect 6557 6408 6603 6422
rect 6617 6408 6663 6422
rect 6663 6408 6669 6422
rect 6551 6342 6557 6394
rect 6557 6342 6603 6394
rect 6617 6342 6663 6394
rect 6663 6342 6669 6394
rect 6551 6275 6557 6327
rect 6557 6275 6603 6327
rect 6617 6275 6663 6327
rect 6663 6275 6669 6327
rect 6551 6208 6557 6260
rect 6557 6208 6603 6260
rect 6617 6208 6663 6260
rect 6663 6208 6669 6260
rect 6828 13877 6880 13892
rect 6828 13843 6834 13877
rect 6834 13843 6868 13877
rect 6868 13843 6880 13877
rect 6828 13840 6880 13843
rect 6894 13877 6946 13892
rect 6894 13843 6906 13877
rect 6906 13843 6940 13877
rect 6940 13843 6946 13877
rect 6894 13840 6946 13843
rect 6828 13799 6880 13826
rect 6828 13774 6834 13799
rect 6834 13774 6868 13799
rect 6868 13774 6880 13799
rect 6894 13799 6946 13826
rect 6894 13774 6906 13799
rect 6906 13774 6940 13799
rect 6940 13774 6946 13799
rect 6828 13722 6880 13760
rect 6828 13708 6834 13722
rect 6834 13708 6868 13722
rect 6868 13708 6880 13722
rect 6894 13722 6946 13760
rect 6894 13708 6906 13722
rect 6906 13708 6940 13722
rect 6940 13708 6946 13722
rect 6828 13688 6834 13694
rect 6834 13688 6868 13694
rect 6868 13688 6880 13694
rect 6828 13645 6880 13688
rect 6828 13642 6834 13645
rect 6834 13642 6868 13645
rect 6868 13642 6880 13645
rect 6894 13688 6906 13694
rect 6906 13688 6940 13694
rect 6940 13688 6946 13694
rect 6894 13645 6946 13688
rect 6894 13642 6906 13645
rect 6906 13642 6940 13645
rect 6940 13642 6946 13645
rect 6828 13611 6834 13628
rect 6834 13611 6868 13628
rect 6868 13611 6880 13628
rect 6828 13576 6880 13611
rect 6894 13611 6906 13628
rect 6906 13611 6940 13628
rect 6940 13611 6946 13628
rect 6894 13576 6946 13611
rect 6828 13534 6834 13562
rect 6834 13534 6868 13562
rect 6868 13534 6880 13562
rect 6828 13510 6880 13534
rect 6894 13534 6906 13562
rect 6906 13534 6940 13562
rect 6940 13534 6946 13562
rect 6894 13510 6946 13534
rect 6828 13491 6880 13495
rect 6828 13457 6834 13491
rect 6834 13457 6868 13491
rect 6868 13457 6880 13491
rect 6828 13443 6880 13457
rect 6894 13491 6946 13495
rect 6894 13457 6906 13491
rect 6906 13457 6940 13491
rect 6940 13457 6946 13491
rect 6894 13443 6946 13457
rect 6828 13414 6880 13428
rect 6828 13380 6834 13414
rect 6834 13380 6868 13414
rect 6868 13380 6880 13414
rect 6828 13376 6880 13380
rect 6894 13414 6946 13428
rect 6894 13380 6906 13414
rect 6906 13380 6940 13414
rect 6940 13380 6946 13414
rect 6894 13376 6946 13380
rect 6828 11840 6834 11892
rect 6834 11840 6880 11892
rect 6894 11840 6940 11892
rect 6940 11840 6946 11892
rect 6828 11774 6834 11826
rect 6834 11774 6880 11826
rect 6894 11774 6940 11826
rect 6940 11774 6946 11826
rect 6828 11708 6834 11760
rect 6834 11708 6880 11760
rect 6894 11708 6940 11760
rect 6940 11708 6946 11760
rect 6828 11642 6834 11694
rect 6834 11642 6880 11694
rect 6894 11642 6940 11694
rect 6940 11642 6946 11694
rect 6828 11576 6834 11628
rect 6834 11576 6880 11628
rect 6894 11576 6940 11628
rect 6940 11576 6946 11628
rect 6828 11510 6834 11562
rect 6834 11510 6880 11562
rect 6894 11510 6940 11562
rect 6940 11510 6946 11562
rect 6828 11443 6834 11495
rect 6834 11443 6880 11495
rect 6894 11443 6940 11495
rect 6940 11443 6946 11495
rect 6828 11380 6834 11428
rect 6834 11380 6880 11428
rect 6894 11380 6940 11428
rect 6940 11380 6946 11428
rect 6828 11376 6880 11380
rect 6894 11376 6946 11380
rect 6828 9844 6834 9896
rect 6834 9844 6880 9896
rect 6894 9844 6940 9896
rect 6940 9844 6946 9896
rect 6828 9778 6834 9830
rect 6834 9778 6880 9830
rect 6894 9778 6940 9830
rect 6940 9778 6946 9830
rect 6828 9712 6834 9764
rect 6834 9712 6880 9764
rect 6894 9712 6940 9764
rect 6940 9712 6946 9764
rect 6828 9646 6834 9698
rect 6834 9646 6880 9698
rect 6894 9646 6940 9698
rect 6940 9646 6946 9698
rect 6828 9580 6834 9632
rect 6834 9580 6880 9632
rect 6894 9580 6940 9632
rect 6940 9580 6946 9632
rect 6828 9514 6834 9566
rect 6834 9514 6880 9566
rect 6894 9514 6940 9566
rect 6940 9514 6946 9566
rect 6828 9447 6834 9499
rect 6834 9447 6880 9499
rect 6894 9447 6940 9499
rect 6940 9447 6946 9499
rect 6828 9380 6834 9432
rect 6834 9380 6880 9432
rect 6894 9380 6940 9432
rect 6940 9380 6946 9432
rect 6828 7840 6834 7892
rect 6834 7840 6880 7892
rect 6894 7840 6940 7892
rect 6940 7840 6946 7892
rect 6828 7774 6834 7826
rect 6834 7774 6880 7826
rect 6894 7774 6940 7826
rect 6940 7774 6946 7826
rect 6828 7708 6834 7760
rect 6834 7708 6880 7760
rect 6894 7708 6940 7760
rect 6940 7708 6946 7760
rect 6828 7642 6834 7694
rect 6834 7642 6880 7694
rect 6894 7642 6940 7694
rect 6940 7642 6946 7694
rect 6828 7576 6834 7628
rect 6834 7576 6880 7628
rect 6894 7576 6940 7628
rect 6940 7576 6946 7628
rect 6828 7510 6834 7562
rect 6834 7510 6880 7562
rect 6894 7510 6940 7562
rect 6940 7510 6946 7562
rect 6828 7443 6834 7495
rect 6834 7443 6880 7495
rect 6894 7443 6940 7495
rect 6940 7443 6946 7495
rect 6828 7380 6834 7428
rect 6834 7380 6880 7428
rect 6894 7380 6940 7428
rect 6940 7380 6946 7428
rect 6828 7376 6880 7380
rect 6894 7376 6946 7380
rect 6828 5844 6834 5896
rect 6834 5844 6880 5896
rect 6894 5844 6940 5896
rect 6940 5844 6946 5896
rect 6828 5778 6834 5830
rect 6834 5778 6880 5830
rect 6894 5778 6940 5830
rect 6940 5778 6946 5830
rect 6828 5712 6834 5764
rect 6834 5712 6880 5764
rect 6894 5712 6940 5764
rect 6940 5712 6946 5764
rect 6828 5646 6834 5698
rect 6834 5646 6880 5698
rect 6894 5646 6940 5698
rect 6940 5646 6946 5698
rect 6828 5580 6834 5632
rect 6834 5580 6880 5632
rect 6894 5580 6940 5632
rect 6940 5580 6946 5632
rect 6828 5514 6834 5566
rect 6834 5514 6880 5566
rect 6894 5514 6940 5566
rect 6940 5514 6946 5566
rect 6828 5447 6834 5499
rect 6834 5447 6880 5499
rect 6894 5447 6940 5499
rect 6940 5447 6946 5499
rect 6828 5380 6834 5432
rect 6834 5380 6880 5432
rect 6894 5380 6940 5432
rect 6940 5380 6946 5432
rect 7105 14345 7157 14390
rect 7105 14338 7111 14345
rect 7111 14338 7145 14345
rect 7145 14338 7157 14345
rect 7171 14345 7223 14390
rect 7659 14668 7711 14720
rect 7725 14668 7777 14720
rect 7659 14602 7711 14654
rect 7725 14602 7777 14654
rect 7659 14536 7711 14588
rect 7725 14536 7777 14588
rect 7659 14470 7711 14522
rect 7725 14470 7777 14522
rect 7659 14404 7711 14456
rect 7725 14404 7777 14456
rect 7171 14338 7183 14345
rect 7183 14338 7217 14345
rect 7217 14338 7223 14345
rect 7105 14311 7111 14323
rect 7111 14311 7145 14323
rect 7145 14311 7157 14323
rect 7105 14271 7157 14311
rect 7171 14311 7183 14323
rect 7183 14311 7217 14323
rect 7217 14311 7223 14323
rect 7171 14271 7223 14311
rect 7105 14233 7111 14256
rect 7111 14233 7145 14256
rect 7145 14233 7157 14256
rect 7105 14204 7157 14233
rect 7171 14233 7183 14256
rect 7183 14233 7217 14256
rect 7217 14233 7223 14256
rect 7171 14204 7223 14233
rect 7105 12714 7157 12720
rect 7105 12680 7111 12714
rect 7111 12680 7145 12714
rect 7145 12680 7157 12714
rect 7105 12668 7157 12680
rect 7171 12714 7223 12720
rect 7171 12680 7183 12714
rect 7183 12680 7217 12714
rect 7217 12680 7223 12714
rect 7171 12668 7223 12680
rect 7105 12641 7157 12654
rect 7105 12607 7111 12641
rect 7111 12607 7145 12641
rect 7145 12607 7157 12641
rect 7105 12602 7157 12607
rect 7171 12641 7223 12654
rect 7171 12607 7183 12641
rect 7183 12607 7217 12641
rect 7217 12607 7223 12641
rect 7171 12602 7223 12607
rect 7105 12568 7157 12588
rect 7105 12536 7111 12568
rect 7111 12536 7145 12568
rect 7145 12536 7157 12568
rect 7171 12568 7223 12588
rect 7171 12536 7183 12568
rect 7183 12536 7217 12568
rect 7217 12536 7223 12568
rect 7105 12495 7157 12522
rect 7105 12470 7111 12495
rect 7111 12470 7145 12495
rect 7145 12470 7157 12495
rect 7171 12495 7223 12522
rect 7171 12470 7183 12495
rect 7183 12470 7217 12495
rect 7217 12470 7223 12495
rect 7105 12422 7157 12456
rect 7171 12422 7223 12456
rect 7105 12404 7111 12422
rect 7111 12404 7157 12422
rect 7171 12404 7217 12422
rect 7217 12404 7223 12422
rect 7105 12338 7111 12390
rect 7111 12338 7157 12390
rect 7171 12338 7217 12390
rect 7217 12338 7223 12390
rect 7105 12271 7111 12323
rect 7111 12271 7157 12323
rect 7171 12271 7217 12323
rect 7217 12271 7223 12323
rect 7105 12204 7111 12256
rect 7111 12204 7157 12256
rect 7171 12204 7217 12256
rect 7217 12204 7223 12256
rect 7105 10714 7157 10724
rect 7105 10680 7111 10714
rect 7111 10680 7145 10714
rect 7145 10680 7157 10714
rect 7105 10672 7157 10680
rect 7171 10714 7223 10724
rect 7171 10680 7183 10714
rect 7183 10680 7217 10714
rect 7217 10680 7223 10714
rect 7171 10672 7223 10680
rect 7105 10641 7157 10658
rect 7105 10607 7111 10641
rect 7111 10607 7145 10641
rect 7145 10607 7157 10641
rect 7105 10606 7157 10607
rect 7171 10641 7223 10658
rect 7171 10607 7183 10641
rect 7183 10607 7217 10641
rect 7217 10607 7223 10641
rect 7171 10606 7223 10607
rect 7105 10568 7157 10592
rect 7105 10540 7111 10568
rect 7111 10540 7145 10568
rect 7145 10540 7157 10568
rect 7171 10568 7223 10592
rect 7171 10540 7183 10568
rect 7183 10540 7217 10568
rect 7217 10540 7223 10568
rect 7105 10495 7157 10526
rect 7105 10474 7111 10495
rect 7111 10474 7145 10495
rect 7145 10474 7157 10495
rect 7171 10495 7223 10526
rect 7171 10474 7183 10495
rect 7183 10474 7217 10495
rect 7217 10474 7223 10495
rect 7105 10422 7157 10460
rect 7171 10422 7223 10460
rect 7105 10408 7111 10422
rect 7111 10408 7157 10422
rect 7171 10408 7217 10422
rect 7217 10408 7223 10422
rect 7105 10342 7111 10394
rect 7111 10342 7157 10394
rect 7171 10342 7217 10394
rect 7217 10342 7223 10394
rect 7105 10275 7111 10327
rect 7111 10275 7157 10327
rect 7171 10275 7217 10327
rect 7217 10275 7223 10327
rect 7105 10208 7111 10260
rect 7111 10208 7157 10260
rect 7171 10208 7217 10260
rect 7217 10208 7223 10260
rect 7105 8714 7157 8720
rect 7105 8680 7111 8714
rect 7111 8680 7145 8714
rect 7145 8680 7157 8714
rect 7105 8668 7157 8680
rect 7171 8714 7223 8720
rect 7171 8680 7183 8714
rect 7183 8680 7217 8714
rect 7217 8680 7223 8714
rect 7171 8668 7223 8680
rect 7105 8641 7157 8654
rect 7105 8607 7111 8641
rect 7111 8607 7145 8641
rect 7145 8607 7157 8641
rect 7105 8602 7157 8607
rect 7171 8641 7223 8654
rect 7171 8607 7183 8641
rect 7183 8607 7217 8641
rect 7217 8607 7223 8641
rect 7171 8602 7223 8607
rect 7105 8568 7157 8588
rect 7105 8536 7111 8568
rect 7111 8536 7145 8568
rect 7145 8536 7157 8568
rect 7171 8568 7223 8588
rect 7171 8536 7183 8568
rect 7183 8536 7217 8568
rect 7217 8536 7223 8568
rect 7105 8495 7157 8522
rect 7105 8470 7111 8495
rect 7111 8470 7145 8495
rect 7145 8470 7157 8495
rect 7171 8495 7223 8522
rect 7171 8470 7183 8495
rect 7183 8470 7217 8495
rect 7217 8470 7223 8495
rect 7105 8422 7157 8456
rect 7171 8422 7223 8456
rect 7105 8404 7111 8422
rect 7111 8404 7157 8422
rect 7171 8404 7217 8422
rect 7217 8404 7223 8422
rect 7105 8338 7111 8390
rect 7111 8338 7157 8390
rect 7171 8338 7217 8390
rect 7217 8338 7223 8390
rect 7105 8271 7111 8323
rect 7111 8271 7157 8323
rect 7171 8271 7217 8323
rect 7217 8271 7223 8323
rect 7105 8204 7111 8256
rect 7111 8204 7157 8256
rect 7171 8204 7217 8256
rect 7217 8204 7223 8256
rect 7105 6714 7157 6724
rect 7105 6680 7111 6714
rect 7111 6680 7145 6714
rect 7145 6680 7157 6714
rect 7105 6672 7157 6680
rect 7171 6714 7223 6724
rect 7171 6680 7183 6714
rect 7183 6680 7217 6714
rect 7217 6680 7223 6714
rect 7171 6672 7223 6680
rect 7105 6641 7157 6658
rect 7105 6607 7111 6641
rect 7111 6607 7145 6641
rect 7145 6607 7157 6641
rect 7105 6606 7157 6607
rect 7171 6641 7223 6658
rect 7171 6607 7183 6641
rect 7183 6607 7217 6641
rect 7217 6607 7223 6641
rect 7171 6606 7223 6607
rect 7105 6568 7157 6592
rect 7105 6540 7111 6568
rect 7111 6540 7145 6568
rect 7145 6540 7157 6568
rect 7171 6568 7223 6592
rect 7171 6540 7183 6568
rect 7183 6540 7217 6568
rect 7217 6540 7223 6568
rect 7105 6495 7157 6526
rect 7105 6474 7111 6495
rect 7111 6474 7145 6495
rect 7145 6474 7157 6495
rect 7171 6495 7223 6526
rect 7171 6474 7183 6495
rect 7183 6474 7217 6495
rect 7217 6474 7223 6495
rect 7105 6422 7157 6460
rect 7171 6422 7223 6460
rect 7105 6408 7111 6422
rect 7111 6408 7157 6422
rect 7171 6408 7217 6422
rect 7217 6408 7223 6422
rect 7105 6342 7111 6394
rect 7111 6342 7157 6394
rect 7171 6342 7217 6394
rect 7217 6342 7223 6394
rect 7105 6275 7111 6327
rect 7111 6275 7157 6327
rect 7171 6275 7217 6327
rect 7217 6275 7223 6327
rect 7105 6208 7111 6260
rect 7111 6208 7157 6260
rect 7171 6208 7217 6260
rect 7217 6208 7223 6260
rect 7382 13877 7434 13892
rect 7382 13843 7388 13877
rect 7388 13843 7422 13877
rect 7422 13843 7434 13877
rect 7382 13840 7434 13843
rect 7448 13877 7500 13892
rect 7448 13843 7460 13877
rect 7460 13843 7494 13877
rect 7494 13843 7500 13877
rect 7448 13840 7500 13843
rect 7382 13799 7434 13826
rect 7382 13774 7388 13799
rect 7388 13774 7422 13799
rect 7422 13774 7434 13799
rect 7448 13799 7500 13826
rect 7448 13774 7460 13799
rect 7460 13774 7494 13799
rect 7494 13774 7500 13799
rect 7382 13722 7434 13760
rect 7382 13708 7388 13722
rect 7388 13708 7422 13722
rect 7422 13708 7434 13722
rect 7448 13722 7500 13760
rect 7448 13708 7460 13722
rect 7460 13708 7494 13722
rect 7494 13708 7500 13722
rect 7382 13688 7388 13694
rect 7388 13688 7422 13694
rect 7422 13688 7434 13694
rect 7382 13645 7434 13688
rect 7382 13642 7388 13645
rect 7388 13642 7422 13645
rect 7422 13642 7434 13645
rect 7448 13688 7460 13694
rect 7460 13688 7494 13694
rect 7494 13688 7500 13694
rect 7448 13645 7500 13688
rect 7448 13642 7460 13645
rect 7460 13642 7494 13645
rect 7494 13642 7500 13645
rect 7382 13611 7388 13628
rect 7388 13611 7422 13628
rect 7422 13611 7434 13628
rect 7382 13576 7434 13611
rect 7448 13611 7460 13628
rect 7460 13611 7494 13628
rect 7494 13611 7500 13628
rect 7448 13576 7500 13611
rect 7382 13534 7388 13562
rect 7388 13534 7422 13562
rect 7422 13534 7434 13562
rect 7382 13510 7434 13534
rect 7448 13534 7460 13562
rect 7460 13534 7494 13562
rect 7494 13534 7500 13562
rect 7448 13510 7500 13534
rect 7382 13491 7434 13495
rect 7382 13457 7388 13491
rect 7388 13457 7422 13491
rect 7422 13457 7434 13491
rect 7382 13443 7434 13457
rect 7448 13491 7500 13495
rect 7448 13457 7460 13491
rect 7460 13457 7494 13491
rect 7494 13457 7500 13491
rect 7448 13443 7500 13457
rect 7382 13414 7434 13428
rect 7382 13380 7388 13414
rect 7388 13380 7422 13414
rect 7422 13380 7434 13414
rect 7382 13376 7434 13380
rect 7448 13414 7500 13428
rect 7448 13380 7460 13414
rect 7460 13380 7494 13414
rect 7494 13380 7500 13414
rect 7448 13376 7500 13380
rect 7382 11840 7388 11892
rect 7388 11840 7434 11892
rect 7448 11840 7494 11892
rect 7494 11840 7500 11892
rect 7382 11774 7388 11826
rect 7388 11774 7434 11826
rect 7448 11774 7494 11826
rect 7494 11774 7500 11826
rect 7382 11708 7388 11760
rect 7388 11708 7434 11760
rect 7448 11708 7494 11760
rect 7494 11708 7500 11760
rect 7382 11642 7388 11694
rect 7388 11642 7434 11694
rect 7448 11642 7494 11694
rect 7494 11642 7500 11694
rect 7382 11576 7388 11628
rect 7388 11576 7434 11628
rect 7448 11576 7494 11628
rect 7494 11576 7500 11628
rect 7382 11510 7388 11562
rect 7388 11510 7434 11562
rect 7448 11510 7494 11562
rect 7494 11510 7500 11562
rect 7382 11443 7388 11495
rect 7388 11443 7434 11495
rect 7448 11443 7494 11495
rect 7494 11443 7500 11495
rect 7382 11380 7388 11428
rect 7388 11380 7434 11428
rect 7448 11380 7494 11428
rect 7494 11380 7500 11428
rect 7382 11376 7434 11380
rect 7448 11376 7500 11380
rect 7382 9844 7388 9896
rect 7388 9844 7434 9896
rect 7448 9844 7494 9896
rect 7494 9844 7500 9896
rect 7382 9778 7388 9830
rect 7388 9778 7434 9830
rect 7448 9778 7494 9830
rect 7494 9778 7500 9830
rect 7382 9712 7388 9764
rect 7388 9712 7434 9764
rect 7448 9712 7494 9764
rect 7494 9712 7500 9764
rect 7382 9646 7388 9698
rect 7388 9646 7434 9698
rect 7448 9646 7494 9698
rect 7494 9646 7500 9698
rect 7382 9580 7388 9632
rect 7388 9580 7434 9632
rect 7448 9580 7494 9632
rect 7494 9580 7500 9632
rect 7382 9514 7388 9566
rect 7388 9514 7434 9566
rect 7448 9514 7494 9566
rect 7494 9514 7500 9566
rect 7382 9447 7388 9499
rect 7388 9447 7434 9499
rect 7448 9447 7494 9499
rect 7494 9447 7500 9499
rect 7382 9380 7388 9432
rect 7388 9380 7434 9432
rect 7448 9380 7494 9432
rect 7494 9380 7500 9432
rect 7382 7840 7388 7892
rect 7388 7840 7434 7892
rect 7448 7840 7494 7892
rect 7494 7840 7500 7892
rect 7382 7774 7388 7826
rect 7388 7774 7434 7826
rect 7448 7774 7494 7826
rect 7494 7774 7500 7826
rect 7382 7708 7388 7760
rect 7388 7708 7434 7760
rect 7448 7708 7494 7760
rect 7494 7708 7500 7760
rect 7382 7642 7388 7694
rect 7388 7642 7434 7694
rect 7448 7642 7494 7694
rect 7494 7642 7500 7694
rect 7382 7576 7388 7628
rect 7388 7576 7434 7628
rect 7448 7576 7494 7628
rect 7494 7576 7500 7628
rect 7382 7510 7388 7562
rect 7388 7510 7434 7562
rect 7448 7510 7494 7562
rect 7494 7510 7500 7562
rect 7382 7443 7388 7495
rect 7388 7443 7434 7495
rect 7448 7443 7494 7495
rect 7494 7443 7500 7495
rect 7382 7380 7388 7428
rect 7388 7380 7434 7428
rect 7448 7380 7494 7428
rect 7494 7380 7500 7428
rect 7382 7376 7434 7380
rect 7448 7376 7500 7380
rect 7382 5844 7388 5896
rect 7388 5844 7434 5896
rect 7448 5844 7494 5896
rect 7494 5844 7500 5896
rect 7382 5778 7388 5830
rect 7388 5778 7434 5830
rect 7448 5778 7494 5830
rect 7494 5778 7500 5830
rect 7382 5712 7388 5764
rect 7388 5712 7434 5764
rect 7448 5712 7494 5764
rect 7494 5712 7500 5764
rect 7382 5646 7388 5698
rect 7388 5646 7434 5698
rect 7448 5646 7494 5698
rect 7494 5646 7500 5698
rect 7382 5580 7388 5632
rect 7388 5580 7434 5632
rect 7448 5580 7494 5632
rect 7494 5580 7500 5632
rect 7382 5514 7388 5566
rect 7388 5514 7434 5566
rect 7448 5514 7494 5566
rect 7494 5514 7500 5566
rect 7382 5447 7388 5499
rect 7388 5447 7434 5499
rect 7448 5447 7494 5499
rect 7494 5447 7500 5499
rect 7382 5380 7388 5432
rect 7388 5380 7434 5432
rect 7448 5380 7494 5432
rect 7494 5380 7500 5432
rect 7659 14345 7711 14390
rect 7659 14338 7665 14345
rect 7665 14338 7699 14345
rect 7699 14338 7711 14345
rect 7725 14345 7777 14390
rect 8213 14668 8265 14720
rect 8279 14668 8331 14720
rect 8213 14602 8265 14654
rect 8279 14602 8331 14654
rect 8213 14536 8265 14588
rect 8279 14536 8331 14588
rect 8213 14470 8265 14522
rect 8279 14470 8331 14522
rect 8213 14404 8265 14456
rect 8279 14404 8331 14456
rect 7725 14338 7737 14345
rect 7737 14338 7771 14345
rect 7771 14338 7777 14345
rect 7659 14311 7665 14323
rect 7665 14311 7699 14323
rect 7699 14311 7711 14323
rect 7659 14271 7711 14311
rect 7725 14311 7737 14323
rect 7737 14311 7771 14323
rect 7771 14311 7777 14323
rect 7725 14271 7777 14311
rect 7659 14233 7665 14256
rect 7665 14233 7699 14256
rect 7699 14233 7711 14256
rect 7659 14204 7711 14233
rect 7725 14233 7737 14256
rect 7737 14233 7771 14256
rect 7771 14233 7777 14256
rect 7725 14204 7777 14233
rect 7659 12714 7711 12720
rect 7659 12680 7665 12714
rect 7665 12680 7699 12714
rect 7699 12680 7711 12714
rect 7659 12668 7711 12680
rect 7725 12714 7777 12720
rect 7725 12680 7737 12714
rect 7737 12680 7771 12714
rect 7771 12680 7777 12714
rect 7725 12668 7777 12680
rect 7659 12641 7711 12654
rect 7659 12607 7665 12641
rect 7665 12607 7699 12641
rect 7699 12607 7711 12641
rect 7659 12602 7711 12607
rect 7725 12641 7777 12654
rect 7725 12607 7737 12641
rect 7737 12607 7771 12641
rect 7771 12607 7777 12641
rect 7725 12602 7777 12607
rect 7659 12568 7711 12588
rect 7659 12536 7665 12568
rect 7665 12536 7699 12568
rect 7699 12536 7711 12568
rect 7725 12568 7777 12588
rect 7725 12536 7737 12568
rect 7737 12536 7771 12568
rect 7771 12536 7777 12568
rect 7659 12495 7711 12522
rect 7659 12470 7665 12495
rect 7665 12470 7699 12495
rect 7699 12470 7711 12495
rect 7725 12495 7777 12522
rect 7725 12470 7737 12495
rect 7737 12470 7771 12495
rect 7771 12470 7777 12495
rect 7659 12422 7711 12456
rect 7725 12422 7777 12456
rect 7659 12404 7665 12422
rect 7665 12404 7711 12422
rect 7725 12404 7771 12422
rect 7771 12404 7777 12422
rect 7659 12338 7665 12390
rect 7665 12338 7711 12390
rect 7725 12338 7771 12390
rect 7771 12338 7777 12390
rect 7659 12271 7665 12323
rect 7665 12271 7711 12323
rect 7725 12271 7771 12323
rect 7771 12271 7777 12323
rect 7659 12204 7665 12256
rect 7665 12204 7711 12256
rect 7725 12204 7771 12256
rect 7771 12204 7777 12256
rect 7659 10714 7711 10724
rect 7659 10680 7665 10714
rect 7665 10680 7699 10714
rect 7699 10680 7711 10714
rect 7659 10672 7711 10680
rect 7725 10714 7777 10724
rect 7725 10680 7737 10714
rect 7737 10680 7771 10714
rect 7771 10680 7777 10714
rect 7725 10672 7777 10680
rect 7659 10641 7711 10658
rect 7659 10607 7665 10641
rect 7665 10607 7699 10641
rect 7699 10607 7711 10641
rect 7659 10606 7711 10607
rect 7725 10641 7777 10658
rect 7725 10607 7737 10641
rect 7737 10607 7771 10641
rect 7771 10607 7777 10641
rect 7725 10606 7777 10607
rect 7659 10568 7711 10592
rect 7659 10540 7665 10568
rect 7665 10540 7699 10568
rect 7699 10540 7711 10568
rect 7725 10568 7777 10592
rect 7725 10540 7737 10568
rect 7737 10540 7771 10568
rect 7771 10540 7777 10568
rect 7659 10495 7711 10526
rect 7659 10474 7665 10495
rect 7665 10474 7699 10495
rect 7699 10474 7711 10495
rect 7725 10495 7777 10526
rect 7725 10474 7737 10495
rect 7737 10474 7771 10495
rect 7771 10474 7777 10495
rect 7659 10422 7711 10460
rect 7725 10422 7777 10460
rect 7659 10408 7665 10422
rect 7665 10408 7711 10422
rect 7725 10408 7771 10422
rect 7771 10408 7777 10422
rect 7659 10342 7665 10394
rect 7665 10342 7711 10394
rect 7725 10342 7771 10394
rect 7771 10342 7777 10394
rect 7659 10275 7665 10327
rect 7665 10275 7711 10327
rect 7725 10275 7771 10327
rect 7771 10275 7777 10327
rect 7659 10208 7665 10260
rect 7665 10208 7711 10260
rect 7725 10208 7771 10260
rect 7771 10208 7777 10260
rect 7659 8714 7711 8720
rect 7659 8680 7665 8714
rect 7665 8680 7699 8714
rect 7699 8680 7711 8714
rect 7659 8668 7711 8680
rect 7725 8714 7777 8720
rect 7725 8680 7737 8714
rect 7737 8680 7771 8714
rect 7771 8680 7777 8714
rect 7725 8668 7777 8680
rect 7659 8641 7711 8654
rect 7659 8607 7665 8641
rect 7665 8607 7699 8641
rect 7699 8607 7711 8641
rect 7659 8602 7711 8607
rect 7725 8641 7777 8654
rect 7725 8607 7737 8641
rect 7737 8607 7771 8641
rect 7771 8607 7777 8641
rect 7725 8602 7777 8607
rect 7659 8568 7711 8588
rect 7659 8536 7665 8568
rect 7665 8536 7699 8568
rect 7699 8536 7711 8568
rect 7725 8568 7777 8588
rect 7725 8536 7737 8568
rect 7737 8536 7771 8568
rect 7771 8536 7777 8568
rect 7659 8495 7711 8522
rect 7659 8470 7665 8495
rect 7665 8470 7699 8495
rect 7699 8470 7711 8495
rect 7725 8495 7777 8522
rect 7725 8470 7737 8495
rect 7737 8470 7771 8495
rect 7771 8470 7777 8495
rect 7659 8422 7711 8456
rect 7725 8422 7777 8456
rect 7659 8404 7665 8422
rect 7665 8404 7711 8422
rect 7725 8404 7771 8422
rect 7771 8404 7777 8422
rect 7659 8338 7665 8390
rect 7665 8338 7711 8390
rect 7725 8338 7771 8390
rect 7771 8338 7777 8390
rect 7659 8271 7665 8323
rect 7665 8271 7711 8323
rect 7725 8271 7771 8323
rect 7771 8271 7777 8323
rect 7659 8204 7665 8256
rect 7665 8204 7711 8256
rect 7725 8204 7771 8256
rect 7771 8204 7777 8256
rect 7659 6714 7711 6724
rect 7659 6680 7665 6714
rect 7665 6680 7699 6714
rect 7699 6680 7711 6714
rect 7659 6672 7711 6680
rect 7725 6714 7777 6724
rect 7725 6680 7737 6714
rect 7737 6680 7771 6714
rect 7771 6680 7777 6714
rect 7725 6672 7777 6680
rect 7659 6641 7711 6658
rect 7659 6607 7665 6641
rect 7665 6607 7699 6641
rect 7699 6607 7711 6641
rect 7659 6606 7711 6607
rect 7725 6641 7777 6658
rect 7725 6607 7737 6641
rect 7737 6607 7771 6641
rect 7771 6607 7777 6641
rect 7725 6606 7777 6607
rect 7659 6568 7711 6592
rect 7659 6540 7665 6568
rect 7665 6540 7699 6568
rect 7699 6540 7711 6568
rect 7725 6568 7777 6592
rect 7725 6540 7737 6568
rect 7737 6540 7771 6568
rect 7771 6540 7777 6568
rect 7659 6495 7711 6526
rect 7659 6474 7665 6495
rect 7665 6474 7699 6495
rect 7699 6474 7711 6495
rect 7725 6495 7777 6526
rect 7725 6474 7737 6495
rect 7737 6474 7771 6495
rect 7771 6474 7777 6495
rect 7659 6422 7711 6460
rect 7725 6422 7777 6460
rect 7659 6408 7665 6422
rect 7665 6408 7711 6422
rect 7725 6408 7771 6422
rect 7771 6408 7777 6422
rect 7659 6342 7665 6394
rect 7665 6342 7711 6394
rect 7725 6342 7771 6394
rect 7771 6342 7777 6394
rect 7659 6275 7665 6327
rect 7665 6275 7711 6327
rect 7725 6275 7771 6327
rect 7771 6275 7777 6327
rect 7659 6208 7665 6260
rect 7665 6208 7711 6260
rect 7725 6208 7771 6260
rect 7771 6208 7777 6260
rect 7936 13877 7988 13892
rect 7936 13843 7942 13877
rect 7942 13843 7976 13877
rect 7976 13843 7988 13877
rect 7936 13840 7988 13843
rect 8002 13877 8054 13892
rect 8002 13843 8014 13877
rect 8014 13843 8048 13877
rect 8048 13843 8054 13877
rect 8002 13840 8054 13843
rect 7936 13799 7988 13826
rect 7936 13774 7942 13799
rect 7942 13774 7976 13799
rect 7976 13774 7988 13799
rect 8002 13799 8054 13826
rect 8002 13774 8014 13799
rect 8014 13774 8048 13799
rect 8048 13774 8054 13799
rect 7936 13722 7988 13760
rect 7936 13708 7942 13722
rect 7942 13708 7976 13722
rect 7976 13708 7988 13722
rect 8002 13722 8054 13760
rect 8002 13708 8014 13722
rect 8014 13708 8048 13722
rect 8048 13708 8054 13722
rect 7936 13688 7942 13694
rect 7942 13688 7976 13694
rect 7976 13688 7988 13694
rect 7936 13645 7988 13688
rect 7936 13642 7942 13645
rect 7942 13642 7976 13645
rect 7976 13642 7988 13645
rect 8002 13688 8014 13694
rect 8014 13688 8048 13694
rect 8048 13688 8054 13694
rect 8002 13645 8054 13688
rect 8002 13642 8014 13645
rect 8014 13642 8048 13645
rect 8048 13642 8054 13645
rect 7936 13611 7942 13628
rect 7942 13611 7976 13628
rect 7976 13611 7988 13628
rect 7936 13576 7988 13611
rect 8002 13611 8014 13628
rect 8014 13611 8048 13628
rect 8048 13611 8054 13628
rect 8002 13576 8054 13611
rect 7936 13534 7942 13562
rect 7942 13534 7976 13562
rect 7976 13534 7988 13562
rect 7936 13510 7988 13534
rect 8002 13534 8014 13562
rect 8014 13534 8048 13562
rect 8048 13534 8054 13562
rect 8002 13510 8054 13534
rect 7936 13491 7988 13495
rect 7936 13457 7942 13491
rect 7942 13457 7976 13491
rect 7976 13457 7988 13491
rect 7936 13443 7988 13457
rect 8002 13491 8054 13495
rect 8002 13457 8014 13491
rect 8014 13457 8048 13491
rect 8048 13457 8054 13491
rect 8002 13443 8054 13457
rect 7936 13414 7988 13428
rect 7936 13380 7942 13414
rect 7942 13380 7976 13414
rect 7976 13380 7988 13414
rect 7936 13376 7988 13380
rect 8002 13414 8054 13428
rect 8002 13380 8014 13414
rect 8014 13380 8048 13414
rect 8048 13380 8054 13414
rect 8002 13376 8054 13380
rect 7936 11840 7942 11892
rect 7942 11840 7988 11892
rect 8002 11840 8048 11892
rect 8048 11840 8054 11892
rect 7936 11774 7942 11826
rect 7942 11774 7988 11826
rect 8002 11774 8048 11826
rect 8048 11774 8054 11826
rect 7936 11708 7942 11760
rect 7942 11708 7988 11760
rect 8002 11708 8048 11760
rect 8048 11708 8054 11760
rect 7936 11642 7942 11694
rect 7942 11642 7988 11694
rect 8002 11642 8048 11694
rect 8048 11642 8054 11694
rect 7936 11576 7942 11628
rect 7942 11576 7988 11628
rect 8002 11576 8048 11628
rect 8048 11576 8054 11628
rect 7936 11510 7942 11562
rect 7942 11510 7988 11562
rect 8002 11510 8048 11562
rect 8048 11510 8054 11562
rect 7936 11443 7942 11495
rect 7942 11443 7988 11495
rect 8002 11443 8048 11495
rect 8048 11443 8054 11495
rect 7936 11380 7942 11428
rect 7942 11380 7988 11428
rect 8002 11380 8048 11428
rect 8048 11380 8054 11428
rect 7936 11376 7988 11380
rect 8002 11376 8054 11380
rect 7936 9844 7942 9896
rect 7942 9844 7988 9896
rect 8002 9844 8048 9896
rect 8048 9844 8054 9896
rect 7936 9778 7942 9830
rect 7942 9778 7988 9830
rect 8002 9778 8048 9830
rect 8048 9778 8054 9830
rect 7936 9712 7942 9764
rect 7942 9712 7988 9764
rect 8002 9712 8048 9764
rect 8048 9712 8054 9764
rect 7936 9646 7942 9698
rect 7942 9646 7988 9698
rect 8002 9646 8048 9698
rect 8048 9646 8054 9698
rect 7936 9580 7942 9632
rect 7942 9580 7988 9632
rect 8002 9580 8048 9632
rect 8048 9580 8054 9632
rect 7936 9514 7942 9566
rect 7942 9514 7988 9566
rect 8002 9514 8048 9566
rect 8048 9514 8054 9566
rect 7936 9447 7942 9499
rect 7942 9447 7988 9499
rect 8002 9447 8048 9499
rect 8048 9447 8054 9499
rect 7936 9380 7942 9432
rect 7942 9380 7988 9432
rect 8002 9380 8048 9432
rect 8048 9380 8054 9432
rect 7936 7840 7942 7892
rect 7942 7840 7988 7892
rect 8002 7840 8048 7892
rect 8048 7840 8054 7892
rect 7936 7774 7942 7826
rect 7942 7774 7988 7826
rect 8002 7774 8048 7826
rect 8048 7774 8054 7826
rect 7936 7708 7942 7760
rect 7942 7708 7988 7760
rect 8002 7708 8048 7760
rect 8048 7708 8054 7760
rect 7936 7642 7942 7694
rect 7942 7642 7988 7694
rect 8002 7642 8048 7694
rect 8048 7642 8054 7694
rect 7936 7576 7942 7628
rect 7942 7576 7988 7628
rect 8002 7576 8048 7628
rect 8048 7576 8054 7628
rect 7936 7510 7942 7562
rect 7942 7510 7988 7562
rect 8002 7510 8048 7562
rect 8048 7510 8054 7562
rect 7936 7443 7942 7495
rect 7942 7443 7988 7495
rect 8002 7443 8048 7495
rect 8048 7443 8054 7495
rect 7936 7380 7942 7428
rect 7942 7380 7988 7428
rect 8002 7380 8048 7428
rect 8048 7380 8054 7428
rect 7936 7376 7988 7380
rect 8002 7376 8054 7380
rect 7936 5844 7942 5896
rect 7942 5844 7988 5896
rect 8002 5844 8048 5896
rect 8048 5844 8054 5896
rect 7936 5778 7942 5830
rect 7942 5778 7988 5830
rect 8002 5778 8048 5830
rect 8048 5778 8054 5830
rect 7936 5712 7942 5764
rect 7942 5712 7988 5764
rect 8002 5712 8048 5764
rect 8048 5712 8054 5764
rect 7936 5646 7942 5698
rect 7942 5646 7988 5698
rect 8002 5646 8048 5698
rect 8048 5646 8054 5698
rect 7936 5580 7942 5632
rect 7942 5580 7988 5632
rect 8002 5580 8048 5632
rect 8048 5580 8054 5632
rect 7936 5514 7942 5566
rect 7942 5514 7988 5566
rect 8002 5514 8048 5566
rect 8048 5514 8054 5566
rect 7936 5447 7942 5499
rect 7942 5447 7988 5499
rect 8002 5447 8048 5499
rect 8048 5447 8054 5499
rect 7936 5380 7942 5432
rect 7942 5380 7988 5432
rect 8002 5380 8048 5432
rect 8048 5380 8054 5432
rect 8213 14345 8265 14390
rect 8213 14338 8219 14345
rect 8219 14338 8253 14345
rect 8253 14338 8265 14345
rect 8279 14345 8331 14390
rect 8767 14668 8819 14720
rect 8833 14668 8885 14720
rect 8767 14602 8819 14654
rect 8833 14602 8885 14654
rect 8767 14536 8819 14588
rect 8833 14536 8885 14588
rect 8767 14470 8819 14522
rect 8833 14470 8885 14522
rect 8767 14404 8819 14456
rect 8833 14404 8885 14456
rect 8279 14338 8291 14345
rect 8291 14338 8325 14345
rect 8325 14338 8331 14345
rect 8213 14311 8219 14323
rect 8219 14311 8253 14323
rect 8253 14311 8265 14323
rect 8213 14271 8265 14311
rect 8279 14311 8291 14323
rect 8291 14311 8325 14323
rect 8325 14311 8331 14323
rect 8279 14271 8331 14311
rect 8213 14233 8219 14256
rect 8219 14233 8253 14256
rect 8253 14233 8265 14256
rect 8213 14204 8265 14233
rect 8279 14233 8291 14256
rect 8291 14233 8325 14256
rect 8325 14233 8331 14256
rect 8279 14204 8331 14233
rect 8213 12714 8265 12720
rect 8213 12680 8219 12714
rect 8219 12680 8253 12714
rect 8253 12680 8265 12714
rect 8213 12668 8265 12680
rect 8279 12714 8331 12720
rect 8279 12680 8291 12714
rect 8291 12680 8325 12714
rect 8325 12680 8331 12714
rect 8279 12668 8331 12680
rect 8213 12641 8265 12654
rect 8213 12607 8219 12641
rect 8219 12607 8253 12641
rect 8253 12607 8265 12641
rect 8213 12602 8265 12607
rect 8279 12641 8331 12654
rect 8279 12607 8291 12641
rect 8291 12607 8325 12641
rect 8325 12607 8331 12641
rect 8279 12602 8331 12607
rect 8213 12568 8265 12588
rect 8213 12536 8219 12568
rect 8219 12536 8253 12568
rect 8253 12536 8265 12568
rect 8279 12568 8331 12588
rect 8279 12536 8291 12568
rect 8291 12536 8325 12568
rect 8325 12536 8331 12568
rect 8213 12495 8265 12522
rect 8213 12470 8219 12495
rect 8219 12470 8253 12495
rect 8253 12470 8265 12495
rect 8279 12495 8331 12522
rect 8279 12470 8291 12495
rect 8291 12470 8325 12495
rect 8325 12470 8331 12495
rect 8213 12422 8265 12456
rect 8279 12422 8331 12456
rect 8213 12404 8219 12422
rect 8219 12404 8265 12422
rect 8279 12404 8325 12422
rect 8325 12404 8331 12422
rect 8213 12338 8219 12390
rect 8219 12338 8265 12390
rect 8279 12338 8325 12390
rect 8325 12338 8331 12390
rect 8213 12271 8219 12323
rect 8219 12271 8265 12323
rect 8279 12271 8325 12323
rect 8325 12271 8331 12323
rect 8213 12204 8219 12256
rect 8219 12204 8265 12256
rect 8279 12204 8325 12256
rect 8325 12204 8331 12256
rect 8213 10714 8265 10724
rect 8213 10680 8219 10714
rect 8219 10680 8253 10714
rect 8253 10680 8265 10714
rect 8213 10672 8265 10680
rect 8279 10714 8331 10724
rect 8279 10680 8291 10714
rect 8291 10680 8325 10714
rect 8325 10680 8331 10714
rect 8279 10672 8331 10680
rect 8213 10641 8265 10658
rect 8213 10607 8219 10641
rect 8219 10607 8253 10641
rect 8253 10607 8265 10641
rect 8213 10606 8265 10607
rect 8279 10641 8331 10658
rect 8279 10607 8291 10641
rect 8291 10607 8325 10641
rect 8325 10607 8331 10641
rect 8279 10606 8331 10607
rect 8213 10568 8265 10592
rect 8213 10540 8219 10568
rect 8219 10540 8253 10568
rect 8253 10540 8265 10568
rect 8279 10568 8331 10592
rect 8279 10540 8291 10568
rect 8291 10540 8325 10568
rect 8325 10540 8331 10568
rect 8213 10495 8265 10526
rect 8213 10474 8219 10495
rect 8219 10474 8253 10495
rect 8253 10474 8265 10495
rect 8279 10495 8331 10526
rect 8279 10474 8291 10495
rect 8291 10474 8325 10495
rect 8325 10474 8331 10495
rect 8213 10422 8265 10460
rect 8279 10422 8331 10460
rect 8213 10408 8219 10422
rect 8219 10408 8265 10422
rect 8279 10408 8325 10422
rect 8325 10408 8331 10422
rect 8213 10342 8219 10394
rect 8219 10342 8265 10394
rect 8279 10342 8325 10394
rect 8325 10342 8331 10394
rect 8213 10275 8219 10327
rect 8219 10275 8265 10327
rect 8279 10275 8325 10327
rect 8325 10275 8331 10327
rect 8213 10208 8219 10260
rect 8219 10208 8265 10260
rect 8279 10208 8325 10260
rect 8325 10208 8331 10260
rect 8213 8714 8265 8720
rect 8213 8680 8219 8714
rect 8219 8680 8253 8714
rect 8253 8680 8265 8714
rect 8213 8668 8265 8680
rect 8279 8714 8331 8720
rect 8279 8680 8291 8714
rect 8291 8680 8325 8714
rect 8325 8680 8331 8714
rect 8279 8668 8331 8680
rect 8213 8641 8265 8654
rect 8213 8607 8219 8641
rect 8219 8607 8253 8641
rect 8253 8607 8265 8641
rect 8213 8602 8265 8607
rect 8279 8641 8331 8654
rect 8279 8607 8291 8641
rect 8291 8607 8325 8641
rect 8325 8607 8331 8641
rect 8279 8602 8331 8607
rect 8213 8568 8265 8588
rect 8213 8536 8219 8568
rect 8219 8536 8253 8568
rect 8253 8536 8265 8568
rect 8279 8568 8331 8588
rect 8279 8536 8291 8568
rect 8291 8536 8325 8568
rect 8325 8536 8331 8568
rect 8213 8495 8265 8522
rect 8213 8470 8219 8495
rect 8219 8470 8253 8495
rect 8253 8470 8265 8495
rect 8279 8495 8331 8522
rect 8279 8470 8291 8495
rect 8291 8470 8325 8495
rect 8325 8470 8331 8495
rect 8213 8422 8265 8456
rect 8279 8422 8331 8456
rect 8213 8404 8219 8422
rect 8219 8404 8265 8422
rect 8279 8404 8325 8422
rect 8325 8404 8331 8422
rect 8213 8338 8219 8390
rect 8219 8338 8265 8390
rect 8279 8338 8325 8390
rect 8325 8338 8331 8390
rect 8213 8271 8219 8323
rect 8219 8271 8265 8323
rect 8279 8271 8325 8323
rect 8325 8271 8331 8323
rect 8213 8204 8219 8256
rect 8219 8204 8265 8256
rect 8279 8204 8325 8256
rect 8325 8204 8331 8256
rect 8213 6714 8265 6724
rect 8213 6680 8219 6714
rect 8219 6680 8253 6714
rect 8253 6680 8265 6714
rect 8213 6672 8265 6680
rect 8279 6714 8331 6724
rect 8279 6680 8291 6714
rect 8291 6680 8325 6714
rect 8325 6680 8331 6714
rect 8279 6672 8331 6680
rect 8213 6641 8265 6658
rect 8213 6607 8219 6641
rect 8219 6607 8253 6641
rect 8253 6607 8265 6641
rect 8213 6606 8265 6607
rect 8279 6641 8331 6658
rect 8279 6607 8291 6641
rect 8291 6607 8325 6641
rect 8325 6607 8331 6641
rect 8279 6606 8331 6607
rect 8213 6568 8265 6592
rect 8213 6540 8219 6568
rect 8219 6540 8253 6568
rect 8253 6540 8265 6568
rect 8279 6568 8331 6592
rect 8279 6540 8291 6568
rect 8291 6540 8325 6568
rect 8325 6540 8331 6568
rect 8213 6495 8265 6526
rect 8213 6474 8219 6495
rect 8219 6474 8253 6495
rect 8253 6474 8265 6495
rect 8279 6495 8331 6526
rect 8279 6474 8291 6495
rect 8291 6474 8325 6495
rect 8325 6474 8331 6495
rect 8213 6422 8265 6460
rect 8279 6422 8331 6460
rect 8213 6408 8219 6422
rect 8219 6408 8265 6422
rect 8279 6408 8325 6422
rect 8325 6408 8331 6422
rect 8213 6342 8219 6394
rect 8219 6342 8265 6394
rect 8279 6342 8325 6394
rect 8325 6342 8331 6394
rect 8213 6275 8219 6327
rect 8219 6275 8265 6327
rect 8279 6275 8325 6327
rect 8325 6275 8331 6327
rect 8213 6208 8219 6260
rect 8219 6208 8265 6260
rect 8279 6208 8325 6260
rect 8325 6208 8331 6260
rect 8490 13877 8542 13892
rect 8490 13843 8496 13877
rect 8496 13843 8530 13877
rect 8530 13843 8542 13877
rect 8490 13840 8542 13843
rect 8556 13877 8608 13892
rect 8556 13843 8568 13877
rect 8568 13843 8602 13877
rect 8602 13843 8608 13877
rect 8556 13840 8608 13843
rect 8490 13799 8542 13826
rect 8490 13774 8496 13799
rect 8496 13774 8530 13799
rect 8530 13774 8542 13799
rect 8556 13799 8608 13826
rect 8556 13774 8568 13799
rect 8568 13774 8602 13799
rect 8602 13774 8608 13799
rect 8490 13722 8542 13760
rect 8490 13708 8496 13722
rect 8496 13708 8530 13722
rect 8530 13708 8542 13722
rect 8556 13722 8608 13760
rect 8556 13708 8568 13722
rect 8568 13708 8602 13722
rect 8602 13708 8608 13722
rect 8490 13688 8496 13694
rect 8496 13688 8530 13694
rect 8530 13688 8542 13694
rect 8490 13645 8542 13688
rect 8490 13642 8496 13645
rect 8496 13642 8530 13645
rect 8530 13642 8542 13645
rect 8556 13688 8568 13694
rect 8568 13688 8602 13694
rect 8602 13688 8608 13694
rect 8556 13645 8608 13688
rect 8556 13642 8568 13645
rect 8568 13642 8602 13645
rect 8602 13642 8608 13645
rect 8490 13611 8496 13628
rect 8496 13611 8530 13628
rect 8530 13611 8542 13628
rect 8490 13576 8542 13611
rect 8556 13611 8568 13628
rect 8568 13611 8602 13628
rect 8602 13611 8608 13628
rect 8556 13576 8608 13611
rect 8490 13534 8496 13562
rect 8496 13534 8530 13562
rect 8530 13534 8542 13562
rect 8490 13510 8542 13534
rect 8556 13534 8568 13562
rect 8568 13534 8602 13562
rect 8602 13534 8608 13562
rect 8556 13510 8608 13534
rect 8490 13491 8542 13495
rect 8490 13457 8496 13491
rect 8496 13457 8530 13491
rect 8530 13457 8542 13491
rect 8490 13443 8542 13457
rect 8556 13491 8608 13495
rect 8556 13457 8568 13491
rect 8568 13457 8602 13491
rect 8602 13457 8608 13491
rect 8556 13443 8608 13457
rect 8490 13414 8542 13428
rect 8490 13380 8496 13414
rect 8496 13380 8530 13414
rect 8530 13380 8542 13414
rect 8490 13376 8542 13380
rect 8556 13414 8608 13428
rect 8556 13380 8568 13414
rect 8568 13380 8602 13414
rect 8602 13380 8608 13414
rect 8556 13376 8608 13380
rect 8490 11840 8496 11892
rect 8496 11840 8542 11892
rect 8556 11840 8602 11892
rect 8602 11840 8608 11892
rect 8490 11774 8496 11826
rect 8496 11774 8542 11826
rect 8556 11774 8602 11826
rect 8602 11774 8608 11826
rect 8490 11708 8496 11760
rect 8496 11708 8542 11760
rect 8556 11708 8602 11760
rect 8602 11708 8608 11760
rect 8490 11642 8496 11694
rect 8496 11642 8542 11694
rect 8556 11642 8602 11694
rect 8602 11642 8608 11694
rect 8490 11576 8496 11628
rect 8496 11576 8542 11628
rect 8556 11576 8602 11628
rect 8602 11576 8608 11628
rect 8490 11510 8496 11562
rect 8496 11510 8542 11562
rect 8556 11510 8602 11562
rect 8602 11510 8608 11562
rect 8490 11443 8496 11495
rect 8496 11443 8542 11495
rect 8556 11443 8602 11495
rect 8602 11443 8608 11495
rect 8490 11380 8496 11428
rect 8496 11380 8542 11428
rect 8556 11380 8602 11428
rect 8602 11380 8608 11428
rect 8490 11376 8542 11380
rect 8556 11376 8608 11380
rect 8490 9844 8496 9896
rect 8496 9844 8542 9896
rect 8556 9844 8602 9896
rect 8602 9844 8608 9896
rect 8490 9778 8496 9830
rect 8496 9778 8542 9830
rect 8556 9778 8602 9830
rect 8602 9778 8608 9830
rect 8490 9712 8496 9764
rect 8496 9712 8542 9764
rect 8556 9712 8602 9764
rect 8602 9712 8608 9764
rect 8490 9646 8496 9698
rect 8496 9646 8542 9698
rect 8556 9646 8602 9698
rect 8602 9646 8608 9698
rect 8490 9580 8496 9632
rect 8496 9580 8542 9632
rect 8556 9580 8602 9632
rect 8602 9580 8608 9632
rect 8490 9514 8496 9566
rect 8496 9514 8542 9566
rect 8556 9514 8602 9566
rect 8602 9514 8608 9566
rect 8490 9447 8496 9499
rect 8496 9447 8542 9499
rect 8556 9447 8602 9499
rect 8602 9447 8608 9499
rect 8490 9380 8496 9432
rect 8496 9380 8542 9432
rect 8556 9380 8602 9432
rect 8602 9380 8608 9432
rect 8490 7840 8496 7892
rect 8496 7840 8542 7892
rect 8556 7840 8602 7892
rect 8602 7840 8608 7892
rect 8490 7774 8496 7826
rect 8496 7774 8542 7826
rect 8556 7774 8602 7826
rect 8602 7774 8608 7826
rect 8490 7708 8496 7760
rect 8496 7708 8542 7760
rect 8556 7708 8602 7760
rect 8602 7708 8608 7760
rect 8490 7642 8496 7694
rect 8496 7642 8542 7694
rect 8556 7642 8602 7694
rect 8602 7642 8608 7694
rect 8490 7576 8496 7628
rect 8496 7576 8542 7628
rect 8556 7576 8602 7628
rect 8602 7576 8608 7628
rect 8490 7510 8496 7562
rect 8496 7510 8542 7562
rect 8556 7510 8602 7562
rect 8602 7510 8608 7562
rect 8490 7443 8496 7495
rect 8496 7443 8542 7495
rect 8556 7443 8602 7495
rect 8602 7443 8608 7495
rect 8490 7380 8496 7428
rect 8496 7380 8542 7428
rect 8556 7380 8602 7428
rect 8602 7380 8608 7428
rect 8490 7376 8542 7380
rect 8556 7376 8608 7380
rect 8490 5844 8496 5896
rect 8496 5844 8542 5896
rect 8556 5844 8602 5896
rect 8602 5844 8608 5896
rect 8490 5778 8496 5830
rect 8496 5778 8542 5830
rect 8556 5778 8602 5830
rect 8602 5778 8608 5830
rect 8490 5712 8496 5764
rect 8496 5712 8542 5764
rect 8556 5712 8602 5764
rect 8602 5712 8608 5764
rect 8490 5646 8496 5698
rect 8496 5646 8542 5698
rect 8556 5646 8602 5698
rect 8602 5646 8608 5698
rect 8490 5580 8496 5632
rect 8496 5580 8542 5632
rect 8556 5580 8602 5632
rect 8602 5580 8608 5632
rect 8490 5514 8496 5566
rect 8496 5514 8542 5566
rect 8556 5514 8602 5566
rect 8602 5514 8608 5566
rect 8490 5447 8496 5499
rect 8496 5447 8542 5499
rect 8556 5447 8602 5499
rect 8602 5447 8608 5499
rect 8490 5380 8496 5432
rect 8496 5380 8542 5432
rect 8556 5380 8602 5432
rect 8602 5380 8608 5432
rect 8767 14345 8819 14390
rect 8767 14338 8773 14345
rect 8773 14338 8807 14345
rect 8807 14338 8819 14345
rect 8833 14345 8885 14390
rect 9321 14668 9373 14720
rect 9387 14668 9439 14720
rect 9321 14602 9373 14654
rect 9387 14602 9439 14654
rect 9321 14536 9373 14588
rect 9387 14536 9439 14588
rect 9321 14470 9373 14522
rect 9387 14470 9439 14522
rect 9321 14404 9373 14456
rect 9387 14404 9439 14456
rect 8833 14338 8845 14345
rect 8845 14338 8879 14345
rect 8879 14338 8885 14345
rect 8767 14311 8773 14323
rect 8773 14311 8807 14323
rect 8807 14311 8819 14323
rect 8767 14271 8819 14311
rect 8833 14311 8845 14323
rect 8845 14311 8879 14323
rect 8879 14311 8885 14323
rect 8833 14271 8885 14311
rect 8767 14233 8773 14256
rect 8773 14233 8807 14256
rect 8807 14233 8819 14256
rect 8767 14204 8819 14233
rect 8833 14233 8845 14256
rect 8845 14233 8879 14256
rect 8879 14233 8885 14256
rect 8833 14204 8885 14233
rect 8767 12714 8819 12720
rect 8767 12680 8773 12714
rect 8773 12680 8807 12714
rect 8807 12680 8819 12714
rect 8767 12668 8819 12680
rect 8833 12714 8885 12720
rect 8833 12680 8845 12714
rect 8845 12680 8879 12714
rect 8879 12680 8885 12714
rect 8833 12668 8885 12680
rect 8767 12641 8819 12654
rect 8767 12607 8773 12641
rect 8773 12607 8807 12641
rect 8807 12607 8819 12641
rect 8767 12602 8819 12607
rect 8833 12641 8885 12654
rect 8833 12607 8845 12641
rect 8845 12607 8879 12641
rect 8879 12607 8885 12641
rect 8833 12602 8885 12607
rect 8767 12568 8819 12588
rect 8767 12536 8773 12568
rect 8773 12536 8807 12568
rect 8807 12536 8819 12568
rect 8833 12568 8885 12588
rect 8833 12536 8845 12568
rect 8845 12536 8879 12568
rect 8879 12536 8885 12568
rect 8767 12495 8819 12522
rect 8767 12470 8773 12495
rect 8773 12470 8807 12495
rect 8807 12470 8819 12495
rect 8833 12495 8885 12522
rect 8833 12470 8845 12495
rect 8845 12470 8879 12495
rect 8879 12470 8885 12495
rect 8767 12422 8819 12456
rect 8833 12422 8885 12456
rect 8767 12404 8773 12422
rect 8773 12404 8819 12422
rect 8833 12404 8879 12422
rect 8879 12404 8885 12422
rect 8767 12338 8773 12390
rect 8773 12338 8819 12390
rect 8833 12338 8879 12390
rect 8879 12338 8885 12390
rect 8767 12271 8773 12323
rect 8773 12271 8819 12323
rect 8833 12271 8879 12323
rect 8879 12271 8885 12323
rect 8767 12204 8773 12256
rect 8773 12204 8819 12256
rect 8833 12204 8879 12256
rect 8879 12204 8885 12256
rect 8767 10714 8819 10724
rect 8767 10680 8773 10714
rect 8773 10680 8807 10714
rect 8807 10680 8819 10714
rect 8767 10672 8819 10680
rect 8833 10714 8885 10724
rect 8833 10680 8845 10714
rect 8845 10680 8879 10714
rect 8879 10680 8885 10714
rect 8833 10672 8885 10680
rect 8767 10641 8819 10658
rect 8767 10607 8773 10641
rect 8773 10607 8807 10641
rect 8807 10607 8819 10641
rect 8767 10606 8819 10607
rect 8833 10641 8885 10658
rect 8833 10607 8845 10641
rect 8845 10607 8879 10641
rect 8879 10607 8885 10641
rect 8833 10606 8885 10607
rect 8767 10568 8819 10592
rect 8767 10540 8773 10568
rect 8773 10540 8807 10568
rect 8807 10540 8819 10568
rect 8833 10568 8885 10592
rect 8833 10540 8845 10568
rect 8845 10540 8879 10568
rect 8879 10540 8885 10568
rect 8767 10495 8819 10526
rect 8767 10474 8773 10495
rect 8773 10474 8807 10495
rect 8807 10474 8819 10495
rect 8833 10495 8885 10526
rect 8833 10474 8845 10495
rect 8845 10474 8879 10495
rect 8879 10474 8885 10495
rect 8767 10422 8819 10460
rect 8833 10422 8885 10460
rect 8767 10408 8773 10422
rect 8773 10408 8819 10422
rect 8833 10408 8879 10422
rect 8879 10408 8885 10422
rect 8767 10342 8773 10394
rect 8773 10342 8819 10394
rect 8833 10342 8879 10394
rect 8879 10342 8885 10394
rect 8767 10275 8773 10327
rect 8773 10275 8819 10327
rect 8833 10275 8879 10327
rect 8879 10275 8885 10327
rect 8767 10208 8773 10260
rect 8773 10208 8819 10260
rect 8833 10208 8879 10260
rect 8879 10208 8885 10260
rect 8767 8714 8819 8720
rect 8767 8680 8773 8714
rect 8773 8680 8807 8714
rect 8807 8680 8819 8714
rect 8767 8668 8819 8680
rect 8833 8714 8885 8720
rect 8833 8680 8845 8714
rect 8845 8680 8879 8714
rect 8879 8680 8885 8714
rect 8833 8668 8885 8680
rect 8767 8641 8819 8654
rect 8767 8607 8773 8641
rect 8773 8607 8807 8641
rect 8807 8607 8819 8641
rect 8767 8602 8819 8607
rect 8833 8641 8885 8654
rect 8833 8607 8845 8641
rect 8845 8607 8879 8641
rect 8879 8607 8885 8641
rect 8833 8602 8885 8607
rect 8767 8568 8819 8588
rect 8767 8536 8773 8568
rect 8773 8536 8807 8568
rect 8807 8536 8819 8568
rect 8833 8568 8885 8588
rect 8833 8536 8845 8568
rect 8845 8536 8879 8568
rect 8879 8536 8885 8568
rect 8767 8495 8819 8522
rect 8767 8470 8773 8495
rect 8773 8470 8807 8495
rect 8807 8470 8819 8495
rect 8833 8495 8885 8522
rect 8833 8470 8845 8495
rect 8845 8470 8879 8495
rect 8879 8470 8885 8495
rect 8767 8422 8819 8456
rect 8833 8422 8885 8456
rect 8767 8404 8773 8422
rect 8773 8404 8819 8422
rect 8833 8404 8879 8422
rect 8879 8404 8885 8422
rect 8767 8338 8773 8390
rect 8773 8338 8819 8390
rect 8833 8338 8879 8390
rect 8879 8338 8885 8390
rect 8767 8271 8773 8323
rect 8773 8271 8819 8323
rect 8833 8271 8879 8323
rect 8879 8271 8885 8323
rect 8767 8204 8773 8256
rect 8773 8204 8819 8256
rect 8833 8204 8879 8256
rect 8879 8204 8885 8256
rect 8767 6714 8819 6724
rect 8767 6680 8773 6714
rect 8773 6680 8807 6714
rect 8807 6680 8819 6714
rect 8767 6672 8819 6680
rect 8833 6714 8885 6724
rect 8833 6680 8845 6714
rect 8845 6680 8879 6714
rect 8879 6680 8885 6714
rect 8833 6672 8885 6680
rect 8767 6641 8819 6658
rect 8767 6607 8773 6641
rect 8773 6607 8807 6641
rect 8807 6607 8819 6641
rect 8767 6606 8819 6607
rect 8833 6641 8885 6658
rect 8833 6607 8845 6641
rect 8845 6607 8879 6641
rect 8879 6607 8885 6641
rect 8833 6606 8885 6607
rect 8767 6568 8819 6592
rect 8767 6540 8773 6568
rect 8773 6540 8807 6568
rect 8807 6540 8819 6568
rect 8833 6568 8885 6592
rect 8833 6540 8845 6568
rect 8845 6540 8879 6568
rect 8879 6540 8885 6568
rect 8767 6495 8819 6526
rect 8767 6474 8773 6495
rect 8773 6474 8807 6495
rect 8807 6474 8819 6495
rect 8833 6495 8885 6526
rect 8833 6474 8845 6495
rect 8845 6474 8879 6495
rect 8879 6474 8885 6495
rect 8767 6422 8819 6460
rect 8833 6422 8885 6460
rect 8767 6408 8773 6422
rect 8773 6408 8819 6422
rect 8833 6408 8879 6422
rect 8879 6408 8885 6422
rect 8767 6342 8773 6394
rect 8773 6342 8819 6394
rect 8833 6342 8879 6394
rect 8879 6342 8885 6394
rect 8767 6275 8773 6327
rect 8773 6275 8819 6327
rect 8833 6275 8879 6327
rect 8879 6275 8885 6327
rect 8767 6208 8773 6260
rect 8773 6208 8819 6260
rect 8833 6208 8879 6260
rect 8879 6208 8885 6260
rect 9044 13877 9096 13892
rect 9044 13843 9050 13877
rect 9050 13843 9084 13877
rect 9084 13843 9096 13877
rect 9044 13840 9096 13843
rect 9110 13877 9162 13892
rect 9110 13843 9122 13877
rect 9122 13843 9156 13877
rect 9156 13843 9162 13877
rect 9110 13840 9162 13843
rect 9044 13799 9096 13826
rect 9044 13774 9050 13799
rect 9050 13774 9084 13799
rect 9084 13774 9096 13799
rect 9110 13799 9162 13826
rect 9110 13774 9122 13799
rect 9122 13774 9156 13799
rect 9156 13774 9162 13799
rect 9044 13722 9096 13760
rect 9044 13708 9050 13722
rect 9050 13708 9084 13722
rect 9084 13708 9096 13722
rect 9110 13722 9162 13760
rect 9110 13708 9122 13722
rect 9122 13708 9156 13722
rect 9156 13708 9162 13722
rect 9044 13688 9050 13694
rect 9050 13688 9084 13694
rect 9084 13688 9096 13694
rect 9044 13645 9096 13688
rect 9044 13642 9050 13645
rect 9050 13642 9084 13645
rect 9084 13642 9096 13645
rect 9110 13688 9122 13694
rect 9122 13688 9156 13694
rect 9156 13688 9162 13694
rect 9110 13645 9162 13688
rect 9110 13642 9122 13645
rect 9122 13642 9156 13645
rect 9156 13642 9162 13645
rect 9044 13611 9050 13628
rect 9050 13611 9084 13628
rect 9084 13611 9096 13628
rect 9044 13576 9096 13611
rect 9110 13611 9122 13628
rect 9122 13611 9156 13628
rect 9156 13611 9162 13628
rect 9110 13576 9162 13611
rect 9044 13534 9050 13562
rect 9050 13534 9084 13562
rect 9084 13534 9096 13562
rect 9044 13510 9096 13534
rect 9110 13534 9122 13562
rect 9122 13534 9156 13562
rect 9156 13534 9162 13562
rect 9110 13510 9162 13534
rect 9044 13491 9096 13495
rect 9044 13457 9050 13491
rect 9050 13457 9084 13491
rect 9084 13457 9096 13491
rect 9044 13443 9096 13457
rect 9110 13491 9162 13495
rect 9110 13457 9122 13491
rect 9122 13457 9156 13491
rect 9156 13457 9162 13491
rect 9110 13443 9162 13457
rect 9044 13414 9096 13428
rect 9044 13380 9050 13414
rect 9050 13380 9084 13414
rect 9084 13380 9096 13414
rect 9044 13376 9096 13380
rect 9110 13414 9162 13428
rect 9110 13380 9122 13414
rect 9122 13380 9156 13414
rect 9156 13380 9162 13414
rect 9110 13376 9162 13380
rect 9044 11840 9050 11892
rect 9050 11840 9096 11892
rect 9110 11840 9156 11892
rect 9156 11840 9162 11892
rect 9044 11774 9050 11826
rect 9050 11774 9096 11826
rect 9110 11774 9156 11826
rect 9156 11774 9162 11826
rect 9044 11708 9050 11760
rect 9050 11708 9096 11760
rect 9110 11708 9156 11760
rect 9156 11708 9162 11760
rect 9044 11642 9050 11694
rect 9050 11642 9096 11694
rect 9110 11642 9156 11694
rect 9156 11642 9162 11694
rect 9044 11576 9050 11628
rect 9050 11576 9096 11628
rect 9110 11576 9156 11628
rect 9156 11576 9162 11628
rect 9044 11510 9050 11562
rect 9050 11510 9096 11562
rect 9110 11510 9156 11562
rect 9156 11510 9162 11562
rect 9044 11443 9050 11495
rect 9050 11443 9096 11495
rect 9110 11443 9156 11495
rect 9156 11443 9162 11495
rect 9044 11380 9050 11428
rect 9050 11380 9096 11428
rect 9110 11380 9156 11428
rect 9156 11380 9162 11428
rect 9044 11376 9096 11380
rect 9110 11376 9162 11380
rect 9044 9844 9050 9896
rect 9050 9844 9096 9896
rect 9110 9844 9156 9896
rect 9156 9844 9162 9896
rect 9044 9778 9050 9830
rect 9050 9778 9096 9830
rect 9110 9778 9156 9830
rect 9156 9778 9162 9830
rect 9044 9712 9050 9764
rect 9050 9712 9096 9764
rect 9110 9712 9156 9764
rect 9156 9712 9162 9764
rect 9044 9646 9050 9698
rect 9050 9646 9096 9698
rect 9110 9646 9156 9698
rect 9156 9646 9162 9698
rect 9044 9580 9050 9632
rect 9050 9580 9096 9632
rect 9110 9580 9156 9632
rect 9156 9580 9162 9632
rect 9044 9514 9050 9566
rect 9050 9514 9096 9566
rect 9110 9514 9156 9566
rect 9156 9514 9162 9566
rect 9044 9447 9050 9499
rect 9050 9447 9096 9499
rect 9110 9447 9156 9499
rect 9156 9447 9162 9499
rect 9044 9380 9050 9432
rect 9050 9380 9096 9432
rect 9110 9380 9156 9432
rect 9156 9380 9162 9432
rect 9044 7840 9050 7892
rect 9050 7840 9096 7892
rect 9110 7840 9156 7892
rect 9156 7840 9162 7892
rect 9044 7774 9050 7826
rect 9050 7774 9096 7826
rect 9110 7774 9156 7826
rect 9156 7774 9162 7826
rect 9044 7708 9050 7760
rect 9050 7708 9096 7760
rect 9110 7708 9156 7760
rect 9156 7708 9162 7760
rect 9044 7642 9050 7694
rect 9050 7642 9096 7694
rect 9110 7642 9156 7694
rect 9156 7642 9162 7694
rect 9044 7576 9050 7628
rect 9050 7576 9096 7628
rect 9110 7576 9156 7628
rect 9156 7576 9162 7628
rect 9044 7510 9050 7562
rect 9050 7510 9096 7562
rect 9110 7510 9156 7562
rect 9156 7510 9162 7562
rect 9044 7443 9050 7495
rect 9050 7443 9096 7495
rect 9110 7443 9156 7495
rect 9156 7443 9162 7495
rect 9044 7380 9050 7428
rect 9050 7380 9096 7428
rect 9110 7380 9156 7428
rect 9156 7380 9162 7428
rect 9044 7376 9096 7380
rect 9110 7376 9162 7380
rect 9044 5844 9050 5896
rect 9050 5844 9096 5896
rect 9110 5844 9156 5896
rect 9156 5844 9162 5896
rect 9044 5778 9050 5830
rect 9050 5778 9096 5830
rect 9110 5778 9156 5830
rect 9156 5778 9162 5830
rect 9044 5712 9050 5764
rect 9050 5712 9096 5764
rect 9110 5712 9156 5764
rect 9156 5712 9162 5764
rect 9044 5646 9050 5698
rect 9050 5646 9096 5698
rect 9110 5646 9156 5698
rect 9156 5646 9162 5698
rect 9044 5580 9050 5632
rect 9050 5580 9096 5632
rect 9110 5580 9156 5632
rect 9156 5580 9162 5632
rect 9044 5514 9050 5566
rect 9050 5514 9096 5566
rect 9110 5514 9156 5566
rect 9156 5514 9162 5566
rect 9044 5447 9050 5499
rect 9050 5447 9096 5499
rect 9110 5447 9156 5499
rect 9156 5447 9162 5499
rect 9044 5380 9050 5432
rect 9050 5380 9096 5432
rect 9110 5380 9156 5432
rect 9156 5380 9162 5432
rect 9321 14345 9373 14390
rect 9321 14338 9327 14345
rect 9327 14338 9361 14345
rect 9361 14338 9373 14345
rect 9387 14345 9439 14390
rect 9875 14668 9927 14720
rect 9941 14668 9993 14720
rect 9875 14602 9927 14654
rect 9941 14602 9993 14654
rect 9875 14536 9927 14588
rect 9941 14536 9993 14588
rect 9875 14470 9927 14522
rect 9941 14470 9993 14522
rect 9875 14404 9927 14456
rect 9941 14404 9993 14456
rect 9387 14338 9399 14345
rect 9399 14338 9433 14345
rect 9433 14338 9439 14345
rect 9321 14311 9327 14323
rect 9327 14311 9361 14323
rect 9361 14311 9373 14323
rect 9321 14271 9373 14311
rect 9387 14311 9399 14323
rect 9399 14311 9433 14323
rect 9433 14311 9439 14323
rect 9387 14271 9439 14311
rect 9321 14233 9327 14256
rect 9327 14233 9361 14256
rect 9361 14233 9373 14256
rect 9321 14204 9373 14233
rect 9387 14233 9399 14256
rect 9399 14233 9433 14256
rect 9433 14233 9439 14256
rect 9387 14204 9439 14233
rect 9321 12714 9373 12720
rect 9321 12680 9327 12714
rect 9327 12680 9361 12714
rect 9361 12680 9373 12714
rect 9321 12668 9373 12680
rect 9387 12714 9439 12720
rect 9387 12680 9399 12714
rect 9399 12680 9433 12714
rect 9433 12680 9439 12714
rect 9387 12668 9439 12680
rect 9321 12641 9373 12654
rect 9321 12607 9327 12641
rect 9327 12607 9361 12641
rect 9361 12607 9373 12641
rect 9321 12602 9373 12607
rect 9387 12641 9439 12654
rect 9387 12607 9399 12641
rect 9399 12607 9433 12641
rect 9433 12607 9439 12641
rect 9387 12602 9439 12607
rect 9321 12568 9373 12588
rect 9321 12536 9327 12568
rect 9327 12536 9361 12568
rect 9361 12536 9373 12568
rect 9387 12568 9439 12588
rect 9387 12536 9399 12568
rect 9399 12536 9433 12568
rect 9433 12536 9439 12568
rect 9321 12495 9373 12522
rect 9321 12470 9327 12495
rect 9327 12470 9361 12495
rect 9361 12470 9373 12495
rect 9387 12495 9439 12522
rect 9387 12470 9399 12495
rect 9399 12470 9433 12495
rect 9433 12470 9439 12495
rect 9321 12422 9373 12456
rect 9387 12422 9439 12456
rect 9321 12404 9327 12422
rect 9327 12404 9373 12422
rect 9387 12404 9433 12422
rect 9433 12404 9439 12422
rect 9321 12338 9327 12390
rect 9327 12338 9373 12390
rect 9387 12338 9433 12390
rect 9433 12338 9439 12390
rect 9321 12271 9327 12323
rect 9327 12271 9373 12323
rect 9387 12271 9433 12323
rect 9433 12271 9439 12323
rect 9321 12204 9327 12256
rect 9327 12204 9373 12256
rect 9387 12204 9433 12256
rect 9433 12204 9439 12256
rect 9321 10714 9373 10724
rect 9321 10680 9327 10714
rect 9327 10680 9361 10714
rect 9361 10680 9373 10714
rect 9321 10672 9373 10680
rect 9387 10714 9439 10724
rect 9387 10680 9399 10714
rect 9399 10680 9433 10714
rect 9433 10680 9439 10714
rect 9387 10672 9439 10680
rect 9321 10641 9373 10658
rect 9321 10607 9327 10641
rect 9327 10607 9361 10641
rect 9361 10607 9373 10641
rect 9321 10606 9373 10607
rect 9387 10641 9439 10658
rect 9387 10607 9399 10641
rect 9399 10607 9433 10641
rect 9433 10607 9439 10641
rect 9387 10606 9439 10607
rect 9321 10568 9373 10592
rect 9321 10540 9327 10568
rect 9327 10540 9361 10568
rect 9361 10540 9373 10568
rect 9387 10568 9439 10592
rect 9387 10540 9399 10568
rect 9399 10540 9433 10568
rect 9433 10540 9439 10568
rect 9321 10495 9373 10526
rect 9321 10474 9327 10495
rect 9327 10474 9361 10495
rect 9361 10474 9373 10495
rect 9387 10495 9439 10526
rect 9387 10474 9399 10495
rect 9399 10474 9433 10495
rect 9433 10474 9439 10495
rect 9321 10422 9373 10460
rect 9387 10422 9439 10460
rect 9321 10408 9327 10422
rect 9327 10408 9373 10422
rect 9387 10408 9433 10422
rect 9433 10408 9439 10422
rect 9321 10342 9327 10394
rect 9327 10342 9373 10394
rect 9387 10342 9433 10394
rect 9433 10342 9439 10394
rect 9321 10275 9327 10327
rect 9327 10275 9373 10327
rect 9387 10275 9433 10327
rect 9433 10275 9439 10327
rect 9321 10208 9327 10260
rect 9327 10208 9373 10260
rect 9387 10208 9433 10260
rect 9433 10208 9439 10260
rect 9321 8714 9373 8720
rect 9321 8680 9327 8714
rect 9327 8680 9361 8714
rect 9361 8680 9373 8714
rect 9321 8668 9373 8680
rect 9387 8714 9439 8720
rect 9387 8680 9399 8714
rect 9399 8680 9433 8714
rect 9433 8680 9439 8714
rect 9387 8668 9439 8680
rect 9321 8641 9373 8654
rect 9321 8607 9327 8641
rect 9327 8607 9361 8641
rect 9361 8607 9373 8641
rect 9321 8602 9373 8607
rect 9387 8641 9439 8654
rect 9387 8607 9399 8641
rect 9399 8607 9433 8641
rect 9433 8607 9439 8641
rect 9387 8602 9439 8607
rect 9321 8568 9373 8588
rect 9321 8536 9327 8568
rect 9327 8536 9361 8568
rect 9361 8536 9373 8568
rect 9387 8568 9439 8588
rect 9387 8536 9399 8568
rect 9399 8536 9433 8568
rect 9433 8536 9439 8568
rect 9321 8495 9373 8522
rect 9321 8470 9327 8495
rect 9327 8470 9361 8495
rect 9361 8470 9373 8495
rect 9387 8495 9439 8522
rect 9387 8470 9399 8495
rect 9399 8470 9433 8495
rect 9433 8470 9439 8495
rect 9321 8422 9373 8456
rect 9387 8422 9439 8456
rect 9321 8404 9327 8422
rect 9327 8404 9373 8422
rect 9387 8404 9433 8422
rect 9433 8404 9439 8422
rect 9321 8338 9327 8390
rect 9327 8338 9373 8390
rect 9387 8338 9433 8390
rect 9433 8338 9439 8390
rect 9321 8271 9327 8323
rect 9327 8271 9373 8323
rect 9387 8271 9433 8323
rect 9433 8271 9439 8323
rect 9321 8204 9327 8256
rect 9327 8204 9373 8256
rect 9387 8204 9433 8256
rect 9433 8204 9439 8256
rect 9321 6714 9373 6724
rect 9321 6680 9327 6714
rect 9327 6680 9361 6714
rect 9361 6680 9373 6714
rect 9321 6672 9373 6680
rect 9387 6714 9439 6724
rect 9387 6680 9399 6714
rect 9399 6680 9433 6714
rect 9433 6680 9439 6714
rect 9387 6672 9439 6680
rect 9321 6641 9373 6658
rect 9321 6607 9327 6641
rect 9327 6607 9361 6641
rect 9361 6607 9373 6641
rect 9321 6606 9373 6607
rect 9387 6641 9439 6658
rect 9387 6607 9399 6641
rect 9399 6607 9433 6641
rect 9433 6607 9439 6641
rect 9387 6606 9439 6607
rect 9321 6568 9373 6592
rect 9321 6540 9327 6568
rect 9327 6540 9361 6568
rect 9361 6540 9373 6568
rect 9387 6568 9439 6592
rect 9387 6540 9399 6568
rect 9399 6540 9433 6568
rect 9433 6540 9439 6568
rect 9321 6495 9373 6526
rect 9321 6474 9327 6495
rect 9327 6474 9361 6495
rect 9361 6474 9373 6495
rect 9387 6495 9439 6526
rect 9387 6474 9399 6495
rect 9399 6474 9433 6495
rect 9433 6474 9439 6495
rect 9321 6422 9373 6460
rect 9387 6422 9439 6460
rect 9321 6408 9327 6422
rect 9327 6408 9373 6422
rect 9387 6408 9433 6422
rect 9433 6408 9439 6422
rect 9321 6342 9327 6394
rect 9327 6342 9373 6394
rect 9387 6342 9433 6394
rect 9433 6342 9439 6394
rect 9321 6275 9327 6327
rect 9327 6275 9373 6327
rect 9387 6275 9433 6327
rect 9433 6275 9439 6327
rect 9321 6208 9327 6260
rect 9327 6208 9373 6260
rect 9387 6208 9433 6260
rect 9433 6208 9439 6260
rect 9598 13877 9650 13892
rect 9598 13843 9604 13877
rect 9604 13843 9638 13877
rect 9638 13843 9650 13877
rect 9598 13840 9650 13843
rect 9664 13877 9716 13892
rect 9664 13843 9676 13877
rect 9676 13843 9710 13877
rect 9710 13843 9716 13877
rect 9664 13840 9716 13843
rect 9598 13799 9650 13826
rect 9598 13774 9604 13799
rect 9604 13774 9638 13799
rect 9638 13774 9650 13799
rect 9664 13799 9716 13826
rect 9664 13774 9676 13799
rect 9676 13774 9710 13799
rect 9710 13774 9716 13799
rect 9598 13722 9650 13760
rect 9598 13708 9604 13722
rect 9604 13708 9638 13722
rect 9638 13708 9650 13722
rect 9664 13722 9716 13760
rect 9664 13708 9676 13722
rect 9676 13708 9710 13722
rect 9710 13708 9716 13722
rect 9598 13688 9604 13694
rect 9604 13688 9638 13694
rect 9638 13688 9650 13694
rect 9598 13645 9650 13688
rect 9598 13642 9604 13645
rect 9604 13642 9638 13645
rect 9638 13642 9650 13645
rect 9664 13688 9676 13694
rect 9676 13688 9710 13694
rect 9710 13688 9716 13694
rect 9664 13645 9716 13688
rect 9664 13642 9676 13645
rect 9676 13642 9710 13645
rect 9710 13642 9716 13645
rect 9598 13611 9604 13628
rect 9604 13611 9638 13628
rect 9638 13611 9650 13628
rect 9598 13576 9650 13611
rect 9664 13611 9676 13628
rect 9676 13611 9710 13628
rect 9710 13611 9716 13628
rect 9664 13576 9716 13611
rect 9598 13534 9604 13562
rect 9604 13534 9638 13562
rect 9638 13534 9650 13562
rect 9598 13510 9650 13534
rect 9664 13534 9676 13562
rect 9676 13534 9710 13562
rect 9710 13534 9716 13562
rect 9664 13510 9716 13534
rect 9598 13491 9650 13495
rect 9598 13457 9604 13491
rect 9604 13457 9638 13491
rect 9638 13457 9650 13491
rect 9598 13443 9650 13457
rect 9664 13491 9716 13495
rect 9664 13457 9676 13491
rect 9676 13457 9710 13491
rect 9710 13457 9716 13491
rect 9664 13443 9716 13457
rect 9598 13414 9650 13428
rect 9598 13380 9604 13414
rect 9604 13380 9638 13414
rect 9638 13380 9650 13414
rect 9598 13376 9650 13380
rect 9664 13414 9716 13428
rect 9664 13380 9676 13414
rect 9676 13380 9710 13414
rect 9710 13380 9716 13414
rect 9664 13376 9716 13380
rect 9598 11840 9604 11892
rect 9604 11840 9650 11892
rect 9664 11840 9710 11892
rect 9710 11840 9716 11892
rect 9598 11774 9604 11826
rect 9604 11774 9650 11826
rect 9664 11774 9710 11826
rect 9710 11774 9716 11826
rect 9598 11708 9604 11760
rect 9604 11708 9650 11760
rect 9664 11708 9710 11760
rect 9710 11708 9716 11760
rect 9598 11642 9604 11694
rect 9604 11642 9650 11694
rect 9664 11642 9710 11694
rect 9710 11642 9716 11694
rect 9598 11576 9604 11628
rect 9604 11576 9650 11628
rect 9664 11576 9710 11628
rect 9710 11576 9716 11628
rect 9598 11510 9604 11562
rect 9604 11510 9650 11562
rect 9664 11510 9710 11562
rect 9710 11510 9716 11562
rect 9598 11443 9604 11495
rect 9604 11443 9650 11495
rect 9664 11443 9710 11495
rect 9710 11443 9716 11495
rect 9598 11380 9604 11428
rect 9604 11380 9650 11428
rect 9664 11380 9710 11428
rect 9710 11380 9716 11428
rect 9598 11376 9650 11380
rect 9664 11376 9716 11380
rect 9598 9844 9604 9896
rect 9604 9844 9650 9896
rect 9664 9844 9710 9896
rect 9710 9844 9716 9896
rect 9598 9778 9604 9830
rect 9604 9778 9650 9830
rect 9664 9778 9710 9830
rect 9710 9778 9716 9830
rect 9598 9712 9604 9764
rect 9604 9712 9650 9764
rect 9664 9712 9710 9764
rect 9710 9712 9716 9764
rect 9598 9646 9604 9698
rect 9604 9646 9650 9698
rect 9664 9646 9710 9698
rect 9710 9646 9716 9698
rect 9598 9580 9604 9632
rect 9604 9580 9650 9632
rect 9664 9580 9710 9632
rect 9710 9580 9716 9632
rect 9598 9514 9604 9566
rect 9604 9514 9650 9566
rect 9664 9514 9710 9566
rect 9710 9514 9716 9566
rect 9598 9447 9604 9499
rect 9604 9447 9650 9499
rect 9664 9447 9710 9499
rect 9710 9447 9716 9499
rect 9598 9380 9604 9432
rect 9604 9380 9650 9432
rect 9664 9380 9710 9432
rect 9710 9380 9716 9432
rect 9598 7840 9604 7892
rect 9604 7840 9650 7892
rect 9664 7840 9710 7892
rect 9710 7840 9716 7892
rect 9598 7774 9604 7826
rect 9604 7774 9650 7826
rect 9664 7774 9710 7826
rect 9710 7774 9716 7826
rect 9598 7708 9604 7760
rect 9604 7708 9650 7760
rect 9664 7708 9710 7760
rect 9710 7708 9716 7760
rect 9598 7642 9604 7694
rect 9604 7642 9650 7694
rect 9664 7642 9710 7694
rect 9710 7642 9716 7694
rect 9598 7576 9604 7628
rect 9604 7576 9650 7628
rect 9664 7576 9710 7628
rect 9710 7576 9716 7628
rect 9598 7510 9604 7562
rect 9604 7510 9650 7562
rect 9664 7510 9710 7562
rect 9710 7510 9716 7562
rect 9598 7443 9604 7495
rect 9604 7443 9650 7495
rect 9664 7443 9710 7495
rect 9710 7443 9716 7495
rect 9598 7380 9604 7428
rect 9604 7380 9650 7428
rect 9664 7380 9710 7428
rect 9710 7380 9716 7428
rect 9598 7376 9650 7380
rect 9664 7376 9716 7380
rect 9598 5844 9604 5896
rect 9604 5844 9650 5896
rect 9664 5844 9710 5896
rect 9710 5844 9716 5896
rect 9598 5778 9604 5830
rect 9604 5778 9650 5830
rect 9664 5778 9710 5830
rect 9710 5778 9716 5830
rect 9598 5712 9604 5764
rect 9604 5712 9650 5764
rect 9664 5712 9710 5764
rect 9710 5712 9716 5764
rect 9598 5646 9604 5698
rect 9604 5646 9650 5698
rect 9664 5646 9710 5698
rect 9710 5646 9716 5698
rect 9598 5580 9604 5632
rect 9604 5580 9650 5632
rect 9664 5580 9710 5632
rect 9710 5580 9716 5632
rect 9598 5514 9604 5566
rect 9604 5514 9650 5566
rect 9664 5514 9710 5566
rect 9710 5514 9716 5566
rect 9598 5447 9604 5499
rect 9604 5447 9650 5499
rect 9664 5447 9710 5499
rect 9710 5447 9716 5499
rect 9598 5380 9604 5432
rect 9604 5380 9650 5432
rect 9664 5380 9710 5432
rect 9710 5380 9716 5432
rect 9875 14345 9927 14390
rect 9875 14338 9881 14345
rect 9881 14338 9915 14345
rect 9915 14338 9927 14345
rect 9941 14345 9993 14390
rect 10429 14668 10481 14720
rect 10495 14668 10547 14720
rect 10429 14602 10481 14654
rect 10495 14602 10547 14654
rect 10429 14536 10481 14588
rect 10495 14536 10547 14588
rect 10429 14470 10481 14522
rect 10495 14470 10547 14522
rect 10429 14404 10481 14456
rect 10495 14404 10547 14456
rect 9941 14338 9953 14345
rect 9953 14338 9987 14345
rect 9987 14338 9993 14345
rect 9875 14311 9881 14323
rect 9881 14311 9915 14323
rect 9915 14311 9927 14323
rect 9875 14271 9927 14311
rect 9941 14311 9953 14323
rect 9953 14311 9987 14323
rect 9987 14311 9993 14323
rect 9941 14271 9993 14311
rect 9875 14233 9881 14256
rect 9881 14233 9915 14256
rect 9915 14233 9927 14256
rect 9875 14204 9927 14233
rect 9941 14233 9953 14256
rect 9953 14233 9987 14256
rect 9987 14233 9993 14256
rect 9941 14204 9993 14233
rect 9875 12714 9927 12720
rect 9875 12680 9881 12714
rect 9881 12680 9915 12714
rect 9915 12680 9927 12714
rect 9875 12668 9927 12680
rect 9941 12714 9993 12720
rect 9941 12680 9953 12714
rect 9953 12680 9987 12714
rect 9987 12680 9993 12714
rect 9941 12668 9993 12680
rect 9875 12641 9927 12654
rect 9875 12607 9881 12641
rect 9881 12607 9915 12641
rect 9915 12607 9927 12641
rect 9875 12602 9927 12607
rect 9941 12641 9993 12654
rect 9941 12607 9953 12641
rect 9953 12607 9987 12641
rect 9987 12607 9993 12641
rect 9941 12602 9993 12607
rect 9875 12568 9927 12588
rect 9875 12536 9881 12568
rect 9881 12536 9915 12568
rect 9915 12536 9927 12568
rect 9941 12568 9993 12588
rect 9941 12536 9953 12568
rect 9953 12536 9987 12568
rect 9987 12536 9993 12568
rect 9875 12495 9927 12522
rect 9875 12470 9881 12495
rect 9881 12470 9915 12495
rect 9915 12470 9927 12495
rect 9941 12495 9993 12522
rect 9941 12470 9953 12495
rect 9953 12470 9987 12495
rect 9987 12470 9993 12495
rect 9875 12422 9927 12456
rect 9941 12422 9993 12456
rect 9875 12404 9881 12422
rect 9881 12404 9927 12422
rect 9941 12404 9987 12422
rect 9987 12404 9993 12422
rect 9875 12338 9881 12390
rect 9881 12338 9927 12390
rect 9941 12338 9987 12390
rect 9987 12338 9993 12390
rect 9875 12271 9881 12323
rect 9881 12271 9927 12323
rect 9941 12271 9987 12323
rect 9987 12271 9993 12323
rect 9875 12204 9881 12256
rect 9881 12204 9927 12256
rect 9941 12204 9987 12256
rect 9987 12204 9993 12256
rect 9875 10714 9927 10724
rect 9875 10680 9881 10714
rect 9881 10680 9915 10714
rect 9915 10680 9927 10714
rect 9875 10672 9927 10680
rect 9941 10714 9993 10724
rect 9941 10680 9953 10714
rect 9953 10680 9987 10714
rect 9987 10680 9993 10714
rect 9941 10672 9993 10680
rect 9875 10641 9927 10658
rect 9875 10607 9881 10641
rect 9881 10607 9915 10641
rect 9915 10607 9927 10641
rect 9875 10606 9927 10607
rect 9941 10641 9993 10658
rect 9941 10607 9953 10641
rect 9953 10607 9987 10641
rect 9987 10607 9993 10641
rect 9941 10606 9993 10607
rect 9875 10568 9927 10592
rect 9875 10540 9881 10568
rect 9881 10540 9915 10568
rect 9915 10540 9927 10568
rect 9941 10568 9993 10592
rect 9941 10540 9953 10568
rect 9953 10540 9987 10568
rect 9987 10540 9993 10568
rect 9875 10495 9927 10526
rect 9875 10474 9881 10495
rect 9881 10474 9915 10495
rect 9915 10474 9927 10495
rect 9941 10495 9993 10526
rect 9941 10474 9953 10495
rect 9953 10474 9987 10495
rect 9987 10474 9993 10495
rect 9875 10422 9927 10460
rect 9941 10422 9993 10460
rect 9875 10408 9881 10422
rect 9881 10408 9927 10422
rect 9941 10408 9987 10422
rect 9987 10408 9993 10422
rect 9875 10342 9881 10394
rect 9881 10342 9927 10394
rect 9941 10342 9987 10394
rect 9987 10342 9993 10394
rect 9875 10275 9881 10327
rect 9881 10275 9927 10327
rect 9941 10275 9987 10327
rect 9987 10275 9993 10327
rect 9875 10208 9881 10260
rect 9881 10208 9927 10260
rect 9941 10208 9987 10260
rect 9987 10208 9993 10260
rect 9875 8714 9927 8720
rect 9875 8680 9881 8714
rect 9881 8680 9915 8714
rect 9915 8680 9927 8714
rect 9875 8668 9927 8680
rect 9941 8714 9993 8720
rect 9941 8680 9953 8714
rect 9953 8680 9987 8714
rect 9987 8680 9993 8714
rect 9941 8668 9993 8680
rect 9875 8641 9927 8654
rect 9875 8607 9881 8641
rect 9881 8607 9915 8641
rect 9915 8607 9927 8641
rect 9875 8602 9927 8607
rect 9941 8641 9993 8654
rect 9941 8607 9953 8641
rect 9953 8607 9987 8641
rect 9987 8607 9993 8641
rect 9941 8602 9993 8607
rect 9875 8568 9927 8588
rect 9875 8536 9881 8568
rect 9881 8536 9915 8568
rect 9915 8536 9927 8568
rect 9941 8568 9993 8588
rect 9941 8536 9953 8568
rect 9953 8536 9987 8568
rect 9987 8536 9993 8568
rect 9875 8495 9927 8522
rect 9875 8470 9881 8495
rect 9881 8470 9915 8495
rect 9915 8470 9927 8495
rect 9941 8495 9993 8522
rect 9941 8470 9953 8495
rect 9953 8470 9987 8495
rect 9987 8470 9993 8495
rect 9875 8422 9927 8456
rect 9941 8422 9993 8456
rect 9875 8404 9881 8422
rect 9881 8404 9927 8422
rect 9941 8404 9987 8422
rect 9987 8404 9993 8422
rect 9875 8338 9881 8390
rect 9881 8338 9927 8390
rect 9941 8338 9987 8390
rect 9987 8338 9993 8390
rect 9875 8271 9881 8323
rect 9881 8271 9927 8323
rect 9941 8271 9987 8323
rect 9987 8271 9993 8323
rect 9875 8204 9881 8256
rect 9881 8204 9927 8256
rect 9941 8204 9987 8256
rect 9987 8204 9993 8256
rect 9875 6714 9927 6724
rect 9875 6680 9881 6714
rect 9881 6680 9915 6714
rect 9915 6680 9927 6714
rect 9875 6672 9927 6680
rect 9941 6714 9993 6724
rect 9941 6680 9953 6714
rect 9953 6680 9987 6714
rect 9987 6680 9993 6714
rect 9941 6672 9993 6680
rect 9875 6641 9927 6658
rect 9875 6607 9881 6641
rect 9881 6607 9915 6641
rect 9915 6607 9927 6641
rect 9875 6606 9927 6607
rect 9941 6641 9993 6658
rect 9941 6607 9953 6641
rect 9953 6607 9987 6641
rect 9987 6607 9993 6641
rect 9941 6606 9993 6607
rect 9875 6568 9927 6592
rect 9875 6540 9881 6568
rect 9881 6540 9915 6568
rect 9915 6540 9927 6568
rect 9941 6568 9993 6592
rect 9941 6540 9953 6568
rect 9953 6540 9987 6568
rect 9987 6540 9993 6568
rect 9875 6495 9927 6526
rect 9875 6474 9881 6495
rect 9881 6474 9915 6495
rect 9915 6474 9927 6495
rect 9941 6495 9993 6526
rect 9941 6474 9953 6495
rect 9953 6474 9987 6495
rect 9987 6474 9993 6495
rect 9875 6422 9927 6460
rect 9941 6422 9993 6460
rect 9875 6408 9881 6422
rect 9881 6408 9927 6422
rect 9941 6408 9987 6422
rect 9987 6408 9993 6422
rect 9875 6342 9881 6394
rect 9881 6342 9927 6394
rect 9941 6342 9987 6394
rect 9987 6342 9993 6394
rect 9875 6275 9881 6327
rect 9881 6275 9927 6327
rect 9941 6275 9987 6327
rect 9987 6275 9993 6327
rect 9875 6208 9881 6260
rect 9881 6208 9927 6260
rect 9941 6208 9987 6260
rect 9987 6208 9993 6260
rect 10152 13877 10204 13892
rect 10152 13843 10158 13877
rect 10158 13843 10192 13877
rect 10192 13843 10204 13877
rect 10152 13840 10204 13843
rect 10218 13877 10270 13892
rect 10218 13843 10230 13877
rect 10230 13843 10264 13877
rect 10264 13843 10270 13877
rect 10218 13840 10270 13843
rect 10152 13799 10204 13826
rect 10152 13774 10158 13799
rect 10158 13774 10192 13799
rect 10192 13774 10204 13799
rect 10218 13799 10270 13826
rect 10218 13774 10230 13799
rect 10230 13774 10264 13799
rect 10264 13774 10270 13799
rect 10152 13722 10204 13760
rect 10152 13708 10158 13722
rect 10158 13708 10192 13722
rect 10192 13708 10204 13722
rect 10218 13722 10270 13760
rect 10218 13708 10230 13722
rect 10230 13708 10264 13722
rect 10264 13708 10270 13722
rect 10152 13688 10158 13694
rect 10158 13688 10192 13694
rect 10192 13688 10204 13694
rect 10152 13645 10204 13688
rect 10152 13642 10158 13645
rect 10158 13642 10192 13645
rect 10192 13642 10204 13645
rect 10218 13688 10230 13694
rect 10230 13688 10264 13694
rect 10264 13688 10270 13694
rect 10218 13645 10270 13688
rect 10218 13642 10230 13645
rect 10230 13642 10264 13645
rect 10264 13642 10270 13645
rect 10152 13611 10158 13628
rect 10158 13611 10192 13628
rect 10192 13611 10204 13628
rect 10152 13576 10204 13611
rect 10218 13611 10230 13628
rect 10230 13611 10264 13628
rect 10264 13611 10270 13628
rect 10218 13576 10270 13611
rect 10152 13534 10158 13562
rect 10158 13534 10192 13562
rect 10192 13534 10204 13562
rect 10152 13510 10204 13534
rect 10218 13534 10230 13562
rect 10230 13534 10264 13562
rect 10264 13534 10270 13562
rect 10218 13510 10270 13534
rect 10152 13491 10204 13495
rect 10152 13457 10158 13491
rect 10158 13457 10192 13491
rect 10192 13457 10204 13491
rect 10152 13443 10204 13457
rect 10218 13491 10270 13495
rect 10218 13457 10230 13491
rect 10230 13457 10264 13491
rect 10264 13457 10270 13491
rect 10218 13443 10270 13457
rect 10152 13414 10204 13428
rect 10152 13380 10158 13414
rect 10158 13380 10192 13414
rect 10192 13380 10204 13414
rect 10152 13376 10204 13380
rect 10218 13414 10270 13428
rect 10218 13380 10230 13414
rect 10230 13380 10264 13414
rect 10264 13380 10270 13414
rect 10218 13376 10270 13380
rect 10152 11840 10158 11892
rect 10158 11840 10204 11892
rect 10218 11840 10264 11892
rect 10264 11840 10270 11892
rect 10152 11774 10158 11826
rect 10158 11774 10204 11826
rect 10218 11774 10264 11826
rect 10264 11774 10270 11826
rect 10152 11708 10158 11760
rect 10158 11708 10204 11760
rect 10218 11708 10264 11760
rect 10264 11708 10270 11760
rect 10152 11642 10158 11694
rect 10158 11642 10204 11694
rect 10218 11642 10264 11694
rect 10264 11642 10270 11694
rect 10152 11576 10158 11628
rect 10158 11576 10204 11628
rect 10218 11576 10264 11628
rect 10264 11576 10270 11628
rect 10152 11510 10158 11562
rect 10158 11510 10204 11562
rect 10218 11510 10264 11562
rect 10264 11510 10270 11562
rect 10152 11443 10158 11495
rect 10158 11443 10204 11495
rect 10218 11443 10264 11495
rect 10264 11443 10270 11495
rect 10152 11380 10158 11428
rect 10158 11380 10204 11428
rect 10218 11380 10264 11428
rect 10264 11380 10270 11428
rect 10152 11376 10204 11380
rect 10218 11376 10270 11380
rect 10152 9844 10158 9896
rect 10158 9844 10204 9896
rect 10218 9844 10264 9896
rect 10264 9844 10270 9896
rect 10152 9778 10158 9830
rect 10158 9778 10204 9830
rect 10218 9778 10264 9830
rect 10264 9778 10270 9830
rect 10152 9712 10158 9764
rect 10158 9712 10204 9764
rect 10218 9712 10264 9764
rect 10264 9712 10270 9764
rect 10152 9646 10158 9698
rect 10158 9646 10204 9698
rect 10218 9646 10264 9698
rect 10264 9646 10270 9698
rect 10152 9580 10158 9632
rect 10158 9580 10204 9632
rect 10218 9580 10264 9632
rect 10264 9580 10270 9632
rect 10152 9514 10158 9566
rect 10158 9514 10204 9566
rect 10218 9514 10264 9566
rect 10264 9514 10270 9566
rect 10152 9447 10158 9499
rect 10158 9447 10204 9499
rect 10218 9447 10264 9499
rect 10264 9447 10270 9499
rect 10152 9380 10158 9432
rect 10158 9380 10204 9432
rect 10218 9380 10264 9432
rect 10264 9380 10270 9432
rect 10152 7840 10158 7892
rect 10158 7840 10204 7892
rect 10218 7840 10264 7892
rect 10264 7840 10270 7892
rect 10152 7774 10158 7826
rect 10158 7774 10204 7826
rect 10218 7774 10264 7826
rect 10264 7774 10270 7826
rect 10152 7708 10158 7760
rect 10158 7708 10204 7760
rect 10218 7708 10264 7760
rect 10264 7708 10270 7760
rect 10152 7642 10158 7694
rect 10158 7642 10204 7694
rect 10218 7642 10264 7694
rect 10264 7642 10270 7694
rect 10152 7576 10158 7628
rect 10158 7576 10204 7628
rect 10218 7576 10264 7628
rect 10264 7576 10270 7628
rect 10152 7510 10158 7562
rect 10158 7510 10204 7562
rect 10218 7510 10264 7562
rect 10264 7510 10270 7562
rect 10152 7443 10158 7495
rect 10158 7443 10204 7495
rect 10218 7443 10264 7495
rect 10264 7443 10270 7495
rect 10152 7380 10158 7428
rect 10158 7380 10204 7428
rect 10218 7380 10264 7428
rect 10264 7380 10270 7428
rect 10152 7376 10204 7380
rect 10218 7376 10270 7380
rect 10152 5844 10158 5896
rect 10158 5844 10204 5896
rect 10218 5844 10264 5896
rect 10264 5844 10270 5896
rect 10152 5778 10158 5830
rect 10158 5778 10204 5830
rect 10218 5778 10264 5830
rect 10264 5778 10270 5830
rect 10152 5712 10158 5764
rect 10158 5712 10204 5764
rect 10218 5712 10264 5764
rect 10264 5712 10270 5764
rect 10152 5646 10158 5698
rect 10158 5646 10204 5698
rect 10218 5646 10264 5698
rect 10264 5646 10270 5698
rect 10152 5580 10158 5632
rect 10158 5580 10204 5632
rect 10218 5580 10264 5632
rect 10264 5580 10270 5632
rect 10152 5514 10158 5566
rect 10158 5514 10204 5566
rect 10218 5514 10264 5566
rect 10264 5514 10270 5566
rect 10152 5447 10158 5499
rect 10158 5447 10204 5499
rect 10218 5447 10264 5499
rect 10264 5447 10270 5499
rect 10152 5380 10158 5432
rect 10158 5380 10204 5432
rect 10218 5380 10264 5432
rect 10264 5380 10270 5432
rect 10429 14345 10481 14390
rect 10429 14338 10435 14345
rect 10435 14338 10469 14345
rect 10469 14338 10481 14345
rect 10495 14345 10547 14390
rect 10983 14668 11035 14720
rect 11049 14668 11101 14720
rect 10983 14602 11035 14654
rect 11049 14602 11101 14654
rect 10983 14536 11035 14588
rect 11049 14536 11101 14588
rect 10983 14470 11035 14522
rect 11049 14470 11101 14522
rect 10983 14404 11035 14456
rect 11049 14404 11101 14456
rect 10495 14338 10507 14345
rect 10507 14338 10541 14345
rect 10541 14338 10547 14345
rect 10429 14311 10435 14323
rect 10435 14311 10469 14323
rect 10469 14311 10481 14323
rect 10429 14271 10481 14311
rect 10495 14311 10507 14323
rect 10507 14311 10541 14323
rect 10541 14311 10547 14323
rect 10495 14271 10547 14311
rect 10429 14233 10435 14256
rect 10435 14233 10469 14256
rect 10469 14233 10481 14256
rect 10429 14204 10481 14233
rect 10495 14233 10507 14256
rect 10507 14233 10541 14256
rect 10541 14233 10547 14256
rect 10495 14204 10547 14233
rect 10429 12714 10481 12720
rect 10429 12680 10435 12714
rect 10435 12680 10469 12714
rect 10469 12680 10481 12714
rect 10429 12668 10481 12680
rect 10495 12714 10547 12720
rect 10495 12680 10507 12714
rect 10507 12680 10541 12714
rect 10541 12680 10547 12714
rect 10495 12668 10547 12680
rect 10429 12641 10481 12654
rect 10429 12607 10435 12641
rect 10435 12607 10469 12641
rect 10469 12607 10481 12641
rect 10429 12602 10481 12607
rect 10495 12641 10547 12654
rect 10495 12607 10507 12641
rect 10507 12607 10541 12641
rect 10541 12607 10547 12641
rect 10495 12602 10547 12607
rect 10429 12568 10481 12588
rect 10429 12536 10435 12568
rect 10435 12536 10469 12568
rect 10469 12536 10481 12568
rect 10495 12568 10547 12588
rect 10495 12536 10507 12568
rect 10507 12536 10541 12568
rect 10541 12536 10547 12568
rect 10429 12495 10481 12522
rect 10429 12470 10435 12495
rect 10435 12470 10469 12495
rect 10469 12470 10481 12495
rect 10495 12495 10547 12522
rect 10495 12470 10507 12495
rect 10507 12470 10541 12495
rect 10541 12470 10547 12495
rect 10429 12422 10481 12456
rect 10495 12422 10547 12456
rect 10429 12404 10435 12422
rect 10435 12404 10481 12422
rect 10495 12404 10541 12422
rect 10541 12404 10547 12422
rect 10429 12338 10435 12390
rect 10435 12338 10481 12390
rect 10495 12338 10541 12390
rect 10541 12338 10547 12390
rect 10429 12271 10435 12323
rect 10435 12271 10481 12323
rect 10495 12271 10541 12323
rect 10541 12271 10547 12323
rect 10429 12204 10435 12256
rect 10435 12204 10481 12256
rect 10495 12204 10541 12256
rect 10541 12204 10547 12256
rect 10429 10714 10481 10724
rect 10429 10680 10435 10714
rect 10435 10680 10469 10714
rect 10469 10680 10481 10714
rect 10429 10672 10481 10680
rect 10495 10714 10547 10724
rect 10495 10680 10507 10714
rect 10507 10680 10541 10714
rect 10541 10680 10547 10714
rect 10495 10672 10547 10680
rect 10429 10641 10481 10658
rect 10429 10607 10435 10641
rect 10435 10607 10469 10641
rect 10469 10607 10481 10641
rect 10429 10606 10481 10607
rect 10495 10641 10547 10658
rect 10495 10607 10507 10641
rect 10507 10607 10541 10641
rect 10541 10607 10547 10641
rect 10495 10606 10547 10607
rect 10429 10568 10481 10592
rect 10429 10540 10435 10568
rect 10435 10540 10469 10568
rect 10469 10540 10481 10568
rect 10495 10568 10547 10592
rect 10495 10540 10507 10568
rect 10507 10540 10541 10568
rect 10541 10540 10547 10568
rect 10429 10495 10481 10526
rect 10429 10474 10435 10495
rect 10435 10474 10469 10495
rect 10469 10474 10481 10495
rect 10495 10495 10547 10526
rect 10495 10474 10507 10495
rect 10507 10474 10541 10495
rect 10541 10474 10547 10495
rect 10429 10422 10481 10460
rect 10495 10422 10547 10460
rect 10429 10408 10435 10422
rect 10435 10408 10481 10422
rect 10495 10408 10541 10422
rect 10541 10408 10547 10422
rect 10429 10342 10435 10394
rect 10435 10342 10481 10394
rect 10495 10342 10541 10394
rect 10541 10342 10547 10394
rect 10429 10275 10435 10327
rect 10435 10275 10481 10327
rect 10495 10275 10541 10327
rect 10541 10275 10547 10327
rect 10429 10208 10435 10260
rect 10435 10208 10481 10260
rect 10495 10208 10541 10260
rect 10541 10208 10547 10260
rect 10429 8714 10481 8720
rect 10429 8680 10435 8714
rect 10435 8680 10469 8714
rect 10469 8680 10481 8714
rect 10429 8668 10481 8680
rect 10495 8714 10547 8720
rect 10495 8680 10507 8714
rect 10507 8680 10541 8714
rect 10541 8680 10547 8714
rect 10495 8668 10547 8680
rect 10429 8641 10481 8654
rect 10429 8607 10435 8641
rect 10435 8607 10469 8641
rect 10469 8607 10481 8641
rect 10429 8602 10481 8607
rect 10495 8641 10547 8654
rect 10495 8607 10507 8641
rect 10507 8607 10541 8641
rect 10541 8607 10547 8641
rect 10495 8602 10547 8607
rect 10429 8568 10481 8588
rect 10429 8536 10435 8568
rect 10435 8536 10469 8568
rect 10469 8536 10481 8568
rect 10495 8568 10547 8588
rect 10495 8536 10507 8568
rect 10507 8536 10541 8568
rect 10541 8536 10547 8568
rect 10429 8495 10481 8522
rect 10429 8470 10435 8495
rect 10435 8470 10469 8495
rect 10469 8470 10481 8495
rect 10495 8495 10547 8522
rect 10495 8470 10507 8495
rect 10507 8470 10541 8495
rect 10541 8470 10547 8495
rect 10429 8422 10481 8456
rect 10495 8422 10547 8456
rect 10429 8404 10435 8422
rect 10435 8404 10481 8422
rect 10495 8404 10541 8422
rect 10541 8404 10547 8422
rect 10429 8338 10435 8390
rect 10435 8338 10481 8390
rect 10495 8338 10541 8390
rect 10541 8338 10547 8390
rect 10429 8271 10435 8323
rect 10435 8271 10481 8323
rect 10495 8271 10541 8323
rect 10541 8271 10547 8323
rect 10429 8204 10435 8256
rect 10435 8204 10481 8256
rect 10495 8204 10541 8256
rect 10541 8204 10547 8256
rect 10429 6714 10481 6724
rect 10429 6680 10435 6714
rect 10435 6680 10469 6714
rect 10469 6680 10481 6714
rect 10429 6672 10481 6680
rect 10495 6714 10547 6724
rect 10495 6680 10507 6714
rect 10507 6680 10541 6714
rect 10541 6680 10547 6714
rect 10495 6672 10547 6680
rect 10429 6641 10481 6658
rect 10429 6607 10435 6641
rect 10435 6607 10469 6641
rect 10469 6607 10481 6641
rect 10429 6606 10481 6607
rect 10495 6641 10547 6658
rect 10495 6607 10507 6641
rect 10507 6607 10541 6641
rect 10541 6607 10547 6641
rect 10495 6606 10547 6607
rect 10429 6568 10481 6592
rect 10429 6540 10435 6568
rect 10435 6540 10469 6568
rect 10469 6540 10481 6568
rect 10495 6568 10547 6592
rect 10495 6540 10507 6568
rect 10507 6540 10541 6568
rect 10541 6540 10547 6568
rect 10429 6495 10481 6526
rect 10429 6474 10435 6495
rect 10435 6474 10469 6495
rect 10469 6474 10481 6495
rect 10495 6495 10547 6526
rect 10495 6474 10507 6495
rect 10507 6474 10541 6495
rect 10541 6474 10547 6495
rect 10429 6422 10481 6460
rect 10495 6422 10547 6460
rect 10429 6408 10435 6422
rect 10435 6408 10481 6422
rect 10495 6408 10541 6422
rect 10541 6408 10547 6422
rect 10429 6342 10435 6394
rect 10435 6342 10481 6394
rect 10495 6342 10541 6394
rect 10541 6342 10547 6394
rect 10429 6275 10435 6327
rect 10435 6275 10481 6327
rect 10495 6275 10541 6327
rect 10541 6275 10547 6327
rect 10429 6208 10435 6260
rect 10435 6208 10481 6260
rect 10495 6208 10541 6260
rect 10541 6208 10547 6260
rect 10706 13877 10758 13892
rect 10706 13843 10712 13877
rect 10712 13843 10746 13877
rect 10746 13843 10758 13877
rect 10706 13840 10758 13843
rect 10772 13877 10824 13892
rect 10772 13843 10784 13877
rect 10784 13843 10818 13877
rect 10818 13843 10824 13877
rect 10772 13840 10824 13843
rect 10706 13799 10758 13826
rect 10706 13774 10712 13799
rect 10712 13774 10746 13799
rect 10746 13774 10758 13799
rect 10772 13799 10824 13826
rect 10772 13774 10784 13799
rect 10784 13774 10818 13799
rect 10818 13774 10824 13799
rect 10706 13722 10758 13760
rect 10706 13708 10712 13722
rect 10712 13708 10746 13722
rect 10746 13708 10758 13722
rect 10772 13722 10824 13760
rect 10772 13708 10784 13722
rect 10784 13708 10818 13722
rect 10818 13708 10824 13722
rect 10706 13688 10712 13694
rect 10712 13688 10746 13694
rect 10746 13688 10758 13694
rect 10706 13645 10758 13688
rect 10706 13642 10712 13645
rect 10712 13642 10746 13645
rect 10746 13642 10758 13645
rect 10772 13688 10784 13694
rect 10784 13688 10818 13694
rect 10818 13688 10824 13694
rect 10772 13645 10824 13688
rect 10772 13642 10784 13645
rect 10784 13642 10818 13645
rect 10818 13642 10824 13645
rect 10706 13611 10712 13628
rect 10712 13611 10746 13628
rect 10746 13611 10758 13628
rect 10706 13576 10758 13611
rect 10772 13611 10784 13628
rect 10784 13611 10818 13628
rect 10818 13611 10824 13628
rect 10772 13576 10824 13611
rect 10706 13534 10712 13562
rect 10712 13534 10746 13562
rect 10746 13534 10758 13562
rect 10706 13510 10758 13534
rect 10772 13534 10784 13562
rect 10784 13534 10818 13562
rect 10818 13534 10824 13562
rect 10772 13510 10824 13534
rect 10706 13491 10758 13495
rect 10706 13457 10712 13491
rect 10712 13457 10746 13491
rect 10746 13457 10758 13491
rect 10706 13443 10758 13457
rect 10772 13491 10824 13495
rect 10772 13457 10784 13491
rect 10784 13457 10818 13491
rect 10818 13457 10824 13491
rect 10772 13443 10824 13457
rect 10706 13414 10758 13428
rect 10706 13380 10712 13414
rect 10712 13380 10746 13414
rect 10746 13380 10758 13414
rect 10706 13376 10758 13380
rect 10772 13414 10824 13428
rect 10772 13380 10784 13414
rect 10784 13380 10818 13414
rect 10818 13380 10824 13414
rect 10772 13376 10824 13380
rect 10706 11840 10712 11892
rect 10712 11840 10758 11892
rect 10772 11840 10818 11892
rect 10818 11840 10824 11892
rect 10706 11774 10712 11826
rect 10712 11774 10758 11826
rect 10772 11774 10818 11826
rect 10818 11774 10824 11826
rect 10706 11708 10712 11760
rect 10712 11708 10758 11760
rect 10772 11708 10818 11760
rect 10818 11708 10824 11760
rect 10706 11642 10712 11694
rect 10712 11642 10758 11694
rect 10772 11642 10818 11694
rect 10818 11642 10824 11694
rect 10706 11576 10712 11628
rect 10712 11576 10758 11628
rect 10772 11576 10818 11628
rect 10818 11576 10824 11628
rect 10706 11510 10712 11562
rect 10712 11510 10758 11562
rect 10772 11510 10818 11562
rect 10818 11510 10824 11562
rect 10706 11443 10712 11495
rect 10712 11443 10758 11495
rect 10772 11443 10818 11495
rect 10818 11443 10824 11495
rect 10706 11380 10712 11428
rect 10712 11380 10758 11428
rect 10772 11380 10818 11428
rect 10818 11380 10824 11428
rect 10706 11376 10758 11380
rect 10772 11376 10824 11380
rect 10706 9844 10712 9896
rect 10712 9844 10758 9896
rect 10772 9844 10818 9896
rect 10818 9844 10824 9896
rect 10706 9778 10712 9830
rect 10712 9778 10758 9830
rect 10772 9778 10818 9830
rect 10818 9778 10824 9830
rect 10706 9712 10712 9764
rect 10712 9712 10758 9764
rect 10772 9712 10818 9764
rect 10818 9712 10824 9764
rect 10706 9646 10712 9698
rect 10712 9646 10758 9698
rect 10772 9646 10818 9698
rect 10818 9646 10824 9698
rect 10706 9580 10712 9632
rect 10712 9580 10758 9632
rect 10772 9580 10818 9632
rect 10818 9580 10824 9632
rect 10706 9514 10712 9566
rect 10712 9514 10758 9566
rect 10772 9514 10818 9566
rect 10818 9514 10824 9566
rect 10706 9447 10712 9499
rect 10712 9447 10758 9499
rect 10772 9447 10818 9499
rect 10818 9447 10824 9499
rect 10706 9380 10712 9432
rect 10712 9380 10758 9432
rect 10772 9380 10818 9432
rect 10818 9380 10824 9432
rect 10706 7840 10712 7892
rect 10712 7840 10758 7892
rect 10772 7840 10818 7892
rect 10818 7840 10824 7892
rect 10706 7774 10712 7826
rect 10712 7774 10758 7826
rect 10772 7774 10818 7826
rect 10818 7774 10824 7826
rect 10706 7708 10712 7760
rect 10712 7708 10758 7760
rect 10772 7708 10818 7760
rect 10818 7708 10824 7760
rect 10706 7642 10712 7694
rect 10712 7642 10758 7694
rect 10772 7642 10818 7694
rect 10818 7642 10824 7694
rect 10706 7576 10712 7628
rect 10712 7576 10758 7628
rect 10772 7576 10818 7628
rect 10818 7576 10824 7628
rect 10706 7510 10712 7562
rect 10712 7510 10758 7562
rect 10772 7510 10818 7562
rect 10818 7510 10824 7562
rect 10706 7443 10712 7495
rect 10712 7443 10758 7495
rect 10772 7443 10818 7495
rect 10818 7443 10824 7495
rect 10706 7380 10712 7428
rect 10712 7380 10758 7428
rect 10772 7380 10818 7428
rect 10818 7380 10824 7428
rect 10706 7376 10758 7380
rect 10772 7376 10824 7380
rect 10706 5844 10712 5896
rect 10712 5844 10758 5896
rect 10772 5844 10818 5896
rect 10818 5844 10824 5896
rect 10706 5778 10712 5830
rect 10712 5778 10758 5830
rect 10772 5778 10818 5830
rect 10818 5778 10824 5830
rect 10706 5712 10712 5764
rect 10712 5712 10758 5764
rect 10772 5712 10818 5764
rect 10818 5712 10824 5764
rect 10706 5646 10712 5698
rect 10712 5646 10758 5698
rect 10772 5646 10818 5698
rect 10818 5646 10824 5698
rect 10706 5580 10712 5632
rect 10712 5580 10758 5632
rect 10772 5580 10818 5632
rect 10818 5580 10824 5632
rect 10706 5514 10712 5566
rect 10712 5514 10758 5566
rect 10772 5514 10818 5566
rect 10818 5514 10824 5566
rect 10706 5447 10712 5499
rect 10712 5447 10758 5499
rect 10772 5447 10818 5499
rect 10818 5447 10824 5499
rect 10706 5380 10712 5432
rect 10712 5380 10758 5432
rect 10772 5380 10818 5432
rect 10818 5380 10824 5432
rect 10983 14345 11035 14390
rect 10983 14338 10989 14345
rect 10989 14338 11023 14345
rect 11023 14338 11035 14345
rect 11049 14345 11101 14390
rect 11537 14668 11589 14720
rect 11603 14668 11655 14720
rect 11537 14602 11589 14654
rect 11603 14602 11655 14654
rect 11537 14536 11589 14588
rect 11603 14536 11655 14588
rect 11537 14470 11589 14522
rect 11603 14470 11655 14522
rect 11537 14404 11589 14456
rect 11603 14404 11655 14456
rect 11049 14338 11061 14345
rect 11061 14338 11095 14345
rect 11095 14338 11101 14345
rect 10983 14311 10989 14323
rect 10989 14311 11023 14323
rect 11023 14311 11035 14323
rect 10983 14271 11035 14311
rect 11049 14311 11061 14323
rect 11061 14311 11095 14323
rect 11095 14311 11101 14323
rect 11049 14271 11101 14311
rect 10983 14233 10989 14256
rect 10989 14233 11023 14256
rect 11023 14233 11035 14256
rect 10983 14204 11035 14233
rect 11049 14233 11061 14256
rect 11061 14233 11095 14256
rect 11095 14233 11101 14256
rect 11049 14204 11101 14233
rect 10983 12714 11035 12720
rect 10983 12680 10989 12714
rect 10989 12680 11023 12714
rect 11023 12680 11035 12714
rect 10983 12668 11035 12680
rect 11049 12714 11101 12720
rect 11049 12680 11061 12714
rect 11061 12680 11095 12714
rect 11095 12680 11101 12714
rect 11049 12668 11101 12680
rect 10983 12641 11035 12654
rect 10983 12607 10989 12641
rect 10989 12607 11023 12641
rect 11023 12607 11035 12641
rect 10983 12602 11035 12607
rect 11049 12641 11101 12654
rect 11049 12607 11061 12641
rect 11061 12607 11095 12641
rect 11095 12607 11101 12641
rect 11049 12602 11101 12607
rect 10983 12568 11035 12588
rect 10983 12536 10989 12568
rect 10989 12536 11023 12568
rect 11023 12536 11035 12568
rect 11049 12568 11101 12588
rect 11049 12536 11061 12568
rect 11061 12536 11095 12568
rect 11095 12536 11101 12568
rect 10983 12495 11035 12522
rect 10983 12470 10989 12495
rect 10989 12470 11023 12495
rect 11023 12470 11035 12495
rect 11049 12495 11101 12522
rect 11049 12470 11061 12495
rect 11061 12470 11095 12495
rect 11095 12470 11101 12495
rect 10983 12422 11035 12456
rect 11049 12422 11101 12456
rect 10983 12404 10989 12422
rect 10989 12404 11035 12422
rect 11049 12404 11095 12422
rect 11095 12404 11101 12422
rect 10983 12338 10989 12390
rect 10989 12338 11035 12390
rect 11049 12338 11095 12390
rect 11095 12338 11101 12390
rect 10983 12271 10989 12323
rect 10989 12271 11035 12323
rect 11049 12271 11095 12323
rect 11095 12271 11101 12323
rect 10983 12204 10989 12256
rect 10989 12204 11035 12256
rect 11049 12204 11095 12256
rect 11095 12204 11101 12256
rect 10983 10714 11035 10724
rect 10983 10680 10989 10714
rect 10989 10680 11023 10714
rect 11023 10680 11035 10714
rect 10983 10672 11035 10680
rect 11049 10714 11101 10724
rect 11049 10680 11061 10714
rect 11061 10680 11095 10714
rect 11095 10680 11101 10714
rect 11049 10672 11101 10680
rect 10983 10641 11035 10658
rect 10983 10607 10989 10641
rect 10989 10607 11023 10641
rect 11023 10607 11035 10641
rect 10983 10606 11035 10607
rect 11049 10641 11101 10658
rect 11049 10607 11061 10641
rect 11061 10607 11095 10641
rect 11095 10607 11101 10641
rect 11049 10606 11101 10607
rect 10983 10568 11035 10592
rect 10983 10540 10989 10568
rect 10989 10540 11023 10568
rect 11023 10540 11035 10568
rect 11049 10568 11101 10592
rect 11049 10540 11061 10568
rect 11061 10540 11095 10568
rect 11095 10540 11101 10568
rect 10983 10495 11035 10526
rect 10983 10474 10989 10495
rect 10989 10474 11023 10495
rect 11023 10474 11035 10495
rect 11049 10495 11101 10526
rect 11049 10474 11061 10495
rect 11061 10474 11095 10495
rect 11095 10474 11101 10495
rect 10983 10422 11035 10460
rect 11049 10422 11101 10460
rect 10983 10408 10989 10422
rect 10989 10408 11035 10422
rect 11049 10408 11095 10422
rect 11095 10408 11101 10422
rect 10983 10342 10989 10394
rect 10989 10342 11035 10394
rect 11049 10342 11095 10394
rect 11095 10342 11101 10394
rect 10983 10275 10989 10327
rect 10989 10275 11035 10327
rect 11049 10275 11095 10327
rect 11095 10275 11101 10327
rect 10983 10208 10989 10260
rect 10989 10208 11035 10260
rect 11049 10208 11095 10260
rect 11095 10208 11101 10260
rect 10983 8714 11035 8720
rect 10983 8680 10989 8714
rect 10989 8680 11023 8714
rect 11023 8680 11035 8714
rect 10983 8668 11035 8680
rect 11049 8714 11101 8720
rect 11049 8680 11061 8714
rect 11061 8680 11095 8714
rect 11095 8680 11101 8714
rect 11049 8668 11101 8680
rect 10983 8641 11035 8654
rect 10983 8607 10989 8641
rect 10989 8607 11023 8641
rect 11023 8607 11035 8641
rect 10983 8602 11035 8607
rect 11049 8641 11101 8654
rect 11049 8607 11061 8641
rect 11061 8607 11095 8641
rect 11095 8607 11101 8641
rect 11049 8602 11101 8607
rect 10983 8568 11035 8588
rect 10983 8536 10989 8568
rect 10989 8536 11023 8568
rect 11023 8536 11035 8568
rect 11049 8568 11101 8588
rect 11049 8536 11061 8568
rect 11061 8536 11095 8568
rect 11095 8536 11101 8568
rect 10983 8495 11035 8522
rect 10983 8470 10989 8495
rect 10989 8470 11023 8495
rect 11023 8470 11035 8495
rect 11049 8495 11101 8522
rect 11049 8470 11061 8495
rect 11061 8470 11095 8495
rect 11095 8470 11101 8495
rect 10983 8422 11035 8456
rect 11049 8422 11101 8456
rect 10983 8404 10989 8422
rect 10989 8404 11035 8422
rect 11049 8404 11095 8422
rect 11095 8404 11101 8422
rect 10983 8338 10989 8390
rect 10989 8338 11035 8390
rect 11049 8338 11095 8390
rect 11095 8338 11101 8390
rect 10983 8271 10989 8323
rect 10989 8271 11035 8323
rect 11049 8271 11095 8323
rect 11095 8271 11101 8323
rect 10983 8204 10989 8256
rect 10989 8204 11035 8256
rect 11049 8204 11095 8256
rect 11095 8204 11101 8256
rect 10983 6714 11035 6724
rect 10983 6680 10989 6714
rect 10989 6680 11023 6714
rect 11023 6680 11035 6714
rect 10983 6672 11035 6680
rect 11049 6714 11101 6724
rect 11049 6680 11061 6714
rect 11061 6680 11095 6714
rect 11095 6680 11101 6714
rect 11049 6672 11101 6680
rect 10983 6641 11035 6658
rect 10983 6607 10989 6641
rect 10989 6607 11023 6641
rect 11023 6607 11035 6641
rect 10983 6606 11035 6607
rect 11049 6641 11101 6658
rect 11049 6607 11061 6641
rect 11061 6607 11095 6641
rect 11095 6607 11101 6641
rect 11049 6606 11101 6607
rect 10983 6568 11035 6592
rect 10983 6540 10989 6568
rect 10989 6540 11023 6568
rect 11023 6540 11035 6568
rect 11049 6568 11101 6592
rect 11049 6540 11061 6568
rect 11061 6540 11095 6568
rect 11095 6540 11101 6568
rect 10983 6495 11035 6526
rect 10983 6474 10989 6495
rect 10989 6474 11023 6495
rect 11023 6474 11035 6495
rect 11049 6495 11101 6526
rect 11049 6474 11061 6495
rect 11061 6474 11095 6495
rect 11095 6474 11101 6495
rect 10983 6422 11035 6460
rect 11049 6422 11101 6460
rect 10983 6408 10989 6422
rect 10989 6408 11035 6422
rect 11049 6408 11095 6422
rect 11095 6408 11101 6422
rect 10983 6342 10989 6394
rect 10989 6342 11035 6394
rect 11049 6342 11095 6394
rect 11095 6342 11101 6394
rect 10983 6275 10989 6327
rect 10989 6275 11035 6327
rect 11049 6275 11095 6327
rect 11095 6275 11101 6327
rect 10983 6208 10989 6260
rect 10989 6208 11035 6260
rect 11049 6208 11095 6260
rect 11095 6208 11101 6260
rect 11260 13877 11312 13892
rect 11260 13843 11266 13877
rect 11266 13843 11300 13877
rect 11300 13843 11312 13877
rect 11260 13840 11312 13843
rect 11326 13877 11378 13892
rect 11326 13843 11338 13877
rect 11338 13843 11372 13877
rect 11372 13843 11378 13877
rect 11326 13840 11378 13843
rect 11260 13799 11312 13826
rect 11260 13774 11266 13799
rect 11266 13774 11300 13799
rect 11300 13774 11312 13799
rect 11326 13799 11378 13826
rect 11326 13774 11338 13799
rect 11338 13774 11372 13799
rect 11372 13774 11378 13799
rect 11260 13722 11312 13760
rect 11260 13708 11266 13722
rect 11266 13708 11300 13722
rect 11300 13708 11312 13722
rect 11326 13722 11378 13760
rect 11326 13708 11338 13722
rect 11338 13708 11372 13722
rect 11372 13708 11378 13722
rect 11260 13688 11266 13694
rect 11266 13688 11300 13694
rect 11300 13688 11312 13694
rect 11260 13645 11312 13688
rect 11260 13642 11266 13645
rect 11266 13642 11300 13645
rect 11300 13642 11312 13645
rect 11326 13688 11338 13694
rect 11338 13688 11372 13694
rect 11372 13688 11378 13694
rect 11326 13645 11378 13688
rect 11326 13642 11338 13645
rect 11338 13642 11372 13645
rect 11372 13642 11378 13645
rect 11260 13611 11266 13628
rect 11266 13611 11300 13628
rect 11300 13611 11312 13628
rect 11260 13576 11312 13611
rect 11326 13611 11338 13628
rect 11338 13611 11372 13628
rect 11372 13611 11378 13628
rect 11326 13576 11378 13611
rect 11260 13534 11266 13562
rect 11266 13534 11300 13562
rect 11300 13534 11312 13562
rect 11260 13510 11312 13534
rect 11326 13534 11338 13562
rect 11338 13534 11372 13562
rect 11372 13534 11378 13562
rect 11326 13510 11378 13534
rect 11260 13491 11312 13495
rect 11260 13457 11266 13491
rect 11266 13457 11300 13491
rect 11300 13457 11312 13491
rect 11260 13443 11312 13457
rect 11326 13491 11378 13495
rect 11326 13457 11338 13491
rect 11338 13457 11372 13491
rect 11372 13457 11378 13491
rect 11326 13443 11378 13457
rect 11260 13414 11312 13428
rect 11260 13380 11266 13414
rect 11266 13380 11300 13414
rect 11300 13380 11312 13414
rect 11260 13376 11312 13380
rect 11326 13414 11378 13428
rect 11326 13380 11338 13414
rect 11338 13380 11372 13414
rect 11372 13380 11378 13414
rect 11326 13376 11378 13380
rect 11260 11840 11266 11892
rect 11266 11840 11312 11892
rect 11326 11840 11372 11892
rect 11372 11840 11378 11892
rect 11260 11774 11266 11826
rect 11266 11774 11312 11826
rect 11326 11774 11372 11826
rect 11372 11774 11378 11826
rect 11260 11708 11266 11760
rect 11266 11708 11312 11760
rect 11326 11708 11372 11760
rect 11372 11708 11378 11760
rect 11260 11642 11266 11694
rect 11266 11642 11312 11694
rect 11326 11642 11372 11694
rect 11372 11642 11378 11694
rect 11260 11576 11266 11628
rect 11266 11576 11312 11628
rect 11326 11576 11372 11628
rect 11372 11576 11378 11628
rect 11260 11510 11266 11562
rect 11266 11510 11312 11562
rect 11326 11510 11372 11562
rect 11372 11510 11378 11562
rect 11260 11443 11266 11495
rect 11266 11443 11312 11495
rect 11326 11443 11372 11495
rect 11372 11443 11378 11495
rect 11260 11380 11266 11428
rect 11266 11380 11312 11428
rect 11326 11380 11372 11428
rect 11372 11380 11378 11428
rect 11260 11376 11312 11380
rect 11326 11376 11378 11380
rect 11260 9844 11266 9896
rect 11266 9844 11312 9896
rect 11326 9844 11372 9896
rect 11372 9844 11378 9896
rect 11260 9778 11266 9830
rect 11266 9778 11312 9830
rect 11326 9778 11372 9830
rect 11372 9778 11378 9830
rect 11260 9712 11266 9764
rect 11266 9712 11312 9764
rect 11326 9712 11372 9764
rect 11372 9712 11378 9764
rect 11260 9646 11266 9698
rect 11266 9646 11312 9698
rect 11326 9646 11372 9698
rect 11372 9646 11378 9698
rect 11260 9580 11266 9632
rect 11266 9580 11312 9632
rect 11326 9580 11372 9632
rect 11372 9580 11378 9632
rect 11260 9514 11266 9566
rect 11266 9514 11312 9566
rect 11326 9514 11372 9566
rect 11372 9514 11378 9566
rect 11260 9447 11266 9499
rect 11266 9447 11312 9499
rect 11326 9447 11372 9499
rect 11372 9447 11378 9499
rect 11260 9380 11266 9432
rect 11266 9380 11312 9432
rect 11326 9380 11372 9432
rect 11372 9380 11378 9432
rect 11260 7840 11266 7892
rect 11266 7840 11312 7892
rect 11326 7840 11372 7892
rect 11372 7840 11378 7892
rect 11260 7774 11266 7826
rect 11266 7774 11312 7826
rect 11326 7774 11372 7826
rect 11372 7774 11378 7826
rect 11260 7708 11266 7760
rect 11266 7708 11312 7760
rect 11326 7708 11372 7760
rect 11372 7708 11378 7760
rect 11260 7642 11266 7694
rect 11266 7642 11312 7694
rect 11326 7642 11372 7694
rect 11372 7642 11378 7694
rect 11260 7576 11266 7628
rect 11266 7576 11312 7628
rect 11326 7576 11372 7628
rect 11372 7576 11378 7628
rect 11260 7510 11266 7562
rect 11266 7510 11312 7562
rect 11326 7510 11372 7562
rect 11372 7510 11378 7562
rect 11260 7443 11266 7495
rect 11266 7443 11312 7495
rect 11326 7443 11372 7495
rect 11372 7443 11378 7495
rect 11260 7380 11266 7428
rect 11266 7380 11312 7428
rect 11326 7380 11372 7428
rect 11372 7380 11378 7428
rect 11260 7376 11312 7380
rect 11326 7376 11378 7380
rect 11260 5844 11266 5896
rect 11266 5844 11312 5896
rect 11326 5844 11372 5896
rect 11372 5844 11378 5896
rect 11260 5778 11266 5830
rect 11266 5778 11312 5830
rect 11326 5778 11372 5830
rect 11372 5778 11378 5830
rect 11260 5712 11266 5764
rect 11266 5712 11312 5764
rect 11326 5712 11372 5764
rect 11372 5712 11378 5764
rect 11260 5646 11266 5698
rect 11266 5646 11312 5698
rect 11326 5646 11372 5698
rect 11372 5646 11378 5698
rect 11260 5580 11266 5632
rect 11266 5580 11312 5632
rect 11326 5580 11372 5632
rect 11372 5580 11378 5632
rect 11260 5514 11266 5566
rect 11266 5514 11312 5566
rect 11326 5514 11372 5566
rect 11372 5514 11378 5566
rect 11260 5447 11266 5499
rect 11266 5447 11312 5499
rect 11326 5447 11372 5499
rect 11372 5447 11378 5499
rect 11260 5380 11266 5432
rect 11266 5380 11312 5432
rect 11326 5380 11372 5432
rect 11372 5380 11378 5432
rect 11537 14345 11589 14390
rect 11537 14338 11543 14345
rect 11543 14338 11577 14345
rect 11577 14338 11589 14345
rect 11603 14345 11655 14390
rect 12091 14668 12143 14720
rect 12157 14668 12209 14720
rect 12091 14602 12143 14654
rect 12157 14602 12209 14654
rect 12091 14536 12143 14588
rect 12157 14536 12209 14588
rect 12091 14470 12143 14522
rect 12157 14470 12209 14522
rect 12091 14404 12143 14456
rect 12157 14404 12209 14456
rect 11603 14338 11615 14345
rect 11615 14338 11649 14345
rect 11649 14338 11655 14345
rect 11537 14311 11543 14323
rect 11543 14311 11577 14323
rect 11577 14311 11589 14323
rect 11537 14271 11589 14311
rect 11603 14311 11615 14323
rect 11615 14311 11649 14323
rect 11649 14311 11655 14323
rect 11603 14271 11655 14311
rect 11537 14233 11543 14256
rect 11543 14233 11577 14256
rect 11577 14233 11589 14256
rect 11537 14204 11589 14233
rect 11603 14233 11615 14256
rect 11615 14233 11649 14256
rect 11649 14233 11655 14256
rect 11603 14204 11655 14233
rect 11537 12714 11589 12720
rect 11537 12680 11543 12714
rect 11543 12680 11577 12714
rect 11577 12680 11589 12714
rect 11537 12668 11589 12680
rect 11603 12714 11655 12720
rect 11603 12680 11615 12714
rect 11615 12680 11649 12714
rect 11649 12680 11655 12714
rect 11603 12668 11655 12680
rect 11537 12641 11589 12654
rect 11537 12607 11543 12641
rect 11543 12607 11577 12641
rect 11577 12607 11589 12641
rect 11537 12602 11589 12607
rect 11603 12641 11655 12654
rect 11603 12607 11615 12641
rect 11615 12607 11649 12641
rect 11649 12607 11655 12641
rect 11603 12602 11655 12607
rect 11537 12568 11589 12588
rect 11537 12536 11543 12568
rect 11543 12536 11577 12568
rect 11577 12536 11589 12568
rect 11603 12568 11655 12588
rect 11603 12536 11615 12568
rect 11615 12536 11649 12568
rect 11649 12536 11655 12568
rect 11537 12495 11589 12522
rect 11537 12470 11543 12495
rect 11543 12470 11577 12495
rect 11577 12470 11589 12495
rect 11603 12495 11655 12522
rect 11603 12470 11615 12495
rect 11615 12470 11649 12495
rect 11649 12470 11655 12495
rect 11537 12422 11589 12456
rect 11603 12422 11655 12456
rect 11537 12404 11543 12422
rect 11543 12404 11589 12422
rect 11603 12404 11649 12422
rect 11649 12404 11655 12422
rect 11537 12338 11543 12390
rect 11543 12338 11589 12390
rect 11603 12338 11649 12390
rect 11649 12338 11655 12390
rect 11537 12271 11543 12323
rect 11543 12271 11589 12323
rect 11603 12271 11649 12323
rect 11649 12271 11655 12323
rect 11537 12204 11543 12256
rect 11543 12204 11589 12256
rect 11603 12204 11649 12256
rect 11649 12204 11655 12256
rect 11537 10714 11589 10724
rect 11537 10680 11543 10714
rect 11543 10680 11577 10714
rect 11577 10680 11589 10714
rect 11537 10672 11589 10680
rect 11603 10714 11655 10724
rect 11603 10680 11615 10714
rect 11615 10680 11649 10714
rect 11649 10680 11655 10714
rect 11603 10672 11655 10680
rect 11537 10641 11589 10658
rect 11537 10607 11543 10641
rect 11543 10607 11577 10641
rect 11577 10607 11589 10641
rect 11537 10606 11589 10607
rect 11603 10641 11655 10658
rect 11603 10607 11615 10641
rect 11615 10607 11649 10641
rect 11649 10607 11655 10641
rect 11603 10606 11655 10607
rect 11537 10568 11589 10592
rect 11537 10540 11543 10568
rect 11543 10540 11577 10568
rect 11577 10540 11589 10568
rect 11603 10568 11655 10592
rect 11603 10540 11615 10568
rect 11615 10540 11649 10568
rect 11649 10540 11655 10568
rect 11537 10495 11589 10526
rect 11537 10474 11543 10495
rect 11543 10474 11577 10495
rect 11577 10474 11589 10495
rect 11603 10495 11655 10526
rect 11603 10474 11615 10495
rect 11615 10474 11649 10495
rect 11649 10474 11655 10495
rect 11537 10422 11589 10460
rect 11603 10422 11655 10460
rect 11537 10408 11543 10422
rect 11543 10408 11589 10422
rect 11603 10408 11649 10422
rect 11649 10408 11655 10422
rect 11537 10342 11543 10394
rect 11543 10342 11589 10394
rect 11603 10342 11649 10394
rect 11649 10342 11655 10394
rect 11537 10275 11543 10327
rect 11543 10275 11589 10327
rect 11603 10275 11649 10327
rect 11649 10275 11655 10327
rect 11537 10208 11543 10260
rect 11543 10208 11589 10260
rect 11603 10208 11649 10260
rect 11649 10208 11655 10260
rect 11537 8714 11589 8720
rect 11537 8680 11543 8714
rect 11543 8680 11577 8714
rect 11577 8680 11589 8714
rect 11537 8668 11589 8680
rect 11603 8714 11655 8720
rect 11603 8680 11615 8714
rect 11615 8680 11649 8714
rect 11649 8680 11655 8714
rect 11603 8668 11655 8680
rect 11537 8641 11589 8654
rect 11537 8607 11543 8641
rect 11543 8607 11577 8641
rect 11577 8607 11589 8641
rect 11537 8602 11589 8607
rect 11603 8641 11655 8654
rect 11603 8607 11615 8641
rect 11615 8607 11649 8641
rect 11649 8607 11655 8641
rect 11603 8602 11655 8607
rect 11537 8568 11589 8588
rect 11537 8536 11543 8568
rect 11543 8536 11577 8568
rect 11577 8536 11589 8568
rect 11603 8568 11655 8588
rect 11603 8536 11615 8568
rect 11615 8536 11649 8568
rect 11649 8536 11655 8568
rect 11537 8495 11589 8522
rect 11537 8470 11543 8495
rect 11543 8470 11577 8495
rect 11577 8470 11589 8495
rect 11603 8495 11655 8522
rect 11603 8470 11615 8495
rect 11615 8470 11649 8495
rect 11649 8470 11655 8495
rect 11537 8422 11589 8456
rect 11603 8422 11655 8456
rect 11537 8404 11543 8422
rect 11543 8404 11589 8422
rect 11603 8404 11649 8422
rect 11649 8404 11655 8422
rect 11537 8338 11543 8390
rect 11543 8338 11589 8390
rect 11603 8338 11649 8390
rect 11649 8338 11655 8390
rect 11537 8271 11543 8323
rect 11543 8271 11589 8323
rect 11603 8271 11649 8323
rect 11649 8271 11655 8323
rect 11537 8204 11543 8256
rect 11543 8204 11589 8256
rect 11603 8204 11649 8256
rect 11649 8204 11655 8256
rect 11537 6714 11589 6724
rect 11537 6680 11543 6714
rect 11543 6680 11577 6714
rect 11577 6680 11589 6714
rect 11537 6672 11589 6680
rect 11603 6714 11655 6724
rect 11603 6680 11615 6714
rect 11615 6680 11649 6714
rect 11649 6680 11655 6714
rect 11603 6672 11655 6680
rect 11537 6641 11589 6658
rect 11537 6607 11543 6641
rect 11543 6607 11577 6641
rect 11577 6607 11589 6641
rect 11537 6606 11589 6607
rect 11603 6641 11655 6658
rect 11603 6607 11615 6641
rect 11615 6607 11649 6641
rect 11649 6607 11655 6641
rect 11603 6606 11655 6607
rect 11537 6568 11589 6592
rect 11537 6540 11543 6568
rect 11543 6540 11577 6568
rect 11577 6540 11589 6568
rect 11603 6568 11655 6592
rect 11603 6540 11615 6568
rect 11615 6540 11649 6568
rect 11649 6540 11655 6568
rect 11537 6495 11589 6526
rect 11537 6474 11543 6495
rect 11543 6474 11577 6495
rect 11577 6474 11589 6495
rect 11603 6495 11655 6526
rect 11603 6474 11615 6495
rect 11615 6474 11649 6495
rect 11649 6474 11655 6495
rect 11537 6422 11589 6460
rect 11603 6422 11655 6460
rect 11537 6408 11543 6422
rect 11543 6408 11589 6422
rect 11603 6408 11649 6422
rect 11649 6408 11655 6422
rect 11537 6342 11543 6394
rect 11543 6342 11589 6394
rect 11603 6342 11649 6394
rect 11649 6342 11655 6394
rect 11537 6275 11543 6327
rect 11543 6275 11589 6327
rect 11603 6275 11649 6327
rect 11649 6275 11655 6327
rect 11537 6208 11543 6260
rect 11543 6208 11589 6260
rect 11603 6208 11649 6260
rect 11649 6208 11655 6260
rect 11814 13877 11866 13892
rect 11814 13843 11820 13877
rect 11820 13843 11854 13877
rect 11854 13843 11866 13877
rect 11814 13840 11866 13843
rect 11880 13877 11932 13892
rect 11880 13843 11892 13877
rect 11892 13843 11926 13877
rect 11926 13843 11932 13877
rect 11880 13840 11932 13843
rect 11814 13799 11866 13826
rect 11814 13774 11820 13799
rect 11820 13774 11854 13799
rect 11854 13774 11866 13799
rect 11880 13799 11932 13826
rect 11880 13774 11892 13799
rect 11892 13774 11926 13799
rect 11926 13774 11932 13799
rect 11814 13722 11866 13760
rect 11814 13708 11820 13722
rect 11820 13708 11854 13722
rect 11854 13708 11866 13722
rect 11880 13722 11932 13760
rect 11880 13708 11892 13722
rect 11892 13708 11926 13722
rect 11926 13708 11932 13722
rect 11814 13688 11820 13694
rect 11820 13688 11854 13694
rect 11854 13688 11866 13694
rect 11814 13645 11866 13688
rect 11814 13642 11820 13645
rect 11820 13642 11854 13645
rect 11854 13642 11866 13645
rect 11880 13688 11892 13694
rect 11892 13688 11926 13694
rect 11926 13688 11932 13694
rect 11880 13645 11932 13688
rect 11880 13642 11892 13645
rect 11892 13642 11926 13645
rect 11926 13642 11932 13645
rect 11814 13611 11820 13628
rect 11820 13611 11854 13628
rect 11854 13611 11866 13628
rect 11814 13576 11866 13611
rect 11880 13611 11892 13628
rect 11892 13611 11926 13628
rect 11926 13611 11932 13628
rect 11880 13576 11932 13611
rect 11814 13534 11820 13562
rect 11820 13534 11854 13562
rect 11854 13534 11866 13562
rect 11814 13510 11866 13534
rect 11880 13534 11892 13562
rect 11892 13534 11926 13562
rect 11926 13534 11932 13562
rect 11880 13510 11932 13534
rect 11814 13491 11866 13495
rect 11814 13457 11820 13491
rect 11820 13457 11854 13491
rect 11854 13457 11866 13491
rect 11814 13443 11866 13457
rect 11880 13491 11932 13495
rect 11880 13457 11892 13491
rect 11892 13457 11926 13491
rect 11926 13457 11932 13491
rect 11880 13443 11932 13457
rect 11814 13414 11866 13428
rect 11814 13380 11820 13414
rect 11820 13380 11854 13414
rect 11854 13380 11866 13414
rect 11814 13376 11866 13380
rect 11880 13414 11932 13428
rect 11880 13380 11892 13414
rect 11892 13380 11926 13414
rect 11926 13380 11932 13414
rect 11880 13376 11932 13380
rect 11814 11840 11820 11892
rect 11820 11840 11866 11892
rect 11880 11840 11926 11892
rect 11926 11840 11932 11892
rect 11814 11774 11820 11826
rect 11820 11774 11866 11826
rect 11880 11774 11926 11826
rect 11926 11774 11932 11826
rect 11814 11708 11820 11760
rect 11820 11708 11866 11760
rect 11880 11708 11926 11760
rect 11926 11708 11932 11760
rect 11814 11642 11820 11694
rect 11820 11642 11866 11694
rect 11880 11642 11926 11694
rect 11926 11642 11932 11694
rect 11814 11576 11820 11628
rect 11820 11576 11866 11628
rect 11880 11576 11926 11628
rect 11926 11576 11932 11628
rect 11814 11510 11820 11562
rect 11820 11510 11866 11562
rect 11880 11510 11926 11562
rect 11926 11510 11932 11562
rect 11814 11443 11820 11495
rect 11820 11443 11866 11495
rect 11880 11443 11926 11495
rect 11926 11443 11932 11495
rect 11814 11380 11820 11428
rect 11820 11380 11866 11428
rect 11880 11380 11926 11428
rect 11926 11380 11932 11428
rect 11814 11376 11866 11380
rect 11880 11376 11932 11380
rect 11814 9844 11820 9896
rect 11820 9844 11866 9896
rect 11880 9844 11926 9896
rect 11926 9844 11932 9896
rect 11814 9778 11820 9830
rect 11820 9778 11866 9830
rect 11880 9778 11926 9830
rect 11926 9778 11932 9830
rect 11814 9712 11820 9764
rect 11820 9712 11866 9764
rect 11880 9712 11926 9764
rect 11926 9712 11932 9764
rect 11814 9646 11820 9698
rect 11820 9646 11866 9698
rect 11880 9646 11926 9698
rect 11926 9646 11932 9698
rect 11814 9580 11820 9632
rect 11820 9580 11866 9632
rect 11880 9580 11926 9632
rect 11926 9580 11932 9632
rect 11814 9514 11820 9566
rect 11820 9514 11866 9566
rect 11880 9514 11926 9566
rect 11926 9514 11932 9566
rect 11814 9447 11820 9499
rect 11820 9447 11866 9499
rect 11880 9447 11926 9499
rect 11926 9447 11932 9499
rect 11814 9380 11820 9432
rect 11820 9380 11866 9432
rect 11880 9380 11926 9432
rect 11926 9380 11932 9432
rect 11814 7840 11820 7892
rect 11820 7840 11866 7892
rect 11880 7840 11926 7892
rect 11926 7840 11932 7892
rect 11814 7774 11820 7826
rect 11820 7774 11866 7826
rect 11880 7774 11926 7826
rect 11926 7774 11932 7826
rect 11814 7708 11820 7760
rect 11820 7708 11866 7760
rect 11880 7708 11926 7760
rect 11926 7708 11932 7760
rect 11814 7642 11820 7694
rect 11820 7642 11866 7694
rect 11880 7642 11926 7694
rect 11926 7642 11932 7694
rect 11814 7576 11820 7628
rect 11820 7576 11866 7628
rect 11880 7576 11926 7628
rect 11926 7576 11932 7628
rect 11814 7510 11820 7562
rect 11820 7510 11866 7562
rect 11880 7510 11926 7562
rect 11926 7510 11932 7562
rect 11814 7443 11820 7495
rect 11820 7443 11866 7495
rect 11880 7443 11926 7495
rect 11926 7443 11932 7495
rect 11814 7380 11820 7428
rect 11820 7380 11866 7428
rect 11880 7380 11926 7428
rect 11926 7380 11932 7428
rect 11814 7376 11866 7380
rect 11880 7376 11932 7380
rect 11814 5844 11820 5896
rect 11820 5844 11866 5896
rect 11880 5844 11926 5896
rect 11926 5844 11932 5896
rect 11814 5778 11820 5830
rect 11820 5778 11866 5830
rect 11880 5778 11926 5830
rect 11926 5778 11932 5830
rect 11814 5712 11820 5764
rect 11820 5712 11866 5764
rect 11880 5712 11926 5764
rect 11926 5712 11932 5764
rect 11814 5646 11820 5698
rect 11820 5646 11866 5698
rect 11880 5646 11926 5698
rect 11926 5646 11932 5698
rect 11814 5580 11820 5632
rect 11820 5580 11866 5632
rect 11880 5580 11926 5632
rect 11926 5580 11932 5632
rect 11814 5514 11820 5566
rect 11820 5514 11866 5566
rect 11880 5514 11926 5566
rect 11926 5514 11932 5566
rect 11814 5447 11820 5499
rect 11820 5447 11866 5499
rect 11880 5447 11926 5499
rect 11926 5447 11932 5499
rect 11814 5380 11820 5432
rect 11820 5380 11866 5432
rect 11880 5380 11926 5432
rect 11926 5380 11932 5432
rect 12091 14345 12143 14390
rect 12091 14338 12097 14345
rect 12097 14338 12131 14345
rect 12131 14338 12143 14345
rect 12157 14345 12209 14390
rect 12645 14668 12697 14720
rect 12711 14668 12763 14720
rect 12645 14602 12697 14654
rect 12711 14602 12763 14654
rect 12645 14536 12697 14588
rect 12711 14536 12763 14588
rect 12645 14470 12697 14522
rect 12711 14470 12763 14522
rect 12645 14404 12697 14456
rect 12711 14404 12763 14456
rect 12157 14338 12169 14345
rect 12169 14338 12203 14345
rect 12203 14338 12209 14345
rect 12091 14311 12097 14323
rect 12097 14311 12131 14323
rect 12131 14311 12143 14323
rect 12091 14271 12143 14311
rect 12157 14311 12169 14323
rect 12169 14311 12203 14323
rect 12203 14311 12209 14323
rect 12157 14271 12209 14311
rect 12091 14233 12097 14256
rect 12097 14233 12131 14256
rect 12131 14233 12143 14256
rect 12091 14204 12143 14233
rect 12157 14233 12169 14256
rect 12169 14233 12203 14256
rect 12203 14233 12209 14256
rect 12157 14204 12209 14233
rect 12091 12714 12143 12720
rect 12091 12680 12097 12714
rect 12097 12680 12131 12714
rect 12131 12680 12143 12714
rect 12091 12668 12143 12680
rect 12157 12714 12209 12720
rect 12157 12680 12169 12714
rect 12169 12680 12203 12714
rect 12203 12680 12209 12714
rect 12157 12668 12209 12680
rect 12091 12641 12143 12654
rect 12091 12607 12097 12641
rect 12097 12607 12131 12641
rect 12131 12607 12143 12641
rect 12091 12602 12143 12607
rect 12157 12641 12209 12654
rect 12157 12607 12169 12641
rect 12169 12607 12203 12641
rect 12203 12607 12209 12641
rect 12157 12602 12209 12607
rect 12091 12568 12143 12588
rect 12091 12536 12097 12568
rect 12097 12536 12131 12568
rect 12131 12536 12143 12568
rect 12157 12568 12209 12588
rect 12157 12536 12169 12568
rect 12169 12536 12203 12568
rect 12203 12536 12209 12568
rect 12091 12495 12143 12522
rect 12091 12470 12097 12495
rect 12097 12470 12131 12495
rect 12131 12470 12143 12495
rect 12157 12495 12209 12522
rect 12157 12470 12169 12495
rect 12169 12470 12203 12495
rect 12203 12470 12209 12495
rect 12091 12422 12143 12456
rect 12157 12422 12209 12456
rect 12091 12404 12097 12422
rect 12097 12404 12143 12422
rect 12157 12404 12203 12422
rect 12203 12404 12209 12422
rect 12091 12338 12097 12390
rect 12097 12338 12143 12390
rect 12157 12338 12203 12390
rect 12203 12338 12209 12390
rect 12091 12271 12097 12323
rect 12097 12271 12143 12323
rect 12157 12271 12203 12323
rect 12203 12271 12209 12323
rect 12091 12204 12097 12256
rect 12097 12204 12143 12256
rect 12157 12204 12203 12256
rect 12203 12204 12209 12256
rect 12091 10714 12143 10724
rect 12091 10680 12097 10714
rect 12097 10680 12131 10714
rect 12131 10680 12143 10714
rect 12091 10672 12143 10680
rect 12157 10714 12209 10724
rect 12157 10680 12169 10714
rect 12169 10680 12203 10714
rect 12203 10680 12209 10714
rect 12157 10672 12209 10680
rect 12091 10641 12143 10658
rect 12091 10607 12097 10641
rect 12097 10607 12131 10641
rect 12131 10607 12143 10641
rect 12091 10606 12143 10607
rect 12157 10641 12209 10658
rect 12157 10607 12169 10641
rect 12169 10607 12203 10641
rect 12203 10607 12209 10641
rect 12157 10606 12209 10607
rect 12091 10568 12143 10592
rect 12091 10540 12097 10568
rect 12097 10540 12131 10568
rect 12131 10540 12143 10568
rect 12157 10568 12209 10592
rect 12157 10540 12169 10568
rect 12169 10540 12203 10568
rect 12203 10540 12209 10568
rect 12091 10495 12143 10526
rect 12091 10474 12097 10495
rect 12097 10474 12131 10495
rect 12131 10474 12143 10495
rect 12157 10495 12209 10526
rect 12157 10474 12169 10495
rect 12169 10474 12203 10495
rect 12203 10474 12209 10495
rect 12091 10422 12143 10460
rect 12157 10422 12209 10460
rect 12091 10408 12097 10422
rect 12097 10408 12143 10422
rect 12157 10408 12203 10422
rect 12203 10408 12209 10422
rect 12091 10342 12097 10394
rect 12097 10342 12143 10394
rect 12157 10342 12203 10394
rect 12203 10342 12209 10394
rect 12091 10275 12097 10327
rect 12097 10275 12143 10327
rect 12157 10275 12203 10327
rect 12203 10275 12209 10327
rect 12091 10208 12097 10260
rect 12097 10208 12143 10260
rect 12157 10208 12203 10260
rect 12203 10208 12209 10260
rect 12091 8714 12143 8720
rect 12091 8680 12097 8714
rect 12097 8680 12131 8714
rect 12131 8680 12143 8714
rect 12091 8668 12143 8680
rect 12157 8714 12209 8720
rect 12157 8680 12169 8714
rect 12169 8680 12203 8714
rect 12203 8680 12209 8714
rect 12157 8668 12209 8680
rect 12091 8641 12143 8654
rect 12091 8607 12097 8641
rect 12097 8607 12131 8641
rect 12131 8607 12143 8641
rect 12091 8602 12143 8607
rect 12157 8641 12209 8654
rect 12157 8607 12169 8641
rect 12169 8607 12203 8641
rect 12203 8607 12209 8641
rect 12157 8602 12209 8607
rect 12091 8568 12143 8588
rect 12091 8536 12097 8568
rect 12097 8536 12131 8568
rect 12131 8536 12143 8568
rect 12157 8568 12209 8588
rect 12157 8536 12169 8568
rect 12169 8536 12203 8568
rect 12203 8536 12209 8568
rect 12091 8495 12143 8522
rect 12091 8470 12097 8495
rect 12097 8470 12131 8495
rect 12131 8470 12143 8495
rect 12157 8495 12209 8522
rect 12157 8470 12169 8495
rect 12169 8470 12203 8495
rect 12203 8470 12209 8495
rect 12091 8422 12143 8456
rect 12157 8422 12209 8456
rect 12091 8404 12097 8422
rect 12097 8404 12143 8422
rect 12157 8404 12203 8422
rect 12203 8404 12209 8422
rect 12091 8338 12097 8390
rect 12097 8338 12143 8390
rect 12157 8338 12203 8390
rect 12203 8338 12209 8390
rect 12091 8271 12097 8323
rect 12097 8271 12143 8323
rect 12157 8271 12203 8323
rect 12203 8271 12209 8323
rect 12091 8204 12097 8256
rect 12097 8204 12143 8256
rect 12157 8204 12203 8256
rect 12203 8204 12209 8256
rect 12091 6714 12143 6724
rect 12091 6680 12097 6714
rect 12097 6680 12131 6714
rect 12131 6680 12143 6714
rect 12091 6672 12143 6680
rect 12157 6714 12209 6724
rect 12157 6680 12169 6714
rect 12169 6680 12203 6714
rect 12203 6680 12209 6714
rect 12157 6672 12209 6680
rect 12091 6641 12143 6658
rect 12091 6607 12097 6641
rect 12097 6607 12131 6641
rect 12131 6607 12143 6641
rect 12091 6606 12143 6607
rect 12157 6641 12209 6658
rect 12157 6607 12169 6641
rect 12169 6607 12203 6641
rect 12203 6607 12209 6641
rect 12157 6606 12209 6607
rect 12091 6568 12143 6592
rect 12091 6540 12097 6568
rect 12097 6540 12131 6568
rect 12131 6540 12143 6568
rect 12157 6568 12209 6592
rect 12157 6540 12169 6568
rect 12169 6540 12203 6568
rect 12203 6540 12209 6568
rect 12091 6495 12143 6526
rect 12091 6474 12097 6495
rect 12097 6474 12131 6495
rect 12131 6474 12143 6495
rect 12157 6495 12209 6526
rect 12157 6474 12169 6495
rect 12169 6474 12203 6495
rect 12203 6474 12209 6495
rect 12091 6422 12143 6460
rect 12157 6422 12209 6460
rect 12091 6408 12097 6422
rect 12097 6408 12143 6422
rect 12157 6408 12203 6422
rect 12203 6408 12209 6422
rect 12091 6342 12097 6394
rect 12097 6342 12143 6394
rect 12157 6342 12203 6394
rect 12203 6342 12209 6394
rect 12091 6275 12097 6327
rect 12097 6275 12143 6327
rect 12157 6275 12203 6327
rect 12203 6275 12209 6327
rect 12091 6208 12097 6260
rect 12097 6208 12143 6260
rect 12157 6208 12203 6260
rect 12203 6208 12209 6260
rect 12368 13877 12420 13892
rect 12368 13843 12374 13877
rect 12374 13843 12408 13877
rect 12408 13843 12420 13877
rect 12368 13840 12420 13843
rect 12434 13877 12486 13892
rect 12434 13843 12446 13877
rect 12446 13843 12480 13877
rect 12480 13843 12486 13877
rect 12434 13840 12486 13843
rect 12368 13799 12420 13826
rect 12368 13774 12374 13799
rect 12374 13774 12408 13799
rect 12408 13774 12420 13799
rect 12434 13799 12486 13826
rect 12434 13774 12446 13799
rect 12446 13774 12480 13799
rect 12480 13774 12486 13799
rect 12368 13722 12420 13760
rect 12368 13708 12374 13722
rect 12374 13708 12408 13722
rect 12408 13708 12420 13722
rect 12434 13722 12486 13760
rect 12434 13708 12446 13722
rect 12446 13708 12480 13722
rect 12480 13708 12486 13722
rect 12368 13688 12374 13694
rect 12374 13688 12408 13694
rect 12408 13688 12420 13694
rect 12368 13645 12420 13688
rect 12368 13642 12374 13645
rect 12374 13642 12408 13645
rect 12408 13642 12420 13645
rect 12434 13688 12446 13694
rect 12446 13688 12480 13694
rect 12480 13688 12486 13694
rect 12434 13645 12486 13688
rect 12434 13642 12446 13645
rect 12446 13642 12480 13645
rect 12480 13642 12486 13645
rect 12368 13611 12374 13628
rect 12374 13611 12408 13628
rect 12408 13611 12420 13628
rect 12368 13576 12420 13611
rect 12434 13611 12446 13628
rect 12446 13611 12480 13628
rect 12480 13611 12486 13628
rect 12434 13576 12486 13611
rect 12368 13534 12374 13562
rect 12374 13534 12408 13562
rect 12408 13534 12420 13562
rect 12368 13510 12420 13534
rect 12434 13534 12446 13562
rect 12446 13534 12480 13562
rect 12480 13534 12486 13562
rect 12434 13510 12486 13534
rect 12368 13491 12420 13495
rect 12368 13457 12374 13491
rect 12374 13457 12408 13491
rect 12408 13457 12420 13491
rect 12368 13443 12420 13457
rect 12434 13491 12486 13495
rect 12434 13457 12446 13491
rect 12446 13457 12480 13491
rect 12480 13457 12486 13491
rect 12434 13443 12486 13457
rect 12368 13414 12420 13428
rect 12368 13380 12374 13414
rect 12374 13380 12408 13414
rect 12408 13380 12420 13414
rect 12368 13376 12420 13380
rect 12434 13414 12486 13428
rect 12434 13380 12446 13414
rect 12446 13380 12480 13414
rect 12480 13380 12486 13414
rect 12434 13376 12486 13380
rect 12368 11840 12374 11892
rect 12374 11840 12420 11892
rect 12434 11840 12480 11892
rect 12480 11840 12486 11892
rect 12368 11774 12374 11826
rect 12374 11774 12420 11826
rect 12434 11774 12480 11826
rect 12480 11774 12486 11826
rect 12368 11708 12374 11760
rect 12374 11708 12420 11760
rect 12434 11708 12480 11760
rect 12480 11708 12486 11760
rect 12368 11642 12374 11694
rect 12374 11642 12420 11694
rect 12434 11642 12480 11694
rect 12480 11642 12486 11694
rect 12368 11576 12374 11628
rect 12374 11576 12420 11628
rect 12434 11576 12480 11628
rect 12480 11576 12486 11628
rect 12368 11510 12374 11562
rect 12374 11510 12420 11562
rect 12434 11510 12480 11562
rect 12480 11510 12486 11562
rect 12368 11443 12374 11495
rect 12374 11443 12420 11495
rect 12434 11443 12480 11495
rect 12480 11443 12486 11495
rect 12368 11380 12374 11428
rect 12374 11380 12420 11428
rect 12434 11380 12480 11428
rect 12480 11380 12486 11428
rect 12368 11376 12420 11380
rect 12434 11376 12486 11380
rect 12368 9844 12374 9896
rect 12374 9844 12420 9896
rect 12434 9844 12480 9896
rect 12480 9844 12486 9896
rect 12368 9778 12374 9830
rect 12374 9778 12420 9830
rect 12434 9778 12480 9830
rect 12480 9778 12486 9830
rect 12368 9712 12374 9764
rect 12374 9712 12420 9764
rect 12434 9712 12480 9764
rect 12480 9712 12486 9764
rect 12368 9646 12374 9698
rect 12374 9646 12420 9698
rect 12434 9646 12480 9698
rect 12480 9646 12486 9698
rect 12368 9580 12374 9632
rect 12374 9580 12420 9632
rect 12434 9580 12480 9632
rect 12480 9580 12486 9632
rect 12368 9514 12374 9566
rect 12374 9514 12420 9566
rect 12434 9514 12480 9566
rect 12480 9514 12486 9566
rect 12368 9447 12374 9499
rect 12374 9447 12420 9499
rect 12434 9447 12480 9499
rect 12480 9447 12486 9499
rect 12368 9380 12374 9432
rect 12374 9380 12420 9432
rect 12434 9380 12480 9432
rect 12480 9380 12486 9432
rect 12368 7839 12374 7891
rect 12374 7839 12420 7891
rect 12434 7839 12480 7891
rect 12480 7839 12486 7891
rect 12368 7773 12374 7825
rect 12374 7773 12420 7825
rect 12434 7773 12480 7825
rect 12480 7773 12486 7825
rect 12368 7707 12374 7759
rect 12374 7707 12420 7759
rect 12434 7707 12480 7759
rect 12480 7707 12486 7759
rect 12368 7641 12374 7693
rect 12374 7641 12420 7693
rect 12434 7641 12480 7693
rect 12480 7641 12486 7693
rect 12368 7575 12374 7627
rect 12374 7575 12420 7627
rect 12434 7575 12480 7627
rect 12480 7575 12486 7627
rect 12368 7509 12374 7561
rect 12374 7509 12420 7561
rect 12434 7509 12480 7561
rect 12480 7509 12486 7561
rect 12368 7442 12374 7494
rect 12374 7442 12420 7494
rect 12434 7442 12480 7494
rect 12480 7442 12486 7494
rect 12368 7380 12374 7427
rect 12374 7380 12420 7427
rect 12434 7380 12480 7427
rect 12480 7380 12486 7427
rect 12368 7375 12420 7380
rect 12434 7375 12486 7380
rect 12368 5842 12374 5894
rect 12374 5842 12420 5894
rect 12434 5842 12480 5894
rect 12480 5842 12486 5894
rect 12368 5776 12374 5828
rect 12374 5776 12420 5828
rect 12434 5776 12480 5828
rect 12480 5776 12486 5828
rect 12368 5710 12374 5762
rect 12374 5710 12420 5762
rect 12434 5710 12480 5762
rect 12480 5710 12486 5762
rect 12368 5644 12374 5696
rect 12374 5644 12420 5696
rect 12434 5644 12480 5696
rect 12480 5644 12486 5696
rect 12368 5578 12374 5630
rect 12374 5578 12420 5630
rect 12434 5578 12480 5630
rect 12480 5578 12486 5630
rect 12368 5512 12374 5564
rect 12374 5512 12420 5564
rect 12434 5512 12480 5564
rect 12480 5512 12486 5564
rect 12368 5445 12374 5497
rect 12374 5445 12420 5497
rect 12434 5445 12480 5497
rect 12480 5445 12486 5497
rect 12368 5380 12374 5430
rect 12374 5380 12420 5430
rect 12434 5380 12480 5430
rect 12480 5380 12486 5430
rect 12368 5378 12420 5380
rect 12434 5378 12486 5380
rect 12645 14345 12697 14390
rect 12645 14338 12651 14345
rect 12651 14338 12685 14345
rect 12685 14338 12697 14345
rect 12711 14345 12763 14390
rect 13200 14662 13252 14714
rect 13270 14662 13322 14714
rect 13340 14662 13392 14714
rect 13410 14662 13462 14714
rect 13480 14662 13490 14714
rect 13490 14662 13532 14714
rect 13550 14662 13596 14714
rect 13596 14662 13602 14714
rect 13200 14598 13252 14650
rect 13270 14598 13322 14650
rect 13340 14598 13392 14650
rect 13410 14598 13462 14650
rect 13480 14598 13490 14650
rect 13490 14598 13532 14650
rect 13550 14598 13596 14650
rect 13596 14598 13602 14650
rect 13200 14534 13252 14586
rect 13270 14534 13322 14586
rect 13340 14534 13392 14586
rect 13410 14534 13462 14586
rect 13480 14534 13490 14586
rect 13490 14534 13532 14586
rect 13550 14534 13596 14586
rect 13596 14534 13602 14586
rect 13200 14470 13252 14522
rect 13270 14470 13322 14522
rect 13340 14470 13392 14522
rect 13410 14470 13462 14522
rect 13480 14470 13490 14522
rect 13490 14470 13532 14522
rect 13550 14470 13596 14522
rect 13596 14470 13602 14522
rect 13200 14406 13252 14458
rect 13270 14406 13322 14458
rect 13340 14406 13392 14458
rect 13410 14406 13462 14458
rect 13480 14406 13490 14458
rect 13490 14406 13532 14458
rect 13550 14406 13596 14458
rect 13596 14406 13602 14458
rect 12711 14338 12723 14345
rect 12723 14338 12757 14345
rect 12757 14338 12763 14345
rect 12645 14311 12651 14323
rect 12651 14311 12685 14323
rect 12685 14311 12697 14323
rect 12645 14271 12697 14311
rect 12711 14311 12723 14323
rect 12723 14311 12757 14323
rect 12757 14311 12763 14323
rect 12711 14271 12763 14311
rect 12645 14233 12651 14256
rect 12651 14233 12685 14256
rect 12685 14233 12697 14256
rect 12645 14204 12697 14233
rect 12711 14233 12723 14256
rect 12723 14233 12757 14256
rect 12757 14233 12763 14256
rect 12711 14204 12763 14233
rect 12645 12714 12697 12720
rect 12645 12680 12651 12714
rect 12651 12680 12685 12714
rect 12685 12680 12697 12714
rect 12645 12668 12697 12680
rect 12711 12714 12763 12720
rect 12711 12680 12723 12714
rect 12723 12680 12757 12714
rect 12757 12680 12763 12714
rect 12711 12668 12763 12680
rect 12645 12641 12697 12654
rect 12645 12607 12651 12641
rect 12651 12607 12685 12641
rect 12685 12607 12697 12641
rect 12645 12602 12697 12607
rect 12711 12641 12763 12654
rect 12711 12607 12723 12641
rect 12723 12607 12757 12641
rect 12757 12607 12763 12641
rect 12711 12602 12763 12607
rect 12645 12568 12697 12588
rect 12645 12536 12651 12568
rect 12651 12536 12685 12568
rect 12685 12536 12697 12568
rect 12711 12568 12763 12588
rect 12711 12536 12723 12568
rect 12723 12536 12757 12568
rect 12757 12536 12763 12568
rect 12645 12495 12697 12522
rect 12645 12470 12651 12495
rect 12651 12470 12685 12495
rect 12685 12470 12697 12495
rect 12711 12495 12763 12522
rect 12711 12470 12723 12495
rect 12723 12470 12757 12495
rect 12757 12470 12763 12495
rect 12645 12422 12697 12456
rect 12711 12422 12763 12456
rect 12645 12404 12651 12422
rect 12651 12404 12697 12422
rect 12711 12404 12757 12422
rect 12757 12404 12763 12422
rect 12645 12338 12651 12390
rect 12651 12338 12697 12390
rect 12711 12338 12757 12390
rect 12757 12338 12763 12390
rect 12645 12271 12651 12323
rect 12651 12271 12697 12323
rect 12711 12271 12757 12323
rect 12757 12271 12763 12323
rect 12645 12204 12651 12256
rect 12651 12204 12697 12256
rect 12711 12204 12757 12256
rect 12757 12204 12763 12256
rect 12645 10714 12697 10724
rect 12645 10680 12651 10714
rect 12651 10680 12685 10714
rect 12685 10680 12697 10714
rect 12645 10672 12697 10680
rect 12711 10714 12763 10724
rect 12711 10680 12723 10714
rect 12723 10680 12757 10714
rect 12757 10680 12763 10714
rect 12711 10672 12763 10680
rect 12645 10641 12697 10658
rect 12645 10607 12651 10641
rect 12651 10607 12685 10641
rect 12685 10607 12697 10641
rect 12645 10606 12697 10607
rect 12711 10641 12763 10658
rect 12711 10607 12723 10641
rect 12723 10607 12757 10641
rect 12757 10607 12763 10641
rect 12711 10606 12763 10607
rect 12645 10568 12697 10592
rect 12645 10540 12651 10568
rect 12651 10540 12685 10568
rect 12685 10540 12697 10568
rect 12711 10568 12763 10592
rect 12711 10540 12723 10568
rect 12723 10540 12757 10568
rect 12757 10540 12763 10568
rect 12645 10495 12697 10526
rect 12645 10474 12651 10495
rect 12651 10474 12685 10495
rect 12685 10474 12697 10495
rect 12711 10495 12763 10526
rect 12711 10474 12723 10495
rect 12723 10474 12757 10495
rect 12757 10474 12763 10495
rect 12645 10422 12697 10460
rect 12711 10422 12763 10460
rect 12645 10408 12651 10422
rect 12651 10408 12697 10422
rect 12711 10408 12757 10422
rect 12757 10408 12763 10422
rect 12645 10342 12651 10394
rect 12651 10342 12697 10394
rect 12711 10342 12757 10394
rect 12757 10342 12763 10394
rect 12645 10275 12651 10327
rect 12651 10275 12697 10327
rect 12711 10275 12757 10327
rect 12757 10275 12763 10327
rect 12645 10208 12651 10260
rect 12651 10208 12697 10260
rect 12711 10208 12757 10260
rect 12757 10208 12763 10260
rect 12645 8714 12697 8720
rect 12645 8680 12651 8714
rect 12651 8680 12685 8714
rect 12685 8680 12697 8714
rect 12645 8668 12697 8680
rect 12711 8714 12763 8720
rect 12711 8680 12723 8714
rect 12723 8680 12757 8714
rect 12757 8680 12763 8714
rect 12711 8668 12763 8680
rect 12645 8641 12697 8654
rect 12645 8607 12651 8641
rect 12651 8607 12685 8641
rect 12685 8607 12697 8641
rect 12645 8602 12697 8607
rect 12711 8641 12763 8654
rect 12711 8607 12723 8641
rect 12723 8607 12757 8641
rect 12757 8607 12763 8641
rect 12711 8602 12763 8607
rect 12645 8568 12697 8588
rect 12645 8536 12651 8568
rect 12651 8536 12685 8568
rect 12685 8536 12697 8568
rect 12711 8568 12763 8588
rect 12711 8536 12723 8568
rect 12723 8536 12757 8568
rect 12757 8536 12763 8568
rect 12645 8495 12697 8522
rect 12645 8470 12651 8495
rect 12651 8470 12685 8495
rect 12685 8470 12697 8495
rect 12711 8495 12763 8522
rect 12711 8470 12723 8495
rect 12723 8470 12757 8495
rect 12757 8470 12763 8495
rect 12645 8422 12697 8456
rect 12711 8422 12763 8456
rect 12645 8404 12651 8422
rect 12651 8404 12697 8422
rect 12711 8404 12757 8422
rect 12757 8404 12763 8422
rect 12645 8338 12651 8390
rect 12651 8338 12697 8390
rect 12711 8338 12757 8390
rect 12757 8338 12763 8390
rect 12645 8271 12651 8323
rect 12651 8271 12697 8323
rect 12711 8271 12757 8323
rect 12757 8271 12763 8323
rect 12645 8204 12651 8256
rect 12651 8204 12697 8256
rect 12711 8204 12757 8256
rect 12757 8204 12763 8256
rect 12645 6714 12697 6724
rect 12645 6680 12651 6714
rect 12651 6680 12685 6714
rect 12685 6680 12697 6714
rect 12645 6672 12697 6680
rect 12711 6714 12763 6724
rect 12711 6680 12723 6714
rect 12723 6680 12757 6714
rect 12757 6680 12763 6714
rect 12711 6672 12763 6680
rect 12645 6641 12697 6658
rect 12645 6607 12651 6641
rect 12651 6607 12685 6641
rect 12685 6607 12697 6641
rect 12645 6606 12697 6607
rect 12711 6641 12763 6658
rect 12711 6607 12723 6641
rect 12723 6607 12757 6641
rect 12757 6607 12763 6641
rect 12711 6606 12763 6607
rect 12645 6568 12697 6592
rect 12645 6540 12651 6568
rect 12651 6540 12685 6568
rect 12685 6540 12697 6568
rect 12711 6568 12763 6592
rect 12711 6540 12723 6568
rect 12723 6540 12757 6568
rect 12757 6540 12763 6568
rect 12645 6495 12697 6526
rect 12645 6474 12651 6495
rect 12651 6474 12685 6495
rect 12685 6474 12697 6495
rect 12711 6495 12763 6526
rect 12711 6474 12723 6495
rect 12723 6474 12757 6495
rect 12757 6474 12763 6495
rect 12645 6422 12697 6460
rect 12711 6422 12763 6460
rect 12645 6408 12651 6422
rect 12651 6408 12697 6422
rect 12711 6408 12757 6422
rect 12757 6408 12763 6422
rect 12645 6342 12651 6394
rect 12651 6342 12697 6394
rect 12711 6342 12757 6394
rect 12757 6342 12763 6394
rect 12645 6275 12651 6327
rect 12651 6275 12697 6327
rect 12711 6275 12757 6327
rect 12757 6275 12763 6327
rect 12645 6208 12651 6260
rect 12651 6208 12697 6260
rect 12711 6208 12757 6260
rect 12757 6208 12763 6260
rect 12922 13877 12974 13892
rect 12922 13843 12928 13877
rect 12928 13843 12962 13877
rect 12962 13843 12974 13877
rect 12922 13840 12974 13843
rect 12988 13877 13040 13892
rect 12988 13843 13000 13877
rect 13000 13843 13034 13877
rect 13034 13843 13040 13877
rect 12988 13840 13040 13843
rect 12922 13799 12974 13826
rect 12922 13774 12928 13799
rect 12928 13774 12962 13799
rect 12962 13774 12974 13799
rect 12988 13799 13040 13826
rect 12988 13774 13000 13799
rect 13000 13774 13034 13799
rect 13034 13774 13040 13799
rect 12922 13722 12974 13760
rect 12922 13708 12928 13722
rect 12928 13708 12962 13722
rect 12962 13708 12974 13722
rect 12988 13722 13040 13760
rect 12988 13708 13000 13722
rect 13000 13708 13034 13722
rect 13034 13708 13040 13722
rect 12922 13688 12928 13694
rect 12928 13688 12962 13694
rect 12962 13688 12974 13694
rect 12922 13645 12974 13688
rect 12922 13642 12928 13645
rect 12928 13642 12962 13645
rect 12962 13642 12974 13645
rect 12988 13688 13000 13694
rect 13000 13688 13034 13694
rect 13034 13688 13040 13694
rect 12988 13645 13040 13688
rect 12988 13642 13000 13645
rect 13000 13642 13034 13645
rect 13034 13642 13040 13645
rect 12922 13611 12928 13628
rect 12928 13611 12962 13628
rect 12962 13611 12974 13628
rect 12922 13576 12974 13611
rect 12988 13611 13000 13628
rect 13000 13611 13034 13628
rect 13034 13611 13040 13628
rect 12988 13576 13040 13611
rect 12922 13534 12928 13562
rect 12928 13534 12962 13562
rect 12962 13534 12974 13562
rect 12922 13510 12974 13534
rect 12988 13534 13000 13562
rect 13000 13534 13034 13562
rect 13034 13534 13040 13562
rect 12988 13510 13040 13534
rect 12922 13491 12974 13495
rect 12922 13457 12928 13491
rect 12928 13457 12962 13491
rect 12962 13457 12974 13491
rect 12922 13443 12974 13457
rect 12988 13491 13040 13495
rect 12988 13457 13000 13491
rect 13000 13457 13034 13491
rect 13034 13457 13040 13491
rect 12988 13443 13040 13457
rect 12922 13414 12974 13428
rect 12922 13380 12928 13414
rect 12928 13380 12962 13414
rect 12962 13380 12974 13414
rect 12922 13376 12974 13380
rect 12988 13414 13040 13428
rect 12988 13380 13000 13414
rect 13000 13380 13034 13414
rect 13034 13380 13040 13414
rect 12988 13376 13040 13380
rect 12922 11840 12928 11892
rect 12928 11840 12974 11892
rect 12988 11840 13034 11892
rect 13034 11840 13040 11892
rect 12922 11774 12928 11826
rect 12928 11774 12974 11826
rect 12988 11774 13034 11826
rect 13034 11774 13040 11826
rect 12922 11708 12928 11760
rect 12928 11708 12974 11760
rect 12988 11708 13034 11760
rect 13034 11708 13040 11760
rect 12922 11642 12928 11694
rect 12928 11642 12974 11694
rect 12988 11642 13034 11694
rect 13034 11642 13040 11694
rect 12922 11576 12928 11628
rect 12928 11576 12974 11628
rect 12988 11576 13034 11628
rect 13034 11576 13040 11628
rect 12922 11510 12928 11562
rect 12928 11510 12974 11562
rect 12988 11510 13034 11562
rect 13034 11510 13040 11562
rect 12922 11443 12928 11495
rect 12928 11443 12974 11495
rect 12988 11443 13034 11495
rect 13034 11443 13040 11495
rect 12922 11380 12928 11428
rect 12928 11380 12974 11428
rect 12988 11380 13034 11428
rect 13034 11380 13040 11428
rect 12922 11376 12974 11380
rect 12988 11376 13040 11380
rect 12922 9844 12928 9896
rect 12928 9844 12974 9896
rect 12988 9844 13034 9896
rect 13034 9844 13040 9896
rect 12922 9778 12928 9830
rect 12928 9778 12974 9830
rect 12988 9778 13034 9830
rect 13034 9778 13040 9830
rect 12922 9712 12928 9764
rect 12928 9712 12974 9764
rect 12988 9712 13034 9764
rect 13034 9712 13040 9764
rect 12922 9646 12928 9698
rect 12928 9646 12974 9698
rect 12988 9646 13034 9698
rect 13034 9646 13040 9698
rect 12922 9580 12928 9632
rect 12928 9580 12974 9632
rect 12988 9580 13034 9632
rect 13034 9580 13040 9632
rect 12922 9514 12928 9566
rect 12928 9514 12974 9566
rect 12988 9514 13034 9566
rect 13034 9514 13040 9566
rect 12922 9447 12928 9499
rect 12928 9447 12974 9499
rect 12988 9447 13034 9499
rect 13034 9447 13040 9499
rect 12922 9380 12928 9432
rect 12928 9380 12974 9432
rect 12988 9380 13034 9432
rect 13034 9380 13040 9432
rect 12922 7839 12928 7891
rect 12928 7839 12974 7891
rect 12988 7839 13034 7891
rect 13034 7839 13040 7891
rect 12922 7773 12928 7825
rect 12928 7773 12974 7825
rect 12988 7773 13034 7825
rect 13034 7773 13040 7825
rect 12922 7707 12928 7759
rect 12928 7707 12974 7759
rect 12988 7707 13034 7759
rect 13034 7707 13040 7759
rect 12922 7641 12928 7693
rect 12928 7641 12974 7693
rect 12988 7641 13034 7693
rect 13034 7641 13040 7693
rect 12922 7575 12928 7627
rect 12928 7575 12974 7627
rect 12988 7575 13034 7627
rect 13034 7575 13040 7627
rect 12922 7509 12928 7561
rect 12928 7509 12974 7561
rect 12988 7509 13034 7561
rect 13034 7509 13040 7561
rect 12922 7442 12928 7494
rect 12928 7442 12974 7494
rect 12988 7442 13034 7494
rect 13034 7442 13040 7494
rect 12922 7380 12928 7427
rect 12928 7380 12974 7427
rect 12988 7380 13034 7427
rect 13034 7380 13040 7427
rect 12922 7375 12974 7380
rect 12988 7375 13040 7380
rect 12922 5842 12928 5894
rect 12928 5842 12974 5894
rect 12988 5842 13034 5894
rect 13034 5842 13040 5894
rect 12922 5776 12928 5828
rect 12928 5776 12974 5828
rect 12988 5776 13034 5828
rect 13034 5776 13040 5828
rect 12922 5710 12928 5762
rect 12928 5710 12974 5762
rect 12988 5710 13034 5762
rect 13034 5710 13040 5762
rect 12922 5644 12928 5696
rect 12928 5644 12974 5696
rect 12988 5644 13034 5696
rect 13034 5644 13040 5696
rect 12922 5578 12928 5630
rect 12928 5578 12974 5630
rect 12988 5578 13034 5630
rect 13034 5578 13040 5630
rect 12922 5512 12928 5564
rect 12928 5512 12974 5564
rect 12988 5512 13034 5564
rect 13034 5512 13040 5564
rect 12922 5445 12928 5497
rect 12928 5445 12974 5497
rect 12988 5445 13034 5497
rect 13034 5445 13040 5497
rect 12922 5380 12928 5430
rect 12928 5380 12974 5430
rect 12988 5380 13034 5430
rect 13034 5380 13040 5430
rect 13200 14345 13252 14394
rect 13200 14342 13205 14345
rect 13205 14342 13239 14345
rect 13239 14342 13252 14345
rect 13270 14345 13322 14394
rect 13270 14342 13277 14345
rect 13277 14342 13311 14345
rect 13311 14342 13322 14345
rect 13340 14342 13392 14394
rect 13410 14342 13462 14394
rect 13480 14342 13490 14394
rect 13490 14342 13532 14394
rect 13550 14342 13596 14394
rect 13596 14342 13602 14394
rect 13200 14311 13205 14330
rect 13205 14311 13239 14330
rect 13239 14311 13252 14330
rect 13200 14278 13252 14311
rect 13270 14311 13277 14330
rect 13277 14311 13311 14330
rect 13311 14311 13322 14330
rect 13270 14278 13322 14311
rect 13340 14278 13392 14330
rect 13410 14278 13462 14330
rect 13480 14278 13490 14330
rect 13490 14278 13532 14330
rect 13550 14278 13596 14330
rect 13596 14278 13602 14330
rect 13200 14233 13205 14266
rect 13205 14233 13239 14266
rect 13239 14233 13252 14266
rect 13200 14214 13252 14233
rect 13270 14233 13277 14266
rect 13277 14233 13311 14266
rect 13311 14233 13322 14266
rect 13270 14214 13322 14233
rect 13340 14214 13392 14266
rect 13410 14214 13462 14266
rect 13480 14214 13490 14266
rect 13490 14214 13532 14266
rect 13550 14214 13596 14266
rect 13596 14214 13602 14266
rect 13200 14189 13252 14202
rect 13200 14155 13205 14189
rect 13205 14155 13239 14189
rect 13239 14155 13252 14189
rect 13200 14150 13252 14155
rect 13270 14189 13322 14202
rect 13270 14155 13277 14189
rect 13277 14155 13311 14189
rect 13311 14155 13322 14189
rect 13270 14150 13322 14155
rect 13340 14150 13392 14202
rect 13410 14150 13462 14202
rect 13480 14150 13490 14202
rect 13490 14150 13532 14202
rect 13550 14150 13596 14202
rect 13596 14150 13602 14202
rect 13200 14111 13252 14138
rect 13200 14086 13205 14111
rect 13205 14086 13239 14111
rect 13239 14086 13252 14111
rect 13270 14111 13322 14138
rect 13270 14086 13277 14111
rect 13277 14086 13311 14111
rect 13311 14086 13322 14111
rect 13340 14086 13392 14138
rect 13410 14086 13462 14138
rect 13480 14086 13490 14138
rect 13490 14086 13532 14138
rect 13550 14086 13596 14138
rect 13596 14086 13602 14138
rect 13200 14033 13252 14074
rect 13200 14022 13205 14033
rect 13205 14022 13239 14033
rect 13239 14022 13252 14033
rect 13270 14033 13322 14074
rect 13270 14022 13277 14033
rect 13277 14022 13311 14033
rect 13311 14022 13322 14033
rect 13340 14022 13392 14074
rect 13410 14022 13462 14074
rect 13480 14022 13490 14074
rect 13490 14022 13532 14074
rect 13550 14022 13596 14074
rect 13596 14022 13602 14074
rect 13200 13999 13205 14010
rect 13205 13999 13239 14010
rect 13239 13999 13252 14010
rect 13200 13958 13252 13999
rect 13270 13999 13277 14010
rect 13277 13999 13311 14010
rect 13311 13999 13322 14010
rect 13270 13958 13322 13999
rect 13340 13958 13392 14010
rect 13410 13958 13462 14010
rect 13480 13958 13490 14010
rect 13490 13958 13532 14010
rect 13550 13958 13596 14010
rect 13596 13958 13602 14010
rect 13200 13921 13205 13946
rect 13205 13921 13239 13946
rect 13239 13921 13252 13946
rect 13200 13894 13252 13921
rect 13270 13921 13277 13946
rect 13277 13921 13311 13946
rect 13311 13921 13322 13946
rect 13270 13894 13322 13921
rect 13340 13894 13392 13946
rect 13410 13894 13462 13946
rect 13480 13894 13490 13946
rect 13490 13894 13532 13946
rect 13550 13894 13596 13946
rect 13596 13894 13602 13946
rect 13200 13877 13252 13882
rect 13200 13843 13205 13877
rect 13205 13843 13239 13877
rect 13239 13843 13252 13877
rect 13200 13830 13252 13843
rect 13270 13877 13322 13882
rect 13270 13843 13277 13877
rect 13277 13843 13311 13877
rect 13311 13843 13322 13877
rect 13270 13830 13322 13843
rect 13340 13830 13392 13882
rect 13410 13830 13462 13882
rect 13480 13830 13490 13882
rect 13490 13830 13532 13882
rect 13550 13830 13596 13882
rect 13596 13830 13602 13882
rect 13200 13799 13252 13818
rect 13200 13766 13205 13799
rect 13205 13766 13239 13799
rect 13239 13766 13252 13799
rect 13270 13799 13322 13818
rect 13270 13766 13277 13799
rect 13277 13766 13311 13799
rect 13311 13766 13322 13799
rect 13340 13766 13392 13818
rect 13410 13766 13462 13818
rect 13480 13766 13490 13818
rect 13490 13766 13532 13818
rect 13550 13766 13596 13818
rect 13596 13766 13602 13818
rect 13200 13722 13252 13754
rect 13200 13702 13205 13722
rect 13205 13702 13239 13722
rect 13239 13702 13252 13722
rect 13270 13722 13322 13754
rect 13270 13702 13277 13722
rect 13277 13702 13311 13722
rect 13311 13702 13322 13722
rect 13340 13702 13392 13754
rect 13410 13702 13462 13754
rect 13480 13702 13490 13754
rect 13490 13702 13532 13754
rect 13550 13702 13596 13754
rect 13596 13702 13602 13754
rect 13200 13688 13205 13690
rect 13205 13688 13239 13690
rect 13239 13688 13252 13690
rect 13200 13645 13252 13688
rect 13200 13638 13205 13645
rect 13205 13638 13239 13645
rect 13239 13638 13252 13645
rect 13270 13688 13277 13690
rect 13277 13688 13311 13690
rect 13311 13688 13322 13690
rect 13270 13645 13322 13688
rect 13270 13638 13277 13645
rect 13277 13638 13311 13645
rect 13311 13638 13322 13645
rect 13340 13638 13392 13690
rect 13410 13638 13462 13690
rect 13480 13638 13490 13690
rect 13490 13638 13532 13690
rect 13550 13638 13596 13690
rect 13596 13638 13602 13690
rect 13200 13611 13205 13626
rect 13205 13611 13239 13626
rect 13239 13611 13252 13626
rect 13200 13574 13252 13611
rect 13270 13611 13277 13626
rect 13277 13611 13311 13626
rect 13311 13611 13322 13626
rect 13270 13574 13322 13611
rect 13340 13574 13392 13626
rect 13410 13574 13462 13626
rect 13480 13574 13490 13626
rect 13490 13574 13532 13626
rect 13550 13574 13596 13626
rect 13596 13574 13602 13626
rect 13200 13534 13205 13562
rect 13205 13534 13239 13562
rect 13239 13534 13252 13562
rect 13200 13510 13252 13534
rect 13270 13534 13277 13562
rect 13277 13534 13311 13562
rect 13311 13534 13322 13562
rect 13270 13510 13322 13534
rect 13340 13510 13392 13562
rect 13410 13510 13462 13562
rect 13480 13510 13490 13562
rect 13490 13510 13532 13562
rect 13550 13510 13596 13562
rect 13596 13510 13602 13562
rect 13200 13491 13252 13498
rect 13200 13457 13205 13491
rect 13205 13457 13239 13491
rect 13239 13457 13252 13491
rect 13200 13446 13252 13457
rect 13270 13491 13322 13498
rect 13270 13457 13277 13491
rect 13277 13457 13311 13491
rect 13311 13457 13322 13491
rect 13270 13446 13322 13457
rect 13340 13446 13392 13498
rect 13410 13446 13462 13498
rect 13480 13446 13490 13498
rect 13490 13446 13532 13498
rect 13550 13446 13596 13498
rect 13596 13446 13602 13498
rect 13200 13414 13252 13434
rect 13200 13382 13205 13414
rect 13205 13382 13239 13414
rect 13239 13382 13252 13414
rect 13270 13414 13322 13434
rect 13270 13382 13277 13414
rect 13277 13382 13311 13414
rect 13311 13382 13322 13414
rect 13340 13382 13392 13434
rect 13410 13382 13462 13434
rect 13480 13382 13490 13434
rect 13490 13382 13532 13434
rect 13550 13382 13596 13434
rect 13596 13382 13602 13434
rect 13200 13318 13252 13370
rect 13270 13318 13322 13370
rect 13340 13318 13392 13370
rect 13410 13318 13462 13370
rect 13480 13318 13490 13370
rect 13490 13318 13532 13370
rect 13550 13318 13596 13370
rect 13596 13318 13602 13370
rect 13200 13254 13252 13306
rect 13270 13254 13322 13306
rect 13340 13254 13392 13306
rect 13410 13254 13462 13306
rect 13480 13254 13490 13306
rect 13490 13254 13532 13306
rect 13550 13254 13596 13306
rect 13596 13254 13602 13306
rect 13200 13190 13252 13242
rect 13270 13190 13322 13242
rect 13340 13190 13392 13242
rect 13410 13190 13462 13242
rect 13480 13190 13490 13242
rect 13490 13190 13532 13242
rect 13550 13190 13596 13242
rect 13596 13190 13602 13242
rect 13200 13126 13252 13178
rect 13270 13126 13322 13178
rect 13340 13126 13392 13178
rect 13410 13126 13462 13178
rect 13480 13126 13490 13178
rect 13490 13126 13532 13178
rect 13550 13126 13596 13178
rect 13596 13126 13602 13178
rect 13200 13062 13252 13114
rect 13270 13062 13322 13114
rect 13340 13062 13392 13114
rect 13410 13062 13462 13114
rect 13480 13062 13490 13114
rect 13490 13062 13532 13114
rect 13550 13062 13596 13114
rect 13596 13062 13602 13114
rect 13200 12998 13252 13050
rect 13270 12998 13322 13050
rect 13340 12998 13392 13050
rect 13410 12998 13462 13050
rect 13480 12998 13490 13050
rect 13490 12998 13532 13050
rect 13550 12998 13596 13050
rect 13596 12998 13602 13050
rect 13200 12934 13252 12986
rect 13270 12934 13322 12986
rect 13340 12934 13392 12986
rect 13410 12934 13462 12986
rect 13480 12934 13490 12986
rect 13490 12934 13532 12986
rect 13550 12934 13596 12986
rect 13596 12934 13602 12986
rect 13200 12870 13252 12922
rect 13270 12870 13322 12922
rect 13340 12870 13392 12922
rect 13410 12870 13462 12922
rect 13480 12870 13490 12922
rect 13490 12870 13532 12922
rect 13550 12870 13596 12922
rect 13596 12870 13602 12922
rect 13200 12806 13252 12858
rect 13270 12806 13322 12858
rect 13340 12806 13392 12858
rect 13410 12806 13462 12858
rect 13480 12806 13490 12858
rect 13490 12806 13532 12858
rect 13550 12806 13596 12858
rect 13596 12806 13602 12858
rect 13200 12742 13252 12794
rect 13270 12742 13322 12794
rect 13340 12742 13392 12794
rect 13410 12742 13462 12794
rect 13480 12742 13490 12794
rect 13490 12742 13532 12794
rect 13550 12742 13596 12794
rect 13596 12742 13602 12794
rect 13200 12714 13252 12730
rect 13200 12680 13205 12714
rect 13205 12680 13239 12714
rect 13239 12680 13252 12714
rect 13200 12678 13252 12680
rect 13270 12714 13322 12730
rect 13270 12680 13277 12714
rect 13277 12680 13311 12714
rect 13311 12680 13322 12714
rect 13270 12678 13322 12680
rect 13340 12678 13392 12730
rect 13410 12678 13462 12730
rect 13480 12678 13490 12730
rect 13490 12678 13532 12730
rect 13550 12678 13596 12730
rect 13596 12678 13602 12730
rect 13200 12641 13252 12666
rect 13200 12614 13205 12641
rect 13205 12614 13239 12641
rect 13239 12614 13252 12641
rect 13270 12641 13322 12666
rect 13270 12614 13277 12641
rect 13277 12614 13311 12641
rect 13311 12614 13322 12641
rect 13340 12614 13392 12666
rect 13410 12614 13462 12666
rect 13480 12614 13490 12666
rect 13490 12614 13532 12666
rect 13550 12614 13596 12666
rect 13596 12614 13602 12666
rect 13200 12568 13252 12602
rect 13200 12550 13205 12568
rect 13205 12550 13239 12568
rect 13239 12550 13252 12568
rect 13270 12568 13322 12602
rect 13270 12550 13277 12568
rect 13277 12550 13311 12568
rect 13311 12550 13322 12568
rect 13340 12550 13392 12602
rect 13410 12550 13462 12602
rect 13480 12550 13490 12602
rect 13490 12550 13532 12602
rect 13550 12550 13596 12602
rect 13596 12550 13602 12602
rect 13200 12534 13205 12538
rect 13205 12534 13239 12538
rect 13239 12534 13252 12538
rect 13200 12495 13252 12534
rect 13200 12486 13205 12495
rect 13205 12486 13239 12495
rect 13239 12486 13252 12495
rect 13270 12534 13277 12538
rect 13277 12534 13311 12538
rect 13311 12534 13322 12538
rect 13270 12495 13322 12534
rect 13270 12486 13277 12495
rect 13277 12486 13311 12495
rect 13311 12486 13322 12495
rect 13340 12486 13392 12538
rect 13410 12486 13462 12538
rect 13480 12486 13490 12538
rect 13490 12486 13532 12538
rect 13550 12486 13596 12538
rect 13596 12486 13602 12538
rect 13200 12461 13205 12474
rect 13205 12461 13239 12474
rect 13239 12461 13252 12474
rect 13200 12422 13252 12461
rect 13270 12461 13277 12474
rect 13277 12461 13311 12474
rect 13311 12461 13322 12474
rect 13270 12422 13322 12461
rect 13340 12422 13392 12474
rect 13410 12422 13462 12474
rect 13480 12422 13490 12474
rect 13490 12422 13532 12474
rect 13550 12422 13596 12474
rect 13596 12422 13602 12474
rect 13200 12358 13205 12410
rect 13205 12358 13252 12410
rect 13270 12358 13311 12410
rect 13311 12358 13322 12410
rect 13340 12358 13392 12410
rect 13410 12358 13462 12410
rect 13480 12358 13490 12410
rect 13490 12358 13532 12410
rect 13550 12358 13596 12410
rect 13596 12358 13602 12410
rect 13200 12294 13205 12346
rect 13205 12294 13252 12346
rect 13270 12294 13311 12346
rect 13311 12294 13322 12346
rect 13340 12294 13392 12346
rect 13410 12294 13462 12346
rect 13480 12294 13490 12346
rect 13490 12294 13532 12346
rect 13550 12294 13596 12346
rect 13596 12294 13602 12346
rect 13200 12230 13205 12282
rect 13205 12230 13252 12282
rect 13270 12230 13311 12282
rect 13311 12230 13322 12282
rect 13340 12230 13392 12282
rect 13410 12230 13462 12282
rect 13480 12230 13490 12282
rect 13490 12230 13532 12282
rect 13550 12230 13596 12282
rect 13596 12230 13602 12282
rect 13200 12166 13205 12218
rect 13205 12166 13252 12218
rect 13270 12166 13311 12218
rect 13311 12166 13322 12218
rect 13340 12166 13392 12218
rect 13410 12166 13462 12218
rect 13480 12166 13490 12218
rect 13490 12166 13532 12218
rect 13550 12166 13596 12218
rect 13596 12166 13602 12218
rect 13200 12102 13205 12154
rect 13205 12102 13252 12154
rect 13270 12102 13311 12154
rect 13311 12102 13322 12154
rect 13340 12102 13392 12154
rect 13410 12102 13462 12154
rect 13480 12102 13490 12154
rect 13490 12102 13532 12154
rect 13550 12102 13596 12154
rect 13596 12102 13602 12154
rect 13200 12038 13205 12090
rect 13205 12038 13252 12090
rect 13270 12038 13311 12090
rect 13311 12038 13322 12090
rect 13340 12038 13392 12090
rect 13410 12038 13462 12090
rect 13480 12038 13490 12090
rect 13490 12038 13532 12090
rect 13550 12038 13596 12090
rect 13596 12038 13602 12090
rect 13200 11974 13205 12026
rect 13205 11974 13252 12026
rect 13270 11974 13311 12026
rect 13311 11974 13322 12026
rect 13340 11974 13392 12026
rect 13410 11974 13462 12026
rect 13480 11974 13490 12026
rect 13490 11974 13532 12026
rect 13550 11974 13596 12026
rect 13596 11974 13602 12026
rect 13200 11910 13205 11962
rect 13205 11910 13252 11962
rect 13270 11910 13311 11962
rect 13311 11910 13322 11962
rect 13340 11910 13392 11962
rect 13410 11910 13462 11962
rect 13480 11910 13490 11962
rect 13490 11910 13532 11962
rect 13550 11910 13596 11962
rect 13596 11910 13602 11962
rect 13200 11846 13205 11898
rect 13205 11846 13252 11898
rect 13270 11846 13311 11898
rect 13311 11846 13322 11898
rect 13340 11846 13392 11898
rect 13410 11846 13462 11898
rect 13480 11846 13490 11898
rect 13490 11846 13532 11898
rect 13550 11846 13596 11898
rect 13596 11846 13602 11898
rect 13200 11782 13205 11834
rect 13205 11782 13252 11834
rect 13270 11782 13311 11834
rect 13311 11782 13322 11834
rect 13340 11782 13392 11834
rect 13410 11782 13462 11834
rect 13480 11782 13490 11834
rect 13490 11782 13532 11834
rect 13550 11782 13596 11834
rect 13596 11782 13602 11834
rect 13200 11718 13205 11770
rect 13205 11718 13252 11770
rect 13270 11718 13311 11770
rect 13311 11718 13322 11770
rect 13340 11718 13392 11770
rect 13410 11718 13462 11770
rect 13480 11718 13490 11770
rect 13490 11718 13532 11770
rect 13550 11718 13596 11770
rect 13596 11718 13602 11770
rect 13200 11654 13205 11706
rect 13205 11654 13252 11706
rect 13270 11654 13311 11706
rect 13311 11654 13322 11706
rect 13340 11654 13392 11706
rect 13410 11654 13462 11706
rect 13480 11654 13490 11706
rect 13490 11654 13532 11706
rect 13550 11654 13596 11706
rect 13596 11654 13602 11706
rect 13200 11590 13205 11642
rect 13205 11590 13252 11642
rect 13270 11590 13311 11642
rect 13311 11590 13322 11642
rect 13340 11590 13392 11642
rect 13410 11590 13462 11642
rect 13480 11590 13490 11642
rect 13490 11590 13532 11642
rect 13550 11590 13596 11642
rect 13596 11590 13602 11642
rect 13200 11526 13205 11578
rect 13205 11526 13252 11578
rect 13270 11526 13311 11578
rect 13311 11526 13322 11578
rect 13340 11526 13392 11578
rect 13410 11526 13462 11578
rect 13480 11526 13490 11578
rect 13490 11526 13532 11578
rect 13550 11526 13596 11578
rect 13596 11526 13602 11578
rect 13200 11462 13205 11514
rect 13205 11462 13252 11514
rect 13270 11462 13311 11514
rect 13311 11462 13322 11514
rect 13340 11462 13392 11514
rect 13410 11462 13462 11514
rect 13480 11462 13490 11514
rect 13490 11462 13532 11514
rect 13550 11462 13596 11514
rect 13596 11462 13602 11514
rect 13200 11398 13205 11450
rect 13205 11398 13252 11450
rect 13270 11398 13311 11450
rect 13311 11398 13322 11450
rect 13340 11398 13392 11450
rect 13410 11398 13462 11450
rect 13480 11398 13490 11450
rect 13490 11398 13532 11450
rect 13550 11398 13596 11450
rect 13596 11398 13602 11450
rect 13200 11380 13205 11386
rect 13205 11380 13252 11386
rect 13270 11380 13311 11386
rect 13311 11380 13322 11386
rect 13200 11334 13252 11380
rect 13270 11334 13322 11380
rect 13340 11334 13392 11386
rect 13410 11334 13462 11386
rect 13480 11334 13490 11386
rect 13490 11334 13532 11386
rect 13550 11334 13596 11386
rect 13596 11334 13602 11386
rect 13200 11270 13252 11322
rect 13270 11270 13322 11322
rect 13340 11270 13392 11322
rect 13410 11270 13462 11322
rect 13480 11270 13490 11322
rect 13490 11270 13532 11322
rect 13550 11270 13596 11322
rect 13596 11270 13602 11322
rect 13200 11206 13252 11258
rect 13270 11206 13322 11258
rect 13340 11206 13392 11258
rect 13410 11206 13462 11258
rect 13480 11206 13490 11258
rect 13490 11206 13532 11258
rect 13550 11206 13596 11258
rect 13596 11206 13602 11258
rect 13200 11142 13252 11194
rect 13270 11142 13322 11194
rect 13340 11142 13392 11194
rect 13410 11142 13462 11194
rect 13480 11142 13490 11194
rect 13490 11142 13532 11194
rect 13550 11142 13596 11194
rect 13596 11142 13602 11194
rect 13200 11078 13252 11130
rect 13270 11078 13322 11130
rect 13340 11078 13392 11130
rect 13410 11078 13462 11130
rect 13480 11078 13490 11130
rect 13490 11078 13532 11130
rect 13550 11078 13596 11130
rect 13596 11078 13602 11130
rect 13200 11014 13252 11066
rect 13270 11014 13322 11066
rect 13340 11014 13392 11066
rect 13410 11014 13462 11066
rect 13480 11014 13490 11066
rect 13490 11014 13532 11066
rect 13550 11014 13596 11066
rect 13596 11014 13602 11066
rect 13200 10950 13252 11002
rect 13270 10950 13322 11002
rect 13340 10950 13392 11002
rect 13410 10950 13462 11002
rect 13480 10950 13490 11002
rect 13490 10950 13532 11002
rect 13550 10950 13596 11002
rect 13596 10950 13602 11002
rect 13200 10886 13252 10938
rect 13270 10886 13322 10938
rect 13340 10886 13392 10938
rect 13410 10886 13462 10938
rect 13480 10886 13490 10938
rect 13490 10886 13532 10938
rect 13550 10886 13596 10938
rect 13596 10886 13602 10938
rect 13200 10822 13252 10874
rect 13270 10822 13322 10874
rect 13340 10822 13392 10874
rect 13410 10822 13462 10874
rect 13480 10822 13490 10874
rect 13490 10822 13532 10874
rect 13550 10822 13596 10874
rect 13596 10822 13602 10874
rect 13200 10758 13252 10810
rect 13270 10758 13322 10810
rect 13340 10758 13392 10810
rect 13410 10758 13462 10810
rect 13480 10758 13490 10810
rect 13490 10758 13532 10810
rect 13550 10758 13596 10810
rect 13596 10758 13602 10810
rect 13200 10714 13252 10746
rect 13200 10694 13205 10714
rect 13205 10694 13239 10714
rect 13239 10694 13252 10714
rect 13270 10714 13322 10746
rect 13270 10694 13277 10714
rect 13277 10694 13311 10714
rect 13311 10694 13322 10714
rect 13340 10694 13392 10746
rect 13410 10694 13462 10746
rect 13480 10694 13490 10746
rect 13490 10694 13532 10746
rect 13550 10694 13596 10746
rect 13596 10694 13602 10746
rect 13200 10680 13205 10682
rect 13205 10680 13239 10682
rect 13239 10680 13252 10682
rect 13200 10641 13252 10680
rect 13200 10630 13205 10641
rect 13205 10630 13239 10641
rect 13239 10630 13252 10641
rect 13270 10680 13277 10682
rect 13277 10680 13311 10682
rect 13311 10680 13322 10682
rect 13270 10641 13322 10680
rect 13270 10630 13277 10641
rect 13277 10630 13311 10641
rect 13311 10630 13322 10641
rect 13340 10630 13392 10682
rect 13410 10630 13462 10682
rect 13480 10630 13490 10682
rect 13490 10630 13532 10682
rect 13550 10630 13596 10682
rect 13596 10630 13602 10682
rect 13200 10607 13205 10618
rect 13205 10607 13239 10618
rect 13239 10607 13252 10618
rect 13200 10568 13252 10607
rect 13200 10566 13205 10568
rect 13205 10566 13239 10568
rect 13239 10566 13252 10568
rect 13270 10607 13277 10618
rect 13277 10607 13311 10618
rect 13311 10607 13322 10618
rect 13270 10568 13322 10607
rect 13270 10566 13277 10568
rect 13277 10566 13311 10568
rect 13311 10566 13322 10568
rect 13340 10566 13392 10618
rect 13410 10566 13462 10618
rect 13480 10566 13490 10618
rect 13490 10566 13532 10618
rect 13550 10566 13596 10618
rect 13596 10566 13602 10618
rect 13200 10534 13205 10554
rect 13205 10534 13239 10554
rect 13239 10534 13252 10554
rect 13200 10502 13252 10534
rect 13270 10534 13277 10554
rect 13277 10534 13311 10554
rect 13311 10534 13322 10554
rect 13270 10502 13322 10534
rect 13340 10502 13392 10554
rect 13410 10502 13462 10554
rect 13480 10502 13490 10554
rect 13490 10502 13532 10554
rect 13550 10502 13596 10554
rect 13596 10502 13602 10554
rect 13200 10461 13205 10490
rect 13205 10461 13239 10490
rect 13239 10461 13252 10490
rect 13200 10438 13252 10461
rect 13270 10461 13277 10490
rect 13277 10461 13311 10490
rect 13311 10461 13322 10490
rect 13270 10438 13322 10461
rect 13340 10438 13392 10490
rect 13410 10438 13462 10490
rect 13480 10438 13490 10490
rect 13490 10438 13532 10490
rect 13550 10438 13596 10490
rect 13596 10438 13602 10490
rect 13200 10422 13252 10426
rect 13270 10422 13322 10426
rect 13200 10374 13205 10422
rect 13205 10374 13252 10422
rect 13270 10374 13311 10422
rect 13311 10374 13322 10422
rect 13340 10374 13392 10426
rect 13410 10374 13462 10426
rect 13480 10374 13490 10426
rect 13490 10374 13532 10426
rect 13550 10374 13596 10426
rect 13596 10374 13602 10426
rect 13200 10310 13205 10362
rect 13205 10310 13252 10362
rect 13270 10310 13311 10362
rect 13311 10310 13322 10362
rect 13340 10310 13392 10362
rect 13410 10310 13462 10362
rect 13480 10310 13490 10362
rect 13490 10310 13532 10362
rect 13550 10310 13596 10362
rect 13596 10310 13602 10362
rect 13200 10246 13205 10298
rect 13205 10246 13252 10298
rect 13270 10246 13311 10298
rect 13311 10246 13322 10298
rect 13340 10246 13392 10298
rect 13410 10246 13462 10298
rect 13480 10246 13490 10298
rect 13490 10246 13532 10298
rect 13550 10246 13596 10298
rect 13596 10246 13602 10298
rect 13200 10182 13205 10234
rect 13205 10182 13252 10234
rect 13270 10182 13311 10234
rect 13311 10182 13322 10234
rect 13340 10182 13392 10234
rect 13410 10182 13462 10234
rect 13480 10182 13490 10234
rect 13490 10182 13532 10234
rect 13550 10182 13596 10234
rect 13596 10182 13602 10234
rect 13200 10118 13205 10170
rect 13205 10118 13252 10170
rect 13270 10118 13311 10170
rect 13311 10118 13322 10170
rect 13340 10118 13392 10170
rect 13410 10118 13462 10170
rect 13480 10118 13490 10170
rect 13490 10118 13532 10170
rect 13550 10118 13596 10170
rect 13596 10118 13602 10170
rect 13200 10054 13205 10106
rect 13205 10054 13252 10106
rect 13270 10054 13311 10106
rect 13311 10054 13322 10106
rect 13340 10054 13392 10106
rect 13410 10054 13462 10106
rect 13480 10054 13490 10106
rect 13490 10054 13532 10106
rect 13550 10054 13596 10106
rect 13596 10054 13602 10106
rect 13200 9990 13205 10042
rect 13205 9990 13252 10042
rect 13270 9990 13311 10042
rect 13311 9990 13322 10042
rect 13340 9990 13392 10042
rect 13410 9990 13462 10042
rect 13480 9990 13490 10042
rect 13490 9990 13532 10042
rect 13550 9990 13596 10042
rect 13596 9990 13602 10042
rect 13200 9926 13205 9978
rect 13205 9926 13252 9978
rect 13270 9926 13311 9978
rect 13311 9926 13322 9978
rect 13340 9926 13392 9978
rect 13410 9926 13462 9978
rect 13480 9926 13490 9978
rect 13490 9926 13532 9978
rect 13550 9926 13596 9978
rect 13596 9926 13602 9978
rect 13200 9862 13205 9914
rect 13205 9862 13252 9914
rect 13270 9862 13311 9914
rect 13311 9862 13322 9914
rect 13340 9862 13392 9914
rect 13410 9862 13462 9914
rect 13480 9862 13490 9914
rect 13490 9862 13532 9914
rect 13550 9862 13596 9914
rect 13596 9862 13602 9914
rect 13200 9798 13205 9850
rect 13205 9798 13252 9850
rect 13270 9798 13311 9850
rect 13311 9798 13322 9850
rect 13340 9798 13392 9850
rect 13410 9798 13462 9850
rect 13480 9798 13490 9850
rect 13490 9798 13532 9850
rect 13550 9798 13596 9850
rect 13596 9798 13602 9850
rect 13200 9734 13205 9786
rect 13205 9734 13252 9786
rect 13270 9734 13311 9786
rect 13311 9734 13322 9786
rect 13340 9734 13392 9786
rect 13410 9734 13462 9786
rect 13480 9734 13490 9786
rect 13490 9734 13532 9786
rect 13550 9734 13596 9786
rect 13596 9734 13602 9786
rect 13200 9670 13205 9722
rect 13205 9670 13252 9722
rect 13270 9670 13311 9722
rect 13311 9670 13322 9722
rect 13340 9670 13392 9722
rect 13410 9670 13462 9722
rect 13480 9670 13490 9722
rect 13490 9670 13532 9722
rect 13550 9670 13596 9722
rect 13596 9670 13602 9722
rect 13200 9606 13205 9658
rect 13205 9606 13252 9658
rect 13270 9606 13311 9658
rect 13311 9606 13322 9658
rect 13340 9606 13392 9658
rect 13410 9606 13462 9658
rect 13480 9606 13490 9658
rect 13490 9606 13532 9658
rect 13550 9606 13596 9658
rect 13596 9606 13602 9658
rect 13200 9542 13205 9594
rect 13205 9542 13252 9594
rect 13270 9542 13311 9594
rect 13311 9542 13322 9594
rect 13340 9542 13392 9594
rect 13410 9542 13462 9594
rect 13480 9542 13490 9594
rect 13490 9542 13532 9594
rect 13550 9542 13596 9594
rect 13596 9542 13602 9594
rect 13200 9478 13205 9530
rect 13205 9478 13252 9530
rect 13270 9478 13311 9530
rect 13311 9478 13322 9530
rect 13340 9478 13392 9530
rect 13410 9478 13462 9530
rect 13480 9478 13490 9530
rect 13490 9478 13532 9530
rect 13550 9478 13596 9530
rect 13596 9478 13602 9530
rect 13200 9414 13205 9466
rect 13205 9414 13252 9466
rect 13270 9414 13311 9466
rect 13311 9414 13322 9466
rect 13340 9414 13392 9466
rect 13410 9414 13462 9466
rect 13480 9414 13490 9466
rect 13490 9414 13532 9466
rect 13550 9414 13596 9466
rect 13596 9414 13602 9466
rect 13200 9380 13205 9402
rect 13205 9380 13252 9402
rect 13270 9380 13311 9402
rect 13311 9380 13322 9402
rect 13200 9350 13252 9380
rect 13270 9350 13322 9380
rect 13340 9350 13392 9402
rect 13410 9350 13462 9402
rect 13480 9350 13490 9402
rect 13490 9350 13532 9402
rect 13550 9350 13596 9402
rect 13596 9350 13602 9402
rect 13200 9286 13252 9338
rect 13270 9286 13322 9338
rect 13340 9286 13392 9338
rect 13410 9286 13462 9338
rect 13480 9286 13490 9338
rect 13490 9286 13532 9338
rect 13550 9286 13596 9338
rect 13596 9286 13602 9338
rect 13200 9222 13252 9274
rect 13270 9222 13322 9274
rect 13340 9222 13392 9274
rect 13410 9222 13462 9274
rect 13480 9222 13490 9274
rect 13490 9222 13532 9274
rect 13550 9222 13596 9274
rect 13596 9222 13602 9274
rect 13200 9158 13252 9210
rect 13270 9158 13322 9210
rect 13340 9158 13392 9210
rect 13410 9158 13462 9210
rect 13480 9158 13490 9210
rect 13490 9158 13532 9210
rect 13550 9158 13596 9210
rect 13596 9158 13602 9210
rect 13200 9094 13252 9146
rect 13270 9094 13322 9146
rect 13340 9094 13392 9146
rect 13410 9094 13462 9146
rect 13480 9094 13490 9146
rect 13490 9094 13532 9146
rect 13550 9094 13596 9146
rect 13596 9094 13602 9146
rect 13200 9030 13252 9082
rect 13270 9030 13322 9082
rect 13340 9030 13392 9082
rect 13410 9030 13462 9082
rect 13480 9030 13490 9082
rect 13490 9030 13532 9082
rect 13550 9030 13596 9082
rect 13596 9030 13602 9082
rect 13200 8966 13252 9018
rect 13270 8966 13322 9018
rect 13340 8966 13392 9018
rect 13410 8966 13462 9018
rect 13480 8966 13490 9018
rect 13490 8966 13532 9018
rect 13550 8966 13596 9018
rect 13596 8966 13602 9018
rect 13200 8902 13252 8954
rect 13270 8902 13322 8954
rect 13340 8902 13392 8954
rect 13410 8902 13462 8954
rect 13480 8902 13490 8954
rect 13490 8902 13532 8954
rect 13550 8902 13596 8954
rect 13596 8902 13602 8954
rect 13200 8838 13252 8890
rect 13270 8838 13322 8890
rect 13340 8838 13392 8890
rect 13410 8838 13462 8890
rect 13480 8838 13490 8890
rect 13490 8838 13532 8890
rect 13550 8838 13596 8890
rect 13596 8838 13602 8890
rect 13200 8774 13252 8826
rect 13270 8774 13322 8826
rect 13340 8774 13392 8826
rect 13410 8774 13462 8826
rect 13480 8774 13490 8826
rect 13490 8774 13532 8826
rect 13550 8774 13596 8826
rect 13596 8774 13602 8826
rect 13200 8714 13252 8762
rect 13200 8710 13205 8714
rect 13205 8710 13239 8714
rect 13239 8710 13252 8714
rect 13270 8714 13322 8762
rect 13270 8710 13277 8714
rect 13277 8710 13311 8714
rect 13311 8710 13322 8714
rect 13340 8710 13392 8762
rect 13410 8710 13462 8762
rect 13480 8710 13490 8762
rect 13490 8710 13532 8762
rect 13550 8710 13596 8762
rect 13596 8710 13602 8762
rect 13200 8680 13205 8698
rect 13205 8680 13239 8698
rect 13239 8680 13252 8698
rect 13200 8646 13252 8680
rect 13270 8680 13277 8698
rect 13277 8680 13311 8698
rect 13311 8680 13322 8698
rect 13270 8646 13322 8680
rect 13340 8646 13392 8698
rect 13410 8646 13462 8698
rect 13480 8646 13490 8698
rect 13490 8646 13532 8698
rect 13550 8646 13596 8698
rect 13596 8646 13602 8698
rect 13200 8607 13205 8634
rect 13205 8607 13239 8634
rect 13239 8607 13252 8634
rect 13200 8582 13252 8607
rect 13270 8607 13277 8634
rect 13277 8607 13311 8634
rect 13311 8607 13322 8634
rect 13270 8582 13322 8607
rect 13340 8582 13392 8634
rect 13410 8582 13462 8634
rect 13480 8582 13490 8634
rect 13490 8582 13532 8634
rect 13550 8582 13596 8634
rect 13596 8582 13602 8634
rect 13200 8568 13252 8570
rect 13200 8534 13205 8568
rect 13205 8534 13239 8568
rect 13239 8534 13252 8568
rect 13200 8518 13252 8534
rect 13270 8568 13322 8570
rect 13270 8534 13277 8568
rect 13277 8534 13311 8568
rect 13311 8534 13322 8568
rect 13270 8518 13322 8534
rect 13340 8518 13392 8570
rect 13410 8518 13462 8570
rect 13480 8518 13490 8570
rect 13490 8518 13532 8570
rect 13550 8518 13596 8570
rect 13596 8518 13602 8570
rect 13200 8495 13252 8506
rect 13200 8461 13205 8495
rect 13205 8461 13239 8495
rect 13239 8461 13252 8495
rect 13200 8454 13252 8461
rect 13270 8495 13322 8506
rect 13270 8461 13277 8495
rect 13277 8461 13311 8495
rect 13311 8461 13322 8495
rect 13270 8454 13322 8461
rect 13340 8454 13392 8506
rect 13410 8454 13462 8506
rect 13480 8454 13490 8506
rect 13490 8454 13532 8506
rect 13550 8454 13596 8506
rect 13596 8454 13602 8506
rect 13200 8422 13252 8442
rect 13270 8422 13322 8442
rect 13200 8390 13205 8422
rect 13205 8390 13252 8422
rect 13270 8390 13311 8422
rect 13311 8390 13322 8422
rect 13340 8390 13392 8442
rect 13410 8390 13462 8442
rect 13480 8390 13490 8442
rect 13490 8390 13532 8442
rect 13550 8390 13596 8442
rect 13596 8390 13602 8442
rect 13200 8326 13205 8378
rect 13205 8326 13252 8378
rect 13270 8326 13311 8378
rect 13311 8326 13322 8378
rect 13340 8326 13392 8378
rect 13410 8326 13462 8378
rect 13480 8326 13490 8378
rect 13490 8326 13532 8378
rect 13550 8326 13596 8378
rect 13596 8326 13602 8378
rect 13200 8262 13205 8314
rect 13205 8262 13252 8314
rect 13270 8262 13311 8314
rect 13311 8262 13322 8314
rect 13340 8262 13392 8314
rect 13410 8262 13462 8314
rect 13480 8262 13490 8314
rect 13490 8262 13532 8314
rect 13550 8262 13596 8314
rect 13596 8262 13602 8314
rect 13200 8198 13205 8250
rect 13205 8198 13252 8250
rect 13270 8198 13311 8250
rect 13311 8198 13322 8250
rect 13340 8198 13392 8250
rect 13410 8198 13462 8250
rect 13480 8198 13490 8250
rect 13490 8198 13532 8250
rect 13550 8198 13596 8250
rect 13596 8198 13602 8250
rect 13200 8134 13205 8186
rect 13205 8134 13252 8186
rect 13270 8134 13311 8186
rect 13311 8134 13322 8186
rect 13340 8134 13392 8186
rect 13410 8134 13462 8186
rect 13480 8134 13490 8186
rect 13490 8134 13532 8186
rect 13550 8134 13596 8186
rect 13596 8134 13602 8186
rect 13200 8070 13205 8122
rect 13205 8070 13252 8122
rect 13270 8070 13311 8122
rect 13311 8070 13322 8122
rect 13340 8070 13392 8122
rect 13410 8070 13462 8122
rect 13480 8070 13490 8122
rect 13490 8070 13532 8122
rect 13550 8070 13596 8122
rect 13596 8070 13602 8122
rect 13200 8006 13205 8058
rect 13205 8006 13252 8058
rect 13270 8006 13311 8058
rect 13311 8006 13322 8058
rect 13340 8006 13392 8058
rect 13410 8006 13462 8058
rect 13480 8006 13490 8058
rect 13490 8006 13532 8058
rect 13550 8006 13596 8058
rect 13596 8006 13602 8058
rect 13200 7942 13205 7994
rect 13205 7942 13252 7994
rect 13270 7942 13311 7994
rect 13311 7942 13322 7994
rect 13340 7942 13392 7994
rect 13410 7942 13462 7994
rect 13480 7942 13490 7994
rect 13490 7942 13532 7994
rect 13550 7942 13596 7994
rect 13596 7942 13602 7994
rect 13200 7878 13205 7930
rect 13205 7878 13252 7930
rect 13270 7878 13311 7930
rect 13311 7878 13322 7930
rect 13340 7878 13392 7930
rect 13410 7878 13462 7930
rect 13480 7878 13490 7930
rect 13490 7878 13532 7930
rect 13550 7878 13596 7930
rect 13596 7878 13602 7930
rect 13200 7814 13205 7866
rect 13205 7814 13252 7866
rect 13270 7814 13311 7866
rect 13311 7814 13322 7866
rect 13340 7814 13392 7866
rect 13410 7814 13462 7866
rect 13480 7814 13490 7866
rect 13490 7814 13532 7866
rect 13550 7814 13596 7866
rect 13596 7814 13602 7866
rect 13200 7750 13205 7802
rect 13205 7750 13252 7802
rect 13270 7750 13311 7802
rect 13311 7750 13322 7802
rect 13340 7750 13392 7802
rect 13410 7750 13462 7802
rect 13480 7750 13490 7802
rect 13490 7750 13532 7802
rect 13550 7750 13596 7802
rect 13596 7750 13602 7802
rect 13200 7686 13205 7738
rect 13205 7686 13252 7738
rect 13270 7686 13311 7738
rect 13311 7686 13322 7738
rect 13340 7686 13392 7738
rect 13410 7686 13462 7738
rect 13480 7686 13490 7738
rect 13490 7686 13532 7738
rect 13550 7686 13596 7738
rect 13596 7686 13602 7738
rect 13200 7622 13205 7674
rect 13205 7622 13252 7674
rect 13270 7622 13311 7674
rect 13311 7622 13322 7674
rect 13340 7622 13392 7674
rect 13410 7622 13462 7674
rect 13480 7622 13490 7674
rect 13490 7622 13532 7674
rect 13550 7622 13596 7674
rect 13596 7622 13602 7674
rect 13200 7558 13205 7610
rect 13205 7558 13252 7610
rect 13270 7558 13311 7610
rect 13311 7558 13322 7610
rect 13340 7558 13392 7610
rect 13410 7558 13462 7610
rect 13480 7558 13490 7610
rect 13490 7558 13532 7610
rect 13550 7558 13596 7610
rect 13596 7558 13602 7610
rect 13200 7494 13205 7546
rect 13205 7494 13252 7546
rect 13270 7494 13311 7546
rect 13311 7494 13322 7546
rect 13340 7494 13392 7546
rect 13410 7494 13462 7546
rect 13480 7494 13490 7546
rect 13490 7494 13532 7546
rect 13550 7494 13596 7546
rect 13596 7494 13602 7546
rect 13200 7430 13205 7482
rect 13205 7430 13252 7482
rect 13270 7430 13311 7482
rect 13311 7430 13322 7482
rect 13340 7430 13392 7482
rect 13410 7430 13462 7482
rect 13480 7430 13490 7482
rect 13490 7430 13532 7482
rect 13550 7430 13596 7482
rect 13596 7430 13602 7482
rect 13200 7380 13205 7418
rect 13205 7380 13252 7418
rect 13270 7380 13311 7418
rect 13311 7380 13322 7418
rect 13200 7366 13252 7380
rect 13270 7366 13322 7380
rect 13340 7366 13392 7418
rect 13410 7366 13462 7418
rect 13480 7366 13490 7418
rect 13490 7366 13532 7418
rect 13550 7366 13596 7418
rect 13596 7366 13602 7418
rect 13200 7302 13252 7354
rect 13270 7302 13322 7354
rect 13340 7302 13392 7354
rect 13410 7302 13462 7354
rect 13480 7302 13490 7354
rect 13490 7302 13532 7354
rect 13550 7302 13596 7354
rect 13596 7302 13602 7354
rect 13200 7238 13252 7290
rect 13270 7238 13322 7290
rect 13340 7238 13392 7290
rect 13410 7238 13462 7290
rect 13480 7238 13490 7290
rect 13490 7238 13532 7290
rect 13550 7238 13596 7290
rect 13596 7238 13602 7290
rect 13200 7174 13252 7226
rect 13270 7174 13322 7226
rect 13340 7174 13392 7226
rect 13410 7174 13462 7226
rect 13480 7174 13490 7226
rect 13490 7174 13532 7226
rect 13550 7174 13596 7226
rect 13596 7174 13602 7226
rect 13200 7110 13252 7162
rect 13270 7110 13322 7162
rect 13340 7110 13392 7162
rect 13410 7110 13462 7162
rect 13480 7110 13490 7162
rect 13490 7110 13532 7162
rect 13550 7110 13596 7162
rect 13596 7110 13602 7162
rect 13200 7046 13252 7098
rect 13270 7046 13322 7098
rect 13340 7046 13392 7098
rect 13410 7046 13462 7098
rect 13480 7046 13490 7098
rect 13490 7046 13532 7098
rect 13550 7046 13596 7098
rect 13596 7046 13602 7098
rect 13200 6982 13252 7034
rect 13270 6982 13322 7034
rect 13340 6982 13392 7034
rect 13410 6982 13462 7034
rect 13480 6982 13490 7034
rect 13490 6982 13532 7034
rect 13550 6982 13596 7034
rect 13596 6982 13602 7034
rect 13200 6918 13252 6970
rect 13270 6918 13322 6970
rect 13340 6918 13392 6970
rect 13410 6918 13462 6970
rect 13480 6918 13490 6970
rect 13490 6918 13532 6970
rect 13550 6918 13596 6970
rect 13596 6918 13602 6970
rect 13200 6854 13252 6906
rect 13270 6854 13322 6906
rect 13340 6854 13392 6906
rect 13410 6854 13462 6906
rect 13480 6854 13490 6906
rect 13490 6854 13532 6906
rect 13550 6854 13596 6906
rect 13596 6854 13602 6906
rect 13200 6790 13252 6842
rect 13270 6790 13322 6842
rect 13340 6790 13392 6842
rect 13410 6790 13462 6842
rect 13480 6790 13490 6842
rect 13490 6790 13532 6842
rect 13550 6790 13596 6842
rect 13596 6790 13602 6842
rect 13200 6726 13252 6778
rect 13270 6726 13322 6778
rect 13340 6726 13392 6778
rect 13410 6726 13462 6778
rect 13480 6726 13490 6778
rect 13490 6726 13532 6778
rect 13550 6726 13596 6778
rect 13596 6726 13602 6778
rect 13200 6680 13205 6714
rect 13205 6680 13239 6714
rect 13239 6680 13252 6714
rect 13200 6662 13252 6680
rect 13270 6680 13277 6714
rect 13277 6680 13311 6714
rect 13311 6680 13322 6714
rect 13270 6662 13322 6680
rect 13340 6662 13392 6714
rect 13410 6662 13462 6714
rect 13480 6662 13490 6714
rect 13490 6662 13532 6714
rect 13550 6662 13596 6714
rect 13596 6662 13602 6714
rect 13200 6641 13252 6650
rect 13200 6607 13205 6641
rect 13205 6607 13239 6641
rect 13239 6607 13252 6641
rect 13200 6598 13252 6607
rect 13270 6641 13322 6650
rect 13270 6607 13277 6641
rect 13277 6607 13311 6641
rect 13311 6607 13322 6641
rect 13270 6598 13322 6607
rect 13340 6598 13392 6650
rect 13410 6598 13462 6650
rect 13480 6598 13490 6650
rect 13490 6598 13532 6650
rect 13550 6598 13596 6650
rect 13596 6598 13602 6650
rect 13200 6568 13252 6586
rect 13200 6534 13205 6568
rect 13205 6534 13239 6568
rect 13239 6534 13252 6568
rect 13270 6568 13322 6586
rect 13270 6534 13277 6568
rect 13277 6534 13311 6568
rect 13311 6534 13322 6568
rect 13340 6534 13392 6586
rect 13410 6534 13462 6586
rect 13480 6534 13490 6586
rect 13490 6534 13532 6586
rect 13550 6534 13596 6586
rect 13596 6534 13602 6586
rect 13200 6495 13252 6522
rect 13200 6470 13205 6495
rect 13205 6470 13239 6495
rect 13239 6470 13252 6495
rect 13270 6495 13322 6522
rect 13270 6470 13277 6495
rect 13277 6470 13311 6495
rect 13311 6470 13322 6495
rect 13340 6470 13392 6522
rect 13410 6470 13462 6522
rect 13480 6470 13490 6522
rect 13490 6470 13532 6522
rect 13550 6470 13596 6522
rect 13596 6470 13602 6522
rect 13200 6422 13252 6458
rect 13270 6422 13322 6458
rect 13200 6406 13205 6422
rect 13205 6406 13252 6422
rect 13270 6406 13311 6422
rect 13311 6406 13322 6422
rect 13340 6406 13392 6458
rect 13410 6406 13462 6458
rect 13480 6406 13490 6458
rect 13490 6406 13532 6458
rect 13550 6406 13596 6458
rect 13596 6406 13602 6458
rect 13200 6342 13205 6394
rect 13205 6342 13252 6394
rect 13270 6342 13311 6394
rect 13311 6342 13322 6394
rect 13340 6342 13392 6394
rect 13410 6342 13462 6394
rect 13480 6342 13490 6394
rect 13490 6342 13532 6394
rect 13550 6342 13596 6394
rect 13596 6342 13602 6394
rect 13200 6278 13205 6330
rect 13205 6278 13252 6330
rect 13270 6278 13311 6330
rect 13311 6278 13322 6330
rect 13340 6278 13392 6330
rect 13410 6278 13462 6330
rect 13480 6278 13490 6330
rect 13490 6278 13532 6330
rect 13550 6278 13596 6330
rect 13596 6278 13602 6330
rect 13200 6214 13205 6266
rect 13205 6214 13252 6266
rect 13270 6214 13311 6266
rect 13311 6214 13322 6266
rect 13340 6214 13392 6266
rect 13410 6214 13462 6266
rect 13480 6214 13490 6266
rect 13490 6214 13532 6266
rect 13550 6214 13596 6266
rect 13596 6214 13602 6266
rect 13200 6150 13205 6202
rect 13205 6150 13252 6202
rect 13270 6150 13311 6202
rect 13311 6150 13322 6202
rect 13340 6150 13392 6202
rect 13410 6150 13462 6202
rect 13480 6150 13490 6202
rect 13490 6150 13532 6202
rect 13550 6150 13596 6202
rect 13596 6150 13602 6202
rect 13200 6086 13205 6138
rect 13205 6086 13252 6138
rect 13270 6086 13311 6138
rect 13311 6086 13322 6138
rect 13340 6086 13392 6138
rect 13410 6086 13462 6138
rect 13480 6086 13490 6138
rect 13490 6086 13532 6138
rect 13550 6086 13596 6138
rect 13596 6086 13602 6138
rect 13200 6022 13205 6074
rect 13205 6022 13252 6074
rect 13270 6022 13311 6074
rect 13311 6022 13322 6074
rect 13340 6022 13392 6074
rect 13410 6022 13462 6074
rect 13480 6022 13490 6074
rect 13490 6022 13532 6074
rect 13550 6022 13596 6074
rect 13596 6022 13602 6074
rect 13200 5958 13205 6010
rect 13205 5958 13252 6010
rect 13270 5958 13311 6010
rect 13311 5958 13322 6010
rect 13340 5958 13392 6010
rect 13410 5958 13462 6010
rect 13480 5958 13490 6010
rect 13490 5958 13532 6010
rect 13550 5958 13596 6010
rect 13596 5958 13602 6010
rect 13200 5894 13205 5946
rect 13205 5894 13252 5946
rect 13270 5894 13311 5946
rect 13311 5894 13322 5946
rect 13340 5894 13392 5946
rect 13410 5894 13462 5946
rect 13480 5894 13490 5946
rect 13490 5894 13532 5946
rect 13550 5894 13596 5946
rect 13596 5894 13602 5946
rect 13200 5830 13205 5882
rect 13205 5830 13252 5882
rect 13270 5830 13311 5882
rect 13311 5830 13322 5882
rect 13340 5830 13392 5882
rect 13410 5830 13462 5882
rect 13480 5830 13490 5882
rect 13490 5830 13532 5882
rect 13550 5830 13596 5882
rect 13596 5830 13602 5882
rect 13200 5766 13205 5818
rect 13205 5766 13252 5818
rect 13270 5766 13311 5818
rect 13311 5766 13322 5818
rect 13340 5766 13392 5818
rect 13410 5766 13462 5818
rect 13480 5815 13490 5818
rect 13490 5815 13532 5818
rect 13550 5815 13596 5818
rect 13596 5815 13602 5818
rect 13480 5776 13532 5815
rect 13480 5766 13490 5776
rect 13490 5766 13524 5776
rect 13524 5766 13532 5776
rect 13550 5776 13602 5815
rect 13550 5766 13562 5776
rect 13562 5766 13596 5776
rect 13596 5766 13602 5776
rect 13200 5702 13205 5754
rect 13205 5702 13252 5754
rect 13270 5702 13311 5754
rect 13311 5702 13322 5754
rect 13340 5702 13392 5754
rect 13410 5702 13462 5754
rect 13480 5742 13490 5754
rect 13490 5742 13524 5754
rect 13524 5742 13532 5754
rect 13480 5703 13532 5742
rect 13480 5702 13490 5703
rect 13490 5702 13524 5703
rect 13524 5702 13532 5703
rect 13550 5742 13562 5754
rect 13562 5742 13596 5754
rect 13596 5742 13602 5754
rect 13550 5703 13602 5742
rect 13550 5702 13562 5703
rect 13562 5702 13596 5703
rect 13596 5702 13602 5703
rect 13200 5638 13205 5690
rect 13205 5638 13252 5690
rect 13270 5638 13311 5690
rect 13311 5638 13322 5690
rect 13340 5638 13392 5690
rect 13410 5638 13462 5690
rect 13480 5669 13490 5690
rect 13490 5669 13524 5690
rect 13524 5669 13532 5690
rect 13480 5638 13532 5669
rect 13550 5669 13562 5690
rect 13562 5669 13596 5690
rect 13596 5669 13602 5690
rect 13550 5638 13602 5669
rect 13200 5574 13205 5626
rect 13205 5574 13252 5626
rect 13270 5574 13311 5626
rect 13311 5574 13322 5626
rect 13340 5574 13392 5626
rect 13410 5574 13462 5626
rect 13480 5596 13490 5626
rect 13490 5596 13524 5626
rect 13524 5596 13532 5626
rect 13480 5574 13532 5596
rect 13550 5596 13562 5626
rect 13562 5596 13596 5626
rect 13596 5596 13602 5626
rect 13550 5574 13602 5596
rect 13200 5510 13205 5562
rect 13205 5510 13252 5562
rect 13270 5510 13311 5562
rect 13311 5510 13322 5562
rect 13340 5510 13392 5562
rect 13410 5510 13462 5562
rect 13480 5557 13532 5562
rect 13480 5523 13490 5557
rect 13490 5523 13524 5557
rect 13524 5523 13532 5557
rect 13480 5510 13532 5523
rect 13550 5557 13602 5562
rect 13550 5523 13562 5557
rect 13562 5523 13596 5557
rect 13596 5523 13602 5557
rect 13550 5510 13602 5523
rect 13200 5446 13205 5498
rect 13205 5446 13252 5498
rect 13270 5446 13311 5498
rect 13311 5446 13322 5498
rect 13340 5446 13392 5498
rect 13410 5446 13462 5498
rect 13480 5484 13532 5498
rect 13480 5450 13490 5484
rect 13490 5450 13524 5484
rect 13524 5450 13532 5484
rect 13480 5446 13532 5450
rect 13550 5484 13602 5498
rect 13550 5450 13562 5484
rect 13562 5450 13596 5484
rect 13596 5450 13602 5484
rect 13550 5446 13602 5450
rect 13200 5382 13205 5434
rect 13205 5382 13252 5434
rect 13270 5382 13311 5434
rect 13311 5382 13322 5434
rect 13340 5382 13392 5434
rect 13410 5382 13462 5434
rect 13480 5411 13532 5434
rect 13480 5382 13490 5411
rect 13490 5382 13524 5411
rect 13524 5382 13532 5411
rect 13550 5411 13602 5434
rect 13550 5382 13562 5411
rect 13562 5382 13596 5411
rect 13596 5382 13602 5411
rect 12922 5378 12974 5380
rect 12988 5378 13040 5380
rect 13200 5318 13252 5370
rect 13270 5318 13322 5370
rect 13340 5318 13392 5370
rect 13410 5318 13462 5370
rect 13480 5338 13532 5370
rect 13480 5318 13490 5338
rect 13490 5318 13524 5338
rect 13524 5318 13532 5338
rect 13550 5338 13602 5370
rect 13550 5318 13562 5338
rect 13562 5318 13596 5338
rect 13596 5318 13602 5338
rect 13200 5254 13252 5306
rect 13270 5254 13322 5306
rect 13340 5254 13392 5306
rect 13410 5254 13462 5306
rect 13480 5304 13490 5306
rect 13490 5304 13524 5306
rect 13524 5304 13532 5306
rect 13480 5265 13532 5304
rect 13480 5254 13490 5265
rect 13490 5254 13524 5265
rect 13524 5254 13532 5265
rect 13550 5304 13562 5306
rect 13562 5304 13596 5306
rect 13596 5304 13602 5306
rect 13550 5265 13602 5304
rect 13550 5254 13562 5265
rect 13562 5254 13596 5265
rect 13596 5254 13602 5265
rect 13200 5197 13252 5242
rect 13270 5197 13322 5242
rect 13340 5197 13392 5242
rect 13410 5197 13462 5242
rect 13200 5190 13252 5197
rect 13270 5190 13322 5197
rect 13340 5190 13392 5197
rect 13410 5190 13452 5197
rect 13452 5190 13462 5197
rect 13480 5231 13490 5242
rect 13490 5231 13524 5242
rect 13524 5231 13532 5242
rect 13480 5192 13532 5231
rect 13480 5190 13490 5192
rect 13490 5190 13524 5192
rect 13524 5190 13532 5192
rect 13550 5231 13562 5242
rect 13562 5231 13596 5242
rect 13596 5231 13602 5242
rect 13550 5192 13602 5231
rect 13550 5190 13562 5192
rect 13562 5190 13596 5192
rect 13596 5190 13602 5192
rect 13200 5126 13252 5178
rect 13270 5126 13322 5178
rect 13340 5126 13392 5178
rect 13410 5126 13452 5178
rect 13452 5126 13462 5178
rect 13480 5158 13490 5178
rect 13490 5158 13524 5178
rect 13524 5158 13532 5178
rect 13480 5126 13532 5158
rect 13550 5158 13562 5178
rect 13562 5158 13596 5178
rect 13596 5158 13602 5178
rect 13550 5126 13602 5158
rect 13200 5062 13252 5114
rect 13270 5062 13322 5114
rect 13340 5062 13392 5114
rect 13410 5062 13452 5114
rect 13452 5062 13462 5114
rect 13480 5085 13490 5114
rect 13490 5085 13524 5114
rect 13524 5085 13532 5114
rect 13480 5062 13532 5085
rect 13550 5085 13562 5114
rect 13562 5085 13596 5114
rect 13596 5085 13602 5114
rect 13550 5062 13602 5085
rect 13200 5019 13252 5049
rect 13270 5019 13322 5049
rect 13340 5019 13392 5049
rect 13410 5019 13452 5049
rect 13452 5019 13462 5049
rect 13200 4997 13252 5019
rect 13270 4997 13322 5019
rect 13340 4997 13392 5019
rect 13410 4997 13462 5019
rect 13480 4997 13532 5049
rect 13550 4997 13602 5049
rect 4968 4871 5020 4877
rect 5085 4871 5137 4877
rect 5202 4871 5254 4877
rect 4968 4837 4977 4871
rect 4977 4837 5016 4871
rect 5016 4837 5020 4871
rect 5085 4837 5089 4871
rect 5089 4837 5123 4871
rect 5123 4837 5137 4871
rect 4968 4825 5020 4837
rect 5085 4825 5137 4837
rect 5202 4825 5235 4871
rect 5235 4825 5254 4871
rect 4968 4799 5020 4811
rect 5085 4799 5137 4811
rect 4968 4765 4977 4799
rect 4977 4765 5016 4799
rect 5016 4765 5020 4799
rect 5085 4765 5089 4799
rect 5089 4765 5123 4799
rect 5123 4765 5137 4799
rect 5202 4765 5235 4811
rect 5235 4765 5254 4811
rect 4968 4759 5020 4765
rect 5085 4759 5137 4765
rect 5202 4759 5254 4765
rect 10369 4669 10421 4721
rect 10445 4669 10497 4721
rect 10369 4583 10421 4635
rect 10445 4583 10497 4635
rect 5209 4168 5261 4220
rect 5278 4168 5330 4220
rect 5346 4168 5398 4220
rect 5414 4168 5466 4220
rect 5482 4168 5534 4220
rect 5550 4168 5602 4220
rect 5618 4168 5670 4220
rect 5686 4168 5738 4220
rect 5754 4168 5806 4220
rect 5822 4168 5874 4220
rect 5890 4168 5942 4220
rect 5209 4044 5261 4096
rect 5278 4044 5330 4096
rect 5346 4044 5398 4096
rect 5414 4044 5466 4096
rect 5482 4044 5534 4096
rect 5550 4044 5602 4096
rect 5618 4044 5670 4096
rect 5686 4044 5738 4096
rect 5754 4044 5806 4096
rect 5822 4044 5874 4096
rect 5890 4044 5942 4096
rect 4820 3664 4872 3666
rect 4885 3664 4937 3666
rect 4820 3630 4840 3664
rect 4840 3630 4872 3664
rect 4885 3630 4912 3664
rect 4912 3630 4937 3664
rect 4820 3614 4872 3630
rect 4885 3614 4937 3630
rect 4950 3664 5002 3666
rect 4950 3630 4984 3664
rect 4984 3630 5002 3664
rect 4950 3614 5002 3630
rect 5015 3664 5067 3666
rect 5015 3630 5022 3664
rect 5022 3630 5056 3664
rect 5056 3630 5067 3664
rect 5015 3614 5067 3630
rect 5080 3664 5132 3666
rect 5080 3630 5094 3664
rect 5094 3630 5128 3664
rect 5128 3630 5132 3664
rect 5080 3614 5132 3630
rect 5145 3664 5197 3666
rect 5210 3664 5262 3666
rect 5275 3664 5327 3666
rect 5340 3664 5392 3666
rect 5405 3664 5457 3666
rect 5470 3664 5522 3666
rect 5535 3664 5587 3666
rect 5600 3664 5652 3666
rect 5145 3630 5166 3664
rect 5166 3630 5197 3664
rect 5210 3630 5238 3664
rect 5238 3630 5262 3664
rect 5275 3630 5310 3664
rect 5310 3630 5327 3664
rect 5340 3630 5344 3664
rect 5344 3630 5382 3664
rect 5382 3630 5392 3664
rect 5405 3630 5416 3664
rect 5416 3630 5454 3664
rect 5454 3630 5457 3664
rect 5470 3630 5488 3664
rect 5488 3630 5522 3664
rect 5535 3630 5560 3664
rect 5560 3630 5587 3664
rect 5600 3630 5632 3664
rect 5632 3630 5652 3664
rect 5145 3614 5197 3630
rect 5210 3614 5262 3630
rect 5275 3614 5327 3630
rect 5340 3614 5392 3630
rect 5405 3614 5457 3630
rect 5470 3614 5522 3630
rect 5535 3614 5587 3630
rect 5600 3614 5652 3630
rect 5665 3664 5717 3666
rect 5665 3630 5670 3664
rect 5670 3630 5704 3664
rect 5704 3630 5717 3664
rect 5665 3614 5717 3630
rect 5730 3664 5782 3666
rect 5730 3630 5742 3664
rect 5742 3630 5776 3664
rect 5776 3630 5782 3664
rect 5730 3614 5782 3630
rect 5795 3664 5847 3666
rect 5860 3664 5912 3666
rect 5925 3664 5977 3666
rect 5990 3664 6042 3666
rect 6055 3664 6107 3666
rect 6120 3664 6172 3666
rect 6185 3664 6237 3666
rect 6250 3664 6302 3666
rect 5795 3630 5814 3664
rect 5814 3630 5847 3664
rect 5860 3630 5886 3664
rect 5886 3630 5912 3664
rect 5925 3630 5958 3664
rect 5958 3630 5977 3664
rect 5990 3630 5992 3664
rect 5992 3630 6030 3664
rect 6030 3630 6042 3664
rect 6055 3630 6064 3664
rect 6064 3630 6102 3664
rect 6102 3630 6107 3664
rect 6120 3630 6136 3664
rect 6136 3630 6172 3664
rect 6185 3630 6208 3664
rect 6208 3630 6237 3664
rect 6250 3630 6280 3664
rect 6280 3630 6302 3664
rect 5795 3614 5847 3630
rect 5860 3614 5912 3630
rect 5925 3614 5977 3630
rect 5990 3614 6042 3630
rect 6055 3614 6107 3630
rect 6120 3614 6172 3630
rect 6185 3614 6237 3630
rect 6250 3614 6302 3630
rect 6315 3664 6367 3666
rect 6315 3630 6318 3664
rect 6318 3630 6352 3664
rect 6352 3630 6367 3664
rect 6315 3614 6367 3630
rect 6380 3664 6432 3666
rect 6380 3630 6390 3664
rect 6390 3630 6424 3664
rect 6424 3630 6432 3664
rect 6380 3614 6432 3630
rect 6445 3664 6497 3666
rect 6445 3630 6462 3664
rect 6462 3630 6496 3664
rect 6496 3630 6497 3664
rect 6445 3614 6497 3630
rect 6510 3664 6562 3666
rect 6575 3664 6627 3666
rect 6640 3664 6692 3666
rect 6705 3664 6757 3666
rect 6770 3664 6822 3666
rect 6835 3664 6887 3666
rect 6900 3664 6952 3666
rect 6510 3630 6534 3664
rect 6534 3630 6562 3664
rect 6575 3630 6606 3664
rect 6606 3630 6627 3664
rect 6640 3630 6678 3664
rect 6678 3630 6692 3664
rect 6705 3630 6712 3664
rect 6712 3630 6750 3664
rect 6750 3630 6757 3664
rect 6770 3630 6784 3664
rect 6784 3630 6822 3664
rect 6835 3630 6856 3664
rect 6856 3630 6887 3664
rect 6900 3630 6928 3664
rect 6928 3630 6952 3664
rect 6510 3614 6562 3630
rect 6575 3614 6627 3630
rect 6640 3614 6692 3630
rect 6705 3614 6757 3630
rect 6770 3614 6822 3630
rect 6835 3614 6887 3630
rect 6900 3614 6952 3630
rect 6965 3664 7017 3666
rect 6965 3630 6966 3664
rect 6966 3630 7000 3664
rect 7000 3630 7017 3664
rect 6965 3614 7017 3630
rect 7030 3664 7082 3666
rect 7030 3630 7038 3664
rect 7038 3630 7072 3664
rect 7072 3630 7082 3664
rect 7030 3614 7082 3630
rect 7095 3664 7147 3666
rect 7095 3630 7110 3664
rect 7110 3630 7144 3664
rect 7144 3630 7147 3664
rect 7095 3614 7147 3630
rect 7160 3664 7212 3666
rect 7160 3630 7182 3664
rect 7182 3630 7212 3664
rect 7160 3614 7212 3630
rect 7225 3614 7277 3666
rect 7290 3614 7342 3666
rect 7355 3614 7407 3666
rect 7419 3664 7471 3666
rect 7419 3630 7428 3664
rect 7428 3630 7462 3664
rect 7462 3630 7471 3664
rect 7419 3614 7471 3630
rect 7483 3664 7535 3666
rect 7483 3630 7501 3664
rect 7501 3630 7535 3664
rect 7483 3614 7535 3630
rect 7547 3664 7599 3666
rect 7611 3664 7663 3666
rect 7675 3664 7727 3666
rect 7739 3664 7791 3666
rect 7803 3664 7855 3666
rect 7867 3664 7919 3666
rect 7547 3630 7574 3664
rect 7574 3630 7599 3664
rect 7611 3630 7646 3664
rect 7646 3630 7663 3664
rect 7675 3630 7680 3664
rect 7680 3630 7718 3664
rect 7718 3630 7727 3664
rect 7739 3630 7752 3664
rect 7752 3630 7790 3664
rect 7790 3630 7791 3664
rect 7803 3630 7824 3664
rect 7824 3630 7855 3664
rect 7867 3630 7896 3664
rect 7896 3630 7919 3664
rect 7547 3614 7599 3630
rect 7611 3614 7663 3630
rect 7675 3614 7727 3630
rect 7739 3614 7791 3630
rect 7803 3614 7855 3630
rect 7867 3614 7919 3630
rect 7931 3664 7983 3666
rect 7931 3630 7934 3664
rect 7934 3630 7968 3664
rect 7968 3630 7983 3664
rect 7931 3614 7983 3630
rect 7995 3664 8047 3666
rect 7995 3630 8006 3664
rect 8006 3630 8040 3664
rect 8040 3630 8047 3664
rect 7995 3614 8047 3630
rect 8059 3664 8111 3666
rect 8123 3664 8175 3666
rect 8187 3664 8239 3666
rect 8251 3664 8303 3666
rect 8315 3664 8367 3666
rect 8379 3664 8431 3666
rect 8443 3664 8495 3666
rect 8059 3630 8078 3664
rect 8078 3630 8111 3664
rect 8123 3630 8150 3664
rect 8150 3630 8175 3664
rect 8187 3630 8222 3664
rect 8222 3630 8239 3664
rect 8251 3630 8256 3664
rect 8256 3630 8294 3664
rect 8294 3630 8303 3664
rect 8315 3630 8328 3664
rect 8328 3630 8366 3664
rect 8366 3630 8367 3664
rect 8379 3630 8400 3664
rect 8400 3630 8431 3664
rect 8443 3630 8472 3664
rect 8472 3630 8495 3664
rect 8059 3614 8111 3630
rect 8123 3614 8175 3630
rect 8187 3614 8239 3630
rect 8251 3614 8303 3630
rect 8315 3614 8367 3630
rect 8379 3614 8431 3630
rect 8443 3614 8495 3630
rect 8507 3664 8559 3666
rect 8507 3630 8510 3664
rect 8510 3630 8544 3664
rect 8544 3630 8559 3664
rect 8507 3614 8559 3630
rect 8571 3664 8623 3666
rect 8571 3630 8582 3664
rect 8582 3630 8616 3664
rect 8616 3630 8623 3664
rect 8571 3614 8623 3630
rect 8635 3664 8687 3666
rect 8699 3664 8751 3666
rect 8763 3664 8815 3666
rect 8827 3664 8879 3666
rect 8891 3664 8943 3666
rect 8955 3664 9007 3666
rect 9019 3664 9071 3666
rect 8635 3630 8654 3664
rect 8654 3630 8687 3664
rect 8699 3630 8726 3664
rect 8726 3630 8751 3664
rect 8763 3630 8798 3664
rect 8798 3630 8815 3664
rect 8827 3630 8832 3664
rect 8832 3630 8870 3664
rect 8870 3630 8879 3664
rect 8891 3630 8904 3664
rect 8904 3630 8942 3664
rect 8942 3630 8943 3664
rect 8955 3630 8976 3664
rect 8976 3630 9007 3664
rect 9019 3630 9048 3664
rect 9048 3630 9071 3664
rect 8635 3614 8687 3630
rect 8699 3614 8751 3630
rect 8763 3614 8815 3630
rect 8827 3614 8879 3630
rect 8891 3614 8943 3630
rect 8955 3614 9007 3630
rect 9019 3614 9071 3630
rect 9083 3664 9135 3666
rect 9083 3630 9086 3664
rect 9086 3630 9120 3664
rect 9120 3630 9135 3664
rect 9083 3614 9135 3630
rect 9147 3664 9199 3666
rect 9147 3630 9158 3664
rect 9158 3630 9192 3664
rect 9192 3630 9199 3664
rect 9147 3614 9199 3630
rect 9211 3664 9263 3666
rect 9275 3664 9327 3666
rect 9339 3664 9391 3666
rect 9403 3664 9455 3666
rect 9467 3664 9519 3666
rect 9531 3664 9583 3666
rect 9595 3664 9647 3666
rect 9211 3630 9230 3664
rect 9230 3630 9263 3664
rect 9275 3630 9302 3664
rect 9302 3630 9327 3664
rect 9339 3630 9374 3664
rect 9374 3630 9391 3664
rect 9403 3630 9408 3664
rect 9408 3630 9446 3664
rect 9446 3630 9455 3664
rect 9467 3630 9480 3664
rect 9480 3630 9518 3664
rect 9518 3630 9519 3664
rect 9531 3630 9552 3664
rect 9552 3630 9583 3664
rect 9595 3630 9624 3664
rect 9624 3630 9647 3664
rect 9211 3614 9263 3630
rect 9275 3614 9327 3630
rect 9339 3614 9391 3630
rect 9403 3614 9455 3630
rect 9467 3614 9519 3630
rect 9531 3614 9583 3630
rect 9595 3614 9647 3630
rect 9659 3664 9711 3666
rect 9659 3630 9662 3664
rect 9662 3630 9696 3664
rect 9696 3630 9711 3664
rect 9659 3614 9711 3630
rect 9723 3664 9775 3666
rect 9723 3630 9734 3664
rect 9734 3630 9768 3664
rect 9768 3630 9775 3664
rect 9723 3614 9775 3630
rect 9787 3664 9839 3666
rect 9851 3664 9903 3666
rect 9915 3664 9967 3666
rect 9979 3664 10031 3666
rect 10043 3664 10095 3666
rect 10107 3664 10159 3666
rect 10171 3664 10223 3666
rect 9787 3630 9806 3664
rect 9806 3630 9839 3664
rect 9851 3630 9878 3664
rect 9878 3630 9903 3664
rect 9915 3630 9950 3664
rect 9950 3630 9967 3664
rect 9979 3630 9984 3664
rect 9984 3630 10022 3664
rect 10022 3630 10031 3664
rect 10043 3630 10056 3664
rect 10056 3630 10094 3664
rect 10094 3630 10095 3664
rect 10107 3630 10128 3664
rect 10128 3630 10159 3664
rect 10171 3630 10200 3664
rect 10200 3630 10223 3664
rect 9787 3614 9839 3630
rect 9851 3614 9903 3630
rect 9915 3614 9967 3630
rect 9979 3614 10031 3630
rect 10043 3614 10095 3630
rect 10107 3614 10159 3630
rect 10171 3614 10223 3630
rect 10235 3664 10287 3666
rect 10235 3630 10238 3664
rect 10238 3630 10272 3664
rect 10272 3630 10287 3664
rect 10235 3614 10287 3630
rect 10299 3664 10351 3666
rect 10299 3630 10310 3664
rect 10310 3630 10344 3664
rect 10344 3630 10351 3664
rect 10299 3614 10351 3630
rect 10363 3664 10415 3666
rect 10427 3664 10479 3666
rect 10491 3664 10543 3666
rect 10555 3664 10607 3666
rect 10619 3664 10671 3666
rect 10683 3664 10735 3666
rect 10747 3664 10799 3666
rect 10363 3630 10382 3664
rect 10382 3630 10415 3664
rect 10427 3630 10454 3664
rect 10454 3630 10479 3664
rect 10491 3630 10526 3664
rect 10526 3630 10543 3664
rect 10555 3630 10560 3664
rect 10560 3630 10598 3664
rect 10598 3630 10607 3664
rect 10619 3630 10632 3664
rect 10632 3630 10670 3664
rect 10670 3630 10671 3664
rect 10683 3630 10704 3664
rect 10704 3630 10735 3664
rect 10747 3630 10776 3664
rect 10776 3630 10799 3664
rect 10363 3614 10415 3630
rect 10427 3614 10479 3630
rect 10491 3614 10543 3630
rect 10555 3614 10607 3630
rect 10619 3614 10671 3630
rect 10683 3614 10735 3630
rect 10747 3614 10799 3630
rect 10811 3664 10863 3666
rect 10811 3630 10814 3664
rect 10814 3630 10848 3664
rect 10848 3630 10863 3664
rect 10811 3614 10863 3630
rect 4820 3556 4872 3578
rect 4885 3556 4937 3578
rect 4820 3526 4840 3556
rect 4840 3526 4872 3556
rect 4885 3526 4912 3556
rect 4912 3526 4937 3556
rect 4950 3556 5002 3578
rect 4950 3526 4984 3556
rect 4984 3526 5002 3556
rect 5015 3556 5067 3578
rect 5015 3526 5022 3556
rect 5022 3526 5056 3556
rect 5056 3526 5067 3556
rect 5080 3556 5132 3578
rect 5080 3526 5094 3556
rect 5094 3526 5128 3556
rect 5128 3526 5132 3556
rect 5145 3556 5197 3578
rect 5210 3556 5262 3578
rect 5275 3556 5327 3578
rect 5340 3556 5392 3578
rect 5405 3556 5457 3578
rect 5470 3556 5522 3578
rect 5535 3556 5587 3578
rect 5600 3556 5652 3578
rect 5145 3526 5166 3556
rect 5166 3526 5197 3556
rect 5210 3526 5238 3556
rect 5238 3526 5262 3556
rect 5275 3526 5310 3556
rect 5310 3526 5327 3556
rect 5340 3526 5344 3556
rect 5344 3526 5382 3556
rect 5382 3526 5392 3556
rect 5405 3526 5416 3556
rect 5416 3526 5454 3556
rect 5454 3526 5457 3556
rect 5470 3526 5488 3556
rect 5488 3526 5522 3556
rect 5535 3526 5560 3556
rect 5560 3526 5587 3556
rect 5600 3526 5632 3556
rect 5632 3526 5652 3556
rect 5665 3556 5717 3578
rect 5665 3526 5670 3556
rect 5670 3526 5704 3556
rect 5704 3526 5717 3556
rect 5730 3556 5782 3578
rect 5730 3526 5742 3556
rect 5742 3526 5776 3556
rect 5776 3526 5782 3556
rect 5795 3556 5847 3578
rect 5860 3556 5912 3578
rect 5925 3556 5977 3578
rect 5990 3556 6042 3578
rect 6055 3556 6107 3578
rect 6120 3556 6172 3578
rect 6185 3556 6237 3578
rect 6250 3556 6302 3578
rect 5795 3526 5814 3556
rect 5814 3526 5847 3556
rect 5860 3526 5886 3556
rect 5886 3526 5912 3556
rect 5925 3526 5958 3556
rect 5958 3526 5977 3556
rect 5990 3526 5992 3556
rect 5992 3526 6030 3556
rect 6030 3526 6042 3556
rect 6055 3526 6064 3556
rect 6064 3526 6102 3556
rect 6102 3526 6107 3556
rect 6120 3526 6136 3556
rect 6136 3526 6172 3556
rect 6185 3526 6208 3556
rect 6208 3526 6237 3556
rect 6250 3526 6280 3556
rect 6280 3526 6302 3556
rect 6315 3556 6367 3578
rect 6315 3526 6318 3556
rect 6318 3526 6352 3556
rect 6352 3526 6367 3556
rect 6380 3556 6432 3578
rect 6380 3526 6390 3556
rect 6390 3526 6424 3556
rect 6424 3526 6432 3556
rect 6445 3556 6497 3578
rect 6445 3526 6462 3556
rect 6462 3526 6496 3556
rect 6496 3526 6497 3556
rect 6510 3556 6562 3578
rect 6575 3556 6627 3578
rect 6640 3556 6692 3578
rect 6705 3556 6757 3578
rect 6770 3556 6822 3578
rect 6835 3556 6887 3578
rect 6900 3556 6952 3578
rect 6510 3526 6534 3556
rect 6534 3526 6562 3556
rect 6575 3526 6606 3556
rect 6606 3526 6627 3556
rect 6640 3526 6678 3556
rect 6678 3526 6692 3556
rect 6705 3526 6712 3556
rect 6712 3526 6750 3556
rect 6750 3526 6757 3556
rect 6770 3526 6784 3556
rect 6784 3526 6822 3556
rect 6835 3526 6856 3556
rect 6856 3526 6887 3556
rect 6900 3526 6928 3556
rect 6928 3526 6952 3556
rect 6965 3556 7017 3578
rect 6965 3526 6966 3556
rect 6966 3526 7000 3556
rect 7000 3526 7017 3556
rect 7030 3556 7082 3578
rect 7030 3526 7038 3556
rect 7038 3526 7072 3556
rect 7072 3526 7082 3556
rect 7095 3556 7147 3578
rect 7095 3526 7110 3556
rect 7110 3526 7144 3556
rect 7144 3526 7147 3556
rect 7160 3556 7212 3578
rect 7160 3526 7182 3556
rect 7182 3526 7212 3556
rect 7225 3526 7277 3578
rect 7290 3526 7342 3578
rect 7355 3526 7407 3578
rect 7419 3556 7471 3578
rect 7419 3526 7428 3556
rect 7428 3526 7462 3556
rect 7462 3526 7471 3556
rect 7483 3556 7535 3578
rect 7483 3526 7501 3556
rect 7501 3526 7535 3556
rect 7547 3556 7599 3578
rect 7611 3556 7663 3578
rect 7675 3556 7727 3578
rect 7739 3556 7791 3578
rect 7803 3556 7855 3578
rect 7867 3556 7919 3578
rect 7547 3526 7574 3556
rect 7574 3526 7599 3556
rect 7611 3526 7646 3556
rect 7646 3526 7663 3556
rect 7675 3526 7680 3556
rect 7680 3526 7718 3556
rect 7718 3526 7727 3556
rect 7739 3526 7752 3556
rect 7752 3526 7790 3556
rect 7790 3526 7791 3556
rect 7803 3526 7824 3556
rect 7824 3526 7855 3556
rect 7867 3526 7896 3556
rect 7896 3526 7919 3556
rect 7931 3556 7983 3578
rect 7931 3526 7934 3556
rect 7934 3526 7968 3556
rect 7968 3526 7983 3556
rect 7995 3556 8047 3578
rect 7995 3526 8006 3556
rect 8006 3526 8040 3556
rect 8040 3526 8047 3556
rect 8059 3556 8111 3578
rect 8123 3556 8175 3578
rect 8187 3556 8239 3578
rect 8251 3556 8303 3578
rect 8315 3556 8367 3578
rect 8379 3556 8431 3578
rect 8443 3556 8495 3578
rect 8059 3526 8078 3556
rect 8078 3526 8111 3556
rect 8123 3526 8150 3556
rect 8150 3526 8175 3556
rect 8187 3526 8222 3556
rect 8222 3526 8239 3556
rect 8251 3526 8256 3556
rect 8256 3526 8294 3556
rect 8294 3526 8303 3556
rect 8315 3526 8328 3556
rect 8328 3526 8366 3556
rect 8366 3526 8367 3556
rect 8379 3526 8400 3556
rect 8400 3526 8431 3556
rect 8443 3526 8472 3556
rect 8472 3526 8495 3556
rect 8507 3556 8559 3578
rect 8507 3526 8510 3556
rect 8510 3526 8544 3556
rect 8544 3526 8559 3556
rect 8571 3556 8623 3578
rect 8571 3526 8582 3556
rect 8582 3526 8616 3556
rect 8616 3526 8623 3556
rect 8635 3556 8687 3578
rect 8699 3556 8751 3578
rect 8763 3556 8815 3578
rect 8827 3556 8879 3578
rect 8891 3556 8943 3578
rect 8955 3556 9007 3578
rect 9019 3556 9071 3578
rect 8635 3526 8654 3556
rect 8654 3526 8687 3556
rect 8699 3526 8726 3556
rect 8726 3526 8751 3556
rect 8763 3526 8798 3556
rect 8798 3526 8815 3556
rect 8827 3526 8832 3556
rect 8832 3526 8870 3556
rect 8870 3526 8879 3556
rect 8891 3526 8904 3556
rect 8904 3526 8942 3556
rect 8942 3526 8943 3556
rect 8955 3526 8976 3556
rect 8976 3526 9007 3556
rect 9019 3526 9048 3556
rect 9048 3526 9071 3556
rect 9083 3556 9135 3578
rect 9083 3526 9086 3556
rect 9086 3526 9120 3556
rect 9120 3526 9135 3556
rect 9147 3556 9199 3578
rect 9147 3526 9158 3556
rect 9158 3526 9192 3556
rect 9192 3526 9199 3556
rect 9211 3556 9263 3578
rect 9275 3556 9327 3578
rect 9339 3556 9391 3578
rect 9403 3556 9455 3578
rect 9467 3556 9519 3578
rect 9531 3556 9583 3578
rect 9595 3556 9647 3578
rect 9211 3526 9230 3556
rect 9230 3526 9263 3556
rect 9275 3526 9302 3556
rect 9302 3526 9327 3556
rect 9339 3526 9374 3556
rect 9374 3526 9391 3556
rect 9403 3526 9408 3556
rect 9408 3526 9446 3556
rect 9446 3526 9455 3556
rect 9467 3526 9480 3556
rect 9480 3526 9518 3556
rect 9518 3526 9519 3556
rect 9531 3526 9552 3556
rect 9552 3526 9583 3556
rect 9595 3526 9624 3556
rect 9624 3526 9647 3556
rect 9659 3556 9711 3578
rect 9659 3526 9662 3556
rect 9662 3526 9696 3556
rect 9696 3526 9711 3556
rect 9723 3556 9775 3578
rect 9723 3526 9734 3556
rect 9734 3526 9768 3556
rect 9768 3526 9775 3556
rect 9787 3556 9839 3578
rect 9851 3556 9903 3578
rect 9915 3556 9967 3578
rect 9979 3556 10031 3578
rect 10043 3556 10095 3578
rect 10107 3556 10159 3578
rect 10171 3556 10223 3578
rect 9787 3526 9806 3556
rect 9806 3526 9839 3556
rect 9851 3526 9878 3556
rect 9878 3526 9903 3556
rect 9915 3526 9950 3556
rect 9950 3526 9967 3556
rect 9979 3526 9984 3556
rect 9984 3526 10022 3556
rect 10022 3526 10031 3556
rect 10043 3526 10056 3556
rect 10056 3526 10094 3556
rect 10094 3526 10095 3556
rect 10107 3526 10128 3556
rect 10128 3526 10159 3556
rect 10171 3526 10200 3556
rect 10200 3526 10223 3556
rect 10235 3556 10287 3578
rect 10235 3526 10238 3556
rect 10238 3526 10272 3556
rect 10272 3526 10287 3556
rect 10299 3556 10351 3578
rect 10299 3526 10310 3556
rect 10310 3526 10344 3556
rect 10344 3526 10351 3556
rect 10363 3556 10415 3578
rect 10427 3556 10479 3578
rect 10491 3556 10543 3578
rect 10555 3556 10607 3578
rect 10619 3556 10671 3578
rect 10683 3556 10735 3578
rect 10747 3556 10799 3578
rect 10363 3526 10382 3556
rect 10382 3526 10415 3556
rect 10427 3526 10454 3556
rect 10454 3526 10479 3556
rect 10491 3526 10526 3556
rect 10526 3526 10543 3556
rect 10555 3526 10560 3556
rect 10560 3526 10598 3556
rect 10598 3526 10607 3556
rect 10619 3526 10632 3556
rect 10632 3526 10670 3556
rect 10670 3526 10671 3556
rect 10683 3526 10704 3556
rect 10704 3526 10735 3556
rect 10747 3526 10776 3556
rect 10776 3526 10799 3556
rect 10811 3556 10863 3578
rect 10811 3526 10814 3556
rect 10814 3526 10848 3556
rect 10848 3526 10863 3556
rect 3938 3358 3990 3410
rect 4020 3358 4072 3410
rect 4102 3358 4154 3410
rect 4184 3358 4236 3410
rect 3938 3292 3990 3344
rect 4020 3292 4072 3344
rect 4102 3292 4154 3344
rect 4184 3292 4236 3344
rect 3938 3226 3990 3278
rect 4020 3226 4072 3278
rect 4102 3226 4154 3278
rect 4184 3226 4236 3278
rect 3938 3160 3990 3212
rect 4020 3160 4072 3212
rect 4102 3160 4154 3212
rect 4184 3160 4236 3212
rect 3938 3094 3990 3146
rect 4020 3094 4072 3146
rect 4102 3094 4154 3146
rect 4184 3094 4236 3146
rect 1939 2926 2119 3042
rect 2132 2990 2184 3042
rect 2197 2990 2249 3042
rect 2262 2990 2314 3042
rect 2327 2990 2379 3042
rect 2392 2990 2444 3042
rect 2457 2990 2509 3042
rect 2522 2990 2574 3042
rect 2587 2990 2639 3042
rect 2652 2990 2704 3042
rect 2717 2990 2769 3042
rect 2782 2990 2834 3042
rect 2847 2990 2899 3042
rect 2912 2990 2964 3042
rect 2977 2990 3029 3042
rect 3042 2990 3094 3042
rect 3107 2990 3159 3042
rect 2132 2926 2184 2978
rect 2197 2926 2249 2978
rect 2262 2926 2314 2978
rect 2327 2926 2379 2978
rect 2392 2926 2444 2978
rect 2457 2926 2509 2978
rect 2522 2926 2574 2978
rect 2587 2926 2639 2978
rect 2652 2926 2704 2978
rect 2717 2926 2769 2978
rect 2782 2926 2834 2978
rect 2847 2926 2899 2978
rect 2912 2926 2964 2978
rect 2977 2926 3029 2978
rect 3042 2926 3094 2978
rect 1939 2862 2055 2926
rect 3107 2914 3223 2978
rect 2068 2862 2120 2914
rect 2133 2862 2185 2914
rect 2198 2862 2250 2914
rect 2263 2862 2315 2914
rect 2328 2862 2380 2914
rect 2393 2862 2445 2914
rect 2458 2862 2510 2914
rect 2523 2862 2575 2914
rect 2588 2862 2640 2914
rect 2653 2862 2705 2914
rect 2718 2862 2770 2914
rect 2783 2862 2835 2914
rect 2848 2862 2900 2914
rect 2913 2862 2965 2914
rect 2978 2862 3030 2914
rect 3043 2850 3223 2914
rect 1939 2798 1991 2850
rect 2004 2798 2056 2850
rect 2069 2798 2121 2850
rect 2134 2798 2186 2850
rect 2199 2798 2251 2850
rect 2264 2798 2316 2850
rect 2329 2798 2381 2850
rect 2394 2798 2446 2850
rect 2459 2798 2511 2850
rect 2524 2798 2576 2850
rect 2589 2798 2641 2850
rect 2654 2798 2706 2850
rect 2719 2798 2771 2850
rect 2784 2798 2836 2850
rect 2849 2798 2901 2850
rect 2914 2798 2966 2850
rect 2979 2786 3223 2850
rect 1939 2734 1991 2786
rect 2004 2734 2056 2786
rect 2069 2734 2121 2786
rect 2134 2734 2186 2786
rect 2199 2734 2251 2786
rect 2264 2734 2316 2786
rect 2329 2734 2381 2786
rect 2394 2734 2446 2786
rect 2459 2734 2511 2786
rect 2524 2734 2576 2786
rect 2589 2734 2641 2786
rect 2654 2734 2706 2786
rect 2719 2734 2771 2786
rect 2784 2734 2836 2786
rect 2849 2734 2901 2786
rect 2915 2722 3223 2786
rect 1939 2670 1991 2722
rect 2004 2670 2056 2722
rect 2069 2670 2121 2722
rect 2134 2670 2186 2722
rect 2199 2670 2251 2722
rect 2264 2670 2316 2722
rect 2329 2670 2381 2722
rect 2394 2670 2446 2722
rect 2459 2670 2511 2722
rect 2524 2670 2576 2722
rect 2589 2670 2641 2722
rect 2654 2670 2706 2722
rect 2719 2670 2771 2722
rect 2785 2670 2837 2722
rect 2851 2658 3223 2722
rect 1939 2606 1991 2658
rect 2004 2606 2056 2658
rect 2069 2606 2121 2658
rect 2134 2606 2186 2658
rect 2199 2606 2251 2658
rect 2264 2606 2316 2658
rect 2329 2606 2381 2658
rect 2394 2606 2446 2658
rect 2459 2606 2511 2658
rect 2524 2606 2576 2658
rect 2589 2606 2641 2658
rect 2655 2606 2707 2658
rect 2721 2606 2773 2658
rect 2787 2594 3223 2658
rect 1939 2542 1991 2594
rect 2004 2542 2056 2594
rect 2069 2542 2121 2594
rect 2134 2542 2186 2594
rect 2199 2542 2251 2594
rect 2264 2542 2316 2594
rect 2329 2542 2381 2594
rect 2394 2542 2446 2594
rect 2459 2542 2511 2594
rect 2525 2542 2577 2594
rect 2591 2542 2643 2594
rect 2657 2542 2709 2594
rect 2723 2530 3223 2594
rect 1939 2478 1991 2530
rect 2004 2478 2056 2530
rect 2069 2478 2121 2530
rect 2134 2478 2186 2530
rect 2199 2478 2251 2530
rect 2264 2478 2316 2530
rect 2329 2478 2381 2530
rect 2395 2478 2447 2530
rect 2461 2478 2513 2530
rect 2527 2478 2579 2530
rect 2593 2478 2645 2530
rect 1939 2414 1991 2466
rect 2004 2414 2056 2466
rect 2069 2414 2121 2466
rect 2134 2414 2186 2466
rect 2199 2414 2251 2466
rect 2265 2414 2317 2466
rect 2331 2414 2383 2466
rect 2397 2414 2449 2466
rect 2463 2414 2515 2466
rect 2529 2414 2581 2466
rect 2595 2414 2647 2466
rect 1939 2350 1991 2402
rect 2004 2350 2056 2402
rect 2069 2350 2121 2402
rect 2135 2350 2187 2402
rect 2201 2350 2253 2402
rect 2267 2350 2319 2402
rect 2333 2350 2385 2402
rect 2399 2350 2451 2402
rect 2465 2350 2517 2402
rect 2531 2350 2583 2402
rect 2595 2349 2647 2401
rect 2659 2350 3223 2530
rect 1939 2286 1991 2338
rect 2005 2286 2057 2338
rect 2071 2286 2123 2338
rect 2137 2286 2189 2338
rect 2203 2286 2255 2338
rect 2269 2286 2321 2338
rect 2335 2286 2387 2338
rect 2401 2286 2453 2338
rect 2467 2286 2519 2338
rect 2531 2285 2583 2337
rect 2595 2284 2647 2336
rect 2659 2285 2711 2337
rect 2723 2286 3223 2350
rect 1939 2222 1991 2274
rect 2005 2222 2057 2274
rect 2071 2222 2123 2274
rect 2137 2222 2189 2274
rect 2203 2222 2255 2274
rect 2269 2222 2321 2274
rect 2336 2222 2388 2274
rect 2403 2222 2455 2274
rect 2467 2221 2519 2273
rect 2531 2220 2583 2272
rect 2595 2219 2647 2271
rect 2659 2220 2711 2272
rect 2723 2221 2775 2273
rect 2787 2222 3223 2286
rect 2403 2157 2455 2209
rect 2467 2156 2519 2208
rect 2531 2155 2583 2207
rect 2595 2154 2647 2206
rect 2659 2155 2711 2207
rect 2723 2156 2775 2208
rect 2787 2157 2839 2209
rect 2851 2158 3223 2222
rect 2403 2092 2455 2144
rect 2467 2091 2519 2143
rect 2531 2090 2583 2142
rect 2595 2089 2647 2141
rect 2659 2090 2711 2142
rect 2723 2091 2775 2143
rect 2787 2092 2839 2144
rect 2851 2093 2903 2145
rect 2915 2094 3223 2158
rect 2403 2027 2455 2079
rect 2467 2026 2519 2078
rect 2531 2025 2583 2077
rect 2595 2024 2647 2076
rect 2659 2025 2711 2077
rect 2723 2026 2775 2078
rect 2787 2027 2839 2079
rect 2851 2028 2903 2080
rect 2915 2029 2967 2081
rect 2979 2030 3223 2094
rect 2403 1962 2455 2014
rect 2467 1961 2519 2013
rect 2531 1960 2583 2012
rect 2595 1959 2647 2011
rect 2659 1960 2711 2012
rect 2723 1961 2775 2013
rect 2787 1962 2839 2014
rect 2851 1963 2903 2015
rect 2915 1964 2967 2016
rect 2979 1965 3031 2017
rect 3043 1966 3223 2030
rect 3938 3027 3990 3079
rect 4020 3027 4072 3079
rect 4102 3027 4154 3079
rect 4184 3027 4236 3079
rect 3938 2960 3990 3012
rect 4020 2960 4072 3012
rect 4102 2960 4154 3012
rect 4184 2960 4236 3012
rect 3938 2893 3990 2945
rect 4020 2893 4072 2945
rect 4102 2893 4154 2945
rect 4184 2893 4236 2945
rect 3938 2826 3990 2878
rect 4020 2826 4072 2878
rect 4102 2826 4154 2878
rect 4184 2826 4236 2878
rect 3938 2759 3990 2811
rect 4020 2759 4072 2811
rect 4102 2759 4154 2811
rect 4184 2759 4236 2811
rect 3938 2692 3990 2744
rect 4020 2692 4072 2744
rect 4102 2692 4154 2744
rect 4184 2692 4236 2744
rect 3938 2625 3990 2677
rect 4020 2625 4072 2677
rect 4102 2625 4154 2677
rect 4184 2625 4236 2677
rect 3938 2558 3990 2610
rect 4020 2558 4072 2610
rect 4102 2558 4154 2610
rect 4184 2558 4236 2610
rect 3938 2491 3990 2543
rect 4020 2491 4072 2543
rect 4102 2491 4154 2543
rect 4184 2491 4236 2543
rect 3938 2424 3990 2476
rect 4020 2424 4072 2476
rect 4102 2424 4154 2476
rect 4184 2424 4236 2476
rect 3938 2357 3990 2409
rect 4020 2357 4072 2409
rect 4102 2357 4154 2409
rect 4184 2357 4236 2409
rect 3938 2290 3990 2342
rect 4020 2290 4072 2342
rect 4102 2290 4154 2342
rect 4184 2290 4236 2342
rect 3938 2223 3990 2275
rect 4020 2223 4072 2275
rect 4102 2223 4154 2275
rect 4184 2223 4236 2275
rect 3938 2156 3990 2208
rect 4020 2156 4072 2208
rect 4102 2156 4154 2208
rect 4184 2156 4236 2208
rect 3938 2089 3990 2141
rect 4020 2089 4072 2141
rect 4102 2089 4154 2141
rect 4184 2089 4236 2141
rect 3938 2022 3990 2074
rect 4020 2022 4072 2074
rect 4102 2022 4154 2074
rect 4184 2022 4236 2074
rect 4762 3358 4814 3410
rect 4844 3358 4896 3410
rect 4926 3358 4978 3410
rect 5008 3358 5060 3410
rect 4762 3292 4814 3344
rect 4844 3292 4896 3344
rect 4926 3292 4978 3344
rect 5008 3292 5060 3344
rect 4762 3226 4814 3278
rect 4844 3226 4896 3278
rect 4926 3226 4978 3278
rect 5008 3226 5060 3278
rect 4762 3160 4814 3212
rect 4844 3160 4896 3212
rect 4926 3160 4978 3212
rect 5008 3160 5060 3212
rect 4762 3094 4814 3146
rect 4844 3094 4896 3146
rect 4926 3094 4978 3146
rect 5008 3094 5060 3146
rect 4762 3027 4814 3079
rect 4844 3027 4896 3079
rect 4926 3027 4978 3079
rect 5008 3027 5060 3079
rect 4762 2960 4814 3012
rect 4844 2960 4896 3012
rect 4926 2960 4978 3012
rect 5008 2960 5060 3012
rect 4762 2893 4814 2945
rect 4844 2893 4896 2945
rect 4926 2893 4978 2945
rect 5008 2893 5060 2945
rect 4762 2826 4814 2878
rect 4844 2826 4896 2878
rect 4926 2826 4978 2878
rect 5008 2826 5060 2878
rect 4762 2759 4814 2811
rect 4844 2759 4896 2811
rect 4926 2759 4978 2811
rect 5008 2759 5060 2811
rect 4762 2692 4814 2744
rect 4844 2692 4896 2744
rect 4926 2692 4978 2744
rect 5008 2692 5060 2744
rect 4762 2625 4814 2677
rect 4844 2625 4896 2677
rect 4926 2625 4978 2677
rect 5008 2625 5060 2677
rect 4762 2558 4814 2610
rect 4844 2558 4896 2610
rect 4926 2558 4978 2610
rect 5008 2558 5060 2610
rect 4762 2491 4814 2543
rect 4844 2491 4896 2543
rect 4926 2491 4978 2543
rect 5008 2491 5060 2543
rect 4762 2424 4814 2476
rect 4844 2424 4896 2476
rect 4926 2424 4978 2476
rect 5008 2424 5060 2476
rect 4762 2357 4814 2409
rect 4844 2357 4896 2409
rect 4926 2357 4978 2409
rect 5008 2357 5060 2409
rect 4762 2290 4814 2342
rect 4844 2290 4896 2342
rect 4926 2290 4978 2342
rect 5008 2290 5060 2342
rect 4762 2223 4814 2275
rect 4844 2223 4896 2275
rect 4926 2223 4978 2275
rect 5008 2223 5060 2275
rect 4762 2156 4814 2208
rect 4844 2156 4896 2208
rect 4926 2156 4978 2208
rect 5008 2156 5060 2208
rect 4762 2089 4814 2141
rect 4844 2089 4896 2141
rect 4926 2089 4978 2141
rect 5008 2089 5060 2141
rect 4762 2022 4814 2074
rect 4844 2022 4896 2074
rect 4926 2022 4978 2074
rect 5008 2022 5060 2074
rect 5586 3358 5638 3410
rect 5668 3358 5720 3410
rect 5750 3358 5802 3410
rect 5832 3358 5884 3410
rect 5586 3292 5638 3344
rect 5668 3292 5720 3344
rect 5750 3292 5802 3344
rect 5832 3292 5884 3344
rect 5586 3226 5638 3278
rect 5668 3226 5720 3278
rect 5750 3226 5802 3278
rect 5832 3226 5884 3278
rect 5586 3160 5638 3212
rect 5668 3160 5720 3212
rect 5750 3160 5802 3212
rect 5832 3160 5884 3212
rect 5586 3094 5638 3146
rect 5668 3094 5720 3146
rect 5750 3094 5802 3146
rect 5832 3094 5884 3146
rect 5586 3027 5638 3079
rect 5668 3027 5720 3079
rect 5750 3027 5802 3079
rect 5832 3027 5884 3079
rect 5586 2960 5638 3012
rect 5668 2960 5720 3012
rect 5750 2960 5802 3012
rect 5832 2960 5884 3012
rect 5586 2893 5638 2945
rect 5668 2893 5720 2945
rect 5750 2893 5802 2945
rect 5832 2893 5884 2945
rect 5586 2826 5638 2878
rect 5668 2826 5720 2878
rect 5750 2826 5802 2878
rect 5832 2826 5884 2878
rect 5586 2759 5638 2811
rect 5668 2759 5720 2811
rect 5750 2759 5802 2811
rect 5832 2759 5884 2811
rect 5586 2692 5638 2744
rect 5668 2692 5720 2744
rect 5750 2692 5802 2744
rect 5832 2692 5884 2744
rect 5586 2625 5638 2677
rect 5668 2625 5720 2677
rect 5750 2625 5802 2677
rect 5832 2625 5884 2677
rect 5586 2558 5638 2610
rect 5668 2558 5720 2610
rect 5750 2558 5802 2610
rect 5832 2558 5884 2610
rect 5586 2491 5638 2543
rect 5668 2491 5720 2543
rect 5750 2491 5802 2543
rect 5832 2491 5884 2543
rect 5586 2424 5638 2476
rect 5668 2424 5720 2476
rect 5750 2424 5802 2476
rect 5832 2424 5884 2476
rect 5586 2357 5638 2409
rect 5668 2357 5720 2409
rect 5750 2357 5802 2409
rect 5832 2357 5884 2409
rect 5586 2290 5638 2342
rect 5668 2290 5720 2342
rect 5750 2290 5802 2342
rect 5832 2290 5884 2342
rect 5586 2223 5638 2275
rect 5668 2223 5720 2275
rect 5750 2223 5802 2275
rect 5832 2223 5884 2275
rect 5586 2156 5638 2208
rect 5668 2156 5720 2208
rect 5750 2156 5802 2208
rect 5832 2156 5884 2208
rect 5586 2089 5638 2141
rect 5668 2089 5720 2141
rect 5750 2089 5802 2141
rect 5832 2089 5884 2141
rect 5586 2022 5638 2074
rect 5668 2022 5720 2074
rect 5750 2022 5802 2074
rect 5832 2022 5884 2074
rect 6410 3358 6462 3410
rect 6492 3358 6544 3410
rect 6574 3358 6626 3410
rect 6656 3358 6708 3410
rect 6410 3292 6462 3344
rect 6492 3292 6544 3344
rect 6574 3292 6626 3344
rect 6656 3292 6708 3344
rect 6410 3226 6462 3278
rect 6492 3226 6544 3278
rect 6574 3226 6626 3278
rect 6656 3226 6708 3278
rect 6410 3160 6462 3212
rect 6492 3160 6544 3212
rect 6574 3160 6626 3212
rect 6656 3160 6708 3212
rect 6410 3094 6462 3146
rect 6492 3094 6544 3146
rect 6574 3094 6626 3146
rect 6656 3094 6708 3146
rect 6410 3027 6462 3079
rect 6492 3027 6544 3079
rect 6574 3027 6626 3079
rect 6656 3027 6708 3079
rect 6410 2960 6462 3012
rect 6492 2960 6544 3012
rect 6574 2960 6626 3012
rect 6656 2960 6708 3012
rect 6410 2893 6462 2945
rect 6492 2893 6544 2945
rect 6574 2893 6626 2945
rect 6656 2893 6708 2945
rect 6410 2826 6462 2878
rect 6492 2826 6544 2878
rect 6574 2826 6626 2878
rect 6656 2826 6708 2878
rect 6410 2759 6462 2811
rect 6492 2759 6544 2811
rect 6574 2759 6626 2811
rect 6656 2759 6708 2811
rect 6410 2692 6462 2744
rect 6492 2692 6544 2744
rect 6574 2692 6626 2744
rect 6656 2692 6708 2744
rect 6410 2625 6462 2677
rect 6492 2625 6544 2677
rect 6574 2625 6626 2677
rect 6656 2625 6708 2677
rect 6410 2558 6462 2610
rect 6492 2558 6544 2610
rect 6574 2558 6626 2610
rect 6656 2558 6708 2610
rect 6410 2491 6462 2543
rect 6492 2491 6544 2543
rect 6574 2491 6626 2543
rect 6656 2491 6708 2543
rect 6410 2424 6462 2476
rect 6492 2424 6544 2476
rect 6574 2424 6626 2476
rect 6656 2424 6708 2476
rect 6410 2357 6462 2409
rect 6492 2357 6544 2409
rect 6574 2357 6626 2409
rect 6656 2357 6708 2409
rect 6410 2290 6462 2342
rect 6492 2290 6544 2342
rect 6574 2290 6626 2342
rect 6656 2290 6708 2342
rect 6410 2223 6462 2275
rect 6492 2223 6544 2275
rect 6574 2223 6626 2275
rect 6656 2223 6708 2275
rect 6410 2156 6462 2208
rect 6492 2156 6544 2208
rect 6574 2156 6626 2208
rect 6656 2156 6708 2208
rect 6410 2089 6462 2141
rect 6492 2089 6544 2141
rect 6574 2089 6626 2141
rect 6656 2089 6708 2141
rect 6410 2022 6462 2074
rect 6492 2022 6544 2074
rect 6574 2022 6626 2074
rect 6656 2022 6708 2074
rect 7524 3358 7576 3410
rect 7606 3358 7658 3410
rect 7688 3358 7740 3410
rect 7770 3358 7822 3410
rect 7524 3292 7576 3344
rect 7606 3292 7658 3344
rect 7688 3292 7740 3344
rect 7770 3292 7822 3344
rect 7524 3226 7576 3278
rect 7606 3226 7658 3278
rect 7688 3226 7740 3278
rect 7770 3226 7822 3278
rect 7524 3160 7576 3212
rect 7606 3160 7658 3212
rect 7688 3160 7740 3212
rect 7770 3160 7822 3212
rect 7524 3094 7576 3146
rect 7606 3094 7658 3146
rect 7688 3094 7740 3146
rect 7770 3094 7822 3146
rect 7524 3027 7576 3079
rect 7606 3027 7658 3079
rect 7688 3027 7740 3079
rect 7770 3027 7822 3079
rect 7524 2960 7576 3012
rect 7606 2960 7658 3012
rect 7688 2960 7740 3012
rect 7770 2960 7822 3012
rect 7524 2893 7576 2945
rect 7606 2893 7658 2945
rect 7688 2893 7740 2945
rect 7770 2893 7822 2945
rect 7524 2826 7576 2878
rect 7606 2826 7658 2878
rect 7688 2826 7740 2878
rect 7770 2826 7822 2878
rect 7524 2759 7576 2811
rect 7606 2759 7658 2811
rect 7688 2759 7740 2811
rect 7770 2759 7822 2811
rect 7524 2692 7576 2744
rect 7606 2692 7658 2744
rect 7688 2692 7740 2744
rect 7770 2692 7822 2744
rect 7524 2625 7576 2677
rect 7606 2625 7658 2677
rect 7688 2625 7740 2677
rect 7770 2625 7822 2677
rect 7524 2558 7576 2610
rect 7606 2558 7658 2610
rect 7688 2558 7740 2610
rect 7770 2558 7822 2610
rect 7524 2491 7576 2543
rect 7606 2491 7658 2543
rect 7688 2491 7740 2543
rect 7770 2491 7822 2543
rect 7524 2424 7576 2476
rect 7606 2424 7658 2476
rect 7688 2424 7740 2476
rect 7770 2424 7822 2476
rect 7524 2357 7576 2409
rect 7606 2357 7658 2409
rect 7688 2357 7740 2409
rect 7770 2357 7822 2409
rect 7524 2290 7576 2342
rect 7606 2290 7658 2342
rect 7688 2290 7740 2342
rect 7770 2290 7822 2342
rect 7524 2223 7576 2275
rect 7606 2223 7658 2275
rect 7688 2223 7740 2275
rect 7770 2223 7822 2275
rect 7524 2156 7576 2208
rect 7606 2156 7658 2208
rect 7688 2156 7740 2208
rect 7770 2156 7822 2208
rect 7524 2089 7576 2141
rect 7606 2089 7658 2141
rect 7688 2089 7740 2141
rect 7770 2089 7822 2141
rect 7524 2022 7576 2074
rect 7606 2022 7658 2074
rect 7688 2022 7740 2074
rect 7770 2022 7822 2074
rect 8348 3358 8400 3410
rect 8430 3358 8482 3410
rect 8512 3358 8564 3410
rect 8594 3358 8646 3410
rect 8348 3292 8400 3344
rect 8430 3292 8482 3344
rect 8512 3292 8564 3344
rect 8594 3292 8646 3344
rect 8348 3226 8400 3278
rect 8430 3226 8482 3278
rect 8512 3226 8564 3278
rect 8594 3226 8646 3278
rect 8348 3160 8400 3212
rect 8430 3160 8482 3212
rect 8512 3160 8564 3212
rect 8594 3160 8646 3212
rect 8348 3094 8400 3146
rect 8430 3094 8482 3146
rect 8512 3094 8564 3146
rect 8594 3094 8646 3146
rect 8348 3027 8400 3079
rect 8430 3027 8482 3079
rect 8512 3027 8564 3079
rect 8594 3027 8646 3079
rect 8348 2960 8400 3012
rect 8430 2960 8482 3012
rect 8512 2960 8564 3012
rect 8594 2960 8646 3012
rect 8348 2893 8400 2945
rect 8430 2893 8482 2945
rect 8512 2893 8564 2945
rect 8594 2893 8646 2945
rect 8348 2826 8400 2878
rect 8430 2826 8482 2878
rect 8512 2826 8564 2878
rect 8594 2826 8646 2878
rect 8348 2759 8400 2811
rect 8430 2759 8482 2811
rect 8512 2759 8564 2811
rect 8594 2759 8646 2811
rect 8348 2692 8400 2744
rect 8430 2692 8482 2744
rect 8512 2692 8564 2744
rect 8594 2692 8646 2744
rect 8348 2625 8400 2677
rect 8430 2625 8482 2677
rect 8512 2625 8564 2677
rect 8594 2625 8646 2677
rect 8348 2558 8400 2610
rect 8430 2558 8482 2610
rect 8512 2558 8564 2610
rect 8594 2558 8646 2610
rect 8348 2491 8400 2543
rect 8430 2491 8482 2543
rect 8512 2491 8564 2543
rect 8594 2491 8646 2543
rect 8348 2424 8400 2476
rect 8430 2424 8482 2476
rect 8512 2424 8564 2476
rect 8594 2424 8646 2476
rect 8348 2357 8400 2409
rect 8430 2357 8482 2409
rect 8512 2357 8564 2409
rect 8594 2357 8646 2409
rect 8348 2290 8400 2342
rect 8430 2290 8482 2342
rect 8512 2290 8564 2342
rect 8594 2290 8646 2342
rect 8348 2223 8400 2275
rect 8430 2223 8482 2275
rect 8512 2223 8564 2275
rect 8594 2223 8646 2275
rect 8348 2156 8400 2208
rect 8430 2156 8482 2208
rect 8512 2156 8564 2208
rect 8594 2156 8646 2208
rect 8348 2089 8400 2141
rect 8430 2089 8482 2141
rect 8512 2089 8564 2141
rect 8594 2089 8646 2141
rect 8348 2022 8400 2074
rect 8430 2022 8482 2074
rect 8512 2022 8564 2074
rect 8594 2022 8646 2074
rect 9172 3358 9224 3410
rect 9254 3358 9306 3410
rect 9336 3358 9388 3410
rect 9418 3358 9470 3410
rect 9172 3292 9224 3344
rect 9254 3292 9306 3344
rect 9336 3292 9388 3344
rect 9418 3292 9470 3344
rect 9172 3226 9224 3278
rect 9254 3226 9306 3278
rect 9336 3226 9388 3278
rect 9418 3226 9470 3278
rect 9172 3160 9224 3212
rect 9254 3160 9306 3212
rect 9336 3160 9388 3212
rect 9418 3160 9470 3212
rect 9172 3094 9224 3146
rect 9254 3094 9306 3146
rect 9336 3094 9388 3146
rect 9418 3094 9470 3146
rect 9172 3027 9224 3079
rect 9254 3027 9306 3079
rect 9336 3027 9388 3079
rect 9418 3027 9470 3079
rect 9172 2960 9224 3012
rect 9254 2960 9306 3012
rect 9336 2960 9388 3012
rect 9418 2960 9470 3012
rect 9172 2893 9224 2945
rect 9254 2893 9306 2945
rect 9336 2893 9388 2945
rect 9418 2893 9470 2945
rect 9172 2826 9224 2878
rect 9254 2826 9306 2878
rect 9336 2826 9388 2878
rect 9418 2826 9470 2878
rect 9172 2759 9224 2811
rect 9254 2759 9306 2811
rect 9336 2759 9388 2811
rect 9418 2759 9470 2811
rect 9172 2692 9224 2744
rect 9254 2692 9306 2744
rect 9336 2692 9388 2744
rect 9418 2692 9470 2744
rect 9172 2625 9224 2677
rect 9254 2625 9306 2677
rect 9336 2625 9388 2677
rect 9418 2625 9470 2677
rect 9172 2558 9224 2610
rect 9254 2558 9306 2610
rect 9336 2558 9388 2610
rect 9418 2558 9470 2610
rect 9172 2491 9224 2543
rect 9254 2491 9306 2543
rect 9336 2491 9388 2543
rect 9418 2491 9470 2543
rect 9172 2424 9224 2476
rect 9254 2424 9306 2476
rect 9336 2424 9388 2476
rect 9418 2424 9470 2476
rect 9172 2357 9224 2409
rect 9254 2357 9306 2409
rect 9336 2357 9388 2409
rect 9418 2357 9470 2409
rect 9172 2290 9224 2342
rect 9254 2290 9306 2342
rect 9336 2290 9388 2342
rect 9418 2290 9470 2342
rect 9172 2223 9224 2275
rect 9254 2223 9306 2275
rect 9336 2223 9388 2275
rect 9418 2223 9470 2275
rect 9172 2156 9224 2208
rect 9254 2156 9306 2208
rect 9336 2156 9388 2208
rect 9418 2156 9470 2208
rect 9172 2089 9224 2141
rect 9254 2089 9306 2141
rect 9336 2089 9388 2141
rect 9418 2089 9470 2141
rect 9172 2022 9224 2074
rect 9254 2022 9306 2074
rect 9336 2022 9388 2074
rect 9418 2022 9470 2074
rect 9996 3358 10048 3410
rect 10078 3358 10130 3410
rect 10160 3358 10212 3410
rect 10242 3358 10294 3410
rect 9996 3292 10048 3344
rect 10078 3292 10130 3344
rect 10160 3292 10212 3344
rect 10242 3292 10294 3344
rect 9996 3226 10048 3278
rect 10078 3226 10130 3278
rect 10160 3226 10212 3278
rect 10242 3226 10294 3278
rect 9996 3160 10048 3212
rect 10078 3160 10130 3212
rect 10160 3160 10212 3212
rect 10242 3160 10294 3212
rect 9996 3094 10048 3146
rect 10078 3094 10130 3146
rect 10160 3094 10212 3146
rect 10242 3094 10294 3146
rect 9996 3027 10048 3079
rect 10078 3027 10130 3079
rect 10160 3027 10212 3079
rect 10242 3027 10294 3079
rect 9996 2960 10048 3012
rect 10078 2960 10130 3012
rect 10160 2960 10212 3012
rect 10242 2960 10294 3012
rect 9996 2893 10048 2945
rect 10078 2893 10130 2945
rect 10160 2893 10212 2945
rect 10242 2893 10294 2945
rect 9996 2826 10048 2878
rect 10078 2826 10130 2878
rect 10160 2826 10212 2878
rect 10242 2826 10294 2878
rect 9996 2759 10048 2811
rect 10078 2759 10130 2811
rect 10160 2759 10212 2811
rect 10242 2759 10294 2811
rect 9996 2692 10048 2744
rect 10078 2692 10130 2744
rect 10160 2692 10212 2744
rect 10242 2692 10294 2744
rect 9996 2625 10048 2677
rect 10078 2625 10130 2677
rect 10160 2625 10212 2677
rect 10242 2625 10294 2677
rect 9996 2558 10048 2610
rect 10078 2558 10130 2610
rect 10160 2558 10212 2610
rect 10242 2558 10294 2610
rect 9996 2491 10048 2543
rect 10078 2491 10130 2543
rect 10160 2491 10212 2543
rect 10242 2491 10294 2543
rect 9996 2424 10048 2476
rect 10078 2424 10130 2476
rect 10160 2424 10212 2476
rect 10242 2424 10294 2476
rect 9996 2357 10048 2409
rect 10078 2357 10130 2409
rect 10160 2357 10212 2409
rect 10242 2357 10294 2409
rect 9996 2290 10048 2342
rect 10078 2290 10130 2342
rect 10160 2290 10212 2342
rect 10242 2290 10294 2342
rect 9996 2223 10048 2275
rect 10078 2223 10130 2275
rect 10160 2223 10212 2275
rect 10242 2223 10294 2275
rect 9996 2156 10048 2208
rect 10078 2156 10130 2208
rect 10160 2156 10212 2208
rect 10242 2156 10294 2208
rect 9996 2089 10048 2141
rect 10078 2089 10130 2141
rect 10160 2089 10212 2141
rect 10242 2089 10294 2141
rect 9996 2022 10048 2074
rect 10078 2022 10130 2074
rect 10160 2022 10212 2074
rect 10242 2022 10294 2074
rect 10820 3358 10872 3410
rect 10902 3358 10954 3410
rect 10984 3358 11036 3410
rect 11066 3358 11118 3410
rect 10820 3292 10872 3344
rect 10902 3292 10954 3344
rect 10984 3292 11036 3344
rect 11066 3292 11118 3344
rect 10820 3226 10872 3278
rect 10902 3226 10954 3278
rect 10984 3226 11036 3278
rect 11066 3226 11118 3278
rect 10820 3160 10872 3212
rect 10902 3160 10954 3212
rect 10984 3160 11036 3212
rect 11066 3160 11118 3212
rect 10820 3094 10872 3146
rect 10902 3094 10954 3146
rect 10984 3094 11036 3146
rect 11066 3094 11118 3146
rect 10820 3027 10872 3079
rect 10902 3027 10954 3079
rect 10984 3027 11036 3079
rect 11066 3027 11118 3079
rect 10820 2960 10872 3012
rect 10902 2960 10954 3012
rect 10984 2960 11036 3012
rect 11066 2960 11118 3012
rect 10820 2893 10872 2945
rect 10902 2893 10954 2945
rect 10984 2893 11036 2945
rect 11066 2893 11118 2945
rect 10820 2826 10872 2878
rect 10902 2826 10954 2878
rect 10984 2826 11036 2878
rect 11066 2826 11118 2878
rect 10820 2759 10872 2811
rect 10902 2759 10954 2811
rect 10984 2759 11036 2811
rect 11066 2759 11118 2811
rect 10820 2692 10872 2744
rect 10902 2692 10954 2744
rect 10984 2692 11036 2744
rect 11066 2692 11118 2744
rect 10820 2625 10872 2677
rect 10902 2625 10954 2677
rect 10984 2625 11036 2677
rect 11066 2625 11118 2677
rect 10820 2558 10872 2610
rect 10902 2558 10954 2610
rect 10984 2558 11036 2610
rect 11066 2558 11118 2610
rect 10820 2491 10872 2543
rect 10902 2491 10954 2543
rect 10984 2491 11036 2543
rect 11066 2491 11118 2543
rect 10820 2424 10872 2476
rect 10902 2424 10954 2476
rect 10984 2424 11036 2476
rect 11066 2424 11118 2476
rect 10820 2357 10872 2409
rect 10902 2357 10954 2409
rect 10984 2357 11036 2409
rect 11066 2357 11118 2409
rect 10820 2290 10872 2342
rect 10902 2290 10954 2342
rect 10984 2290 11036 2342
rect 11066 2290 11118 2342
rect 10820 2223 10872 2275
rect 10902 2223 10954 2275
rect 10984 2223 11036 2275
rect 11066 2223 11118 2275
rect 10820 2156 10872 2208
rect 10902 2156 10954 2208
rect 10984 2156 11036 2208
rect 11066 2156 11118 2208
rect 10820 2089 10872 2141
rect 10902 2089 10954 2141
rect 10984 2089 11036 2141
rect 11066 2089 11118 2141
rect 10820 2022 10872 2074
rect 10902 2022 10954 2074
rect 10984 2022 11036 2074
rect 11066 2022 11118 2074
rect 2403 1897 2455 1949
rect 2467 1896 2519 1948
rect 2531 1895 2583 1947
rect 2595 1894 2647 1946
rect 2659 1895 2711 1947
rect 2723 1896 2775 1948
rect 2787 1897 2839 1949
rect 2851 1898 2903 1950
rect 2915 1899 2967 1951
rect 2979 1900 3031 1952
rect 3043 1901 3095 1953
rect 3107 1902 3223 1966
rect 2403 1832 2455 1884
rect 2467 1831 2519 1883
rect 2531 1830 2583 1882
rect 2595 1829 2647 1881
rect 2659 1830 2711 1882
rect 2723 1831 2775 1883
rect 2787 1832 2839 1884
rect 2851 1833 2903 1885
rect 2915 1834 2967 1886
rect 2979 1835 3031 1887
rect 3043 1836 3095 1888
rect 3107 1837 3159 1889
rect 3171 1837 3223 1889
rect 2403 1766 2455 1818
rect 2467 1766 2519 1818
rect 2531 1765 2583 1817
rect 2595 1764 2647 1816
rect 2659 1765 2711 1817
rect 2723 1766 2775 1818
rect 2787 1767 2839 1819
rect 2851 1768 2903 1820
rect 2915 1769 2967 1821
rect 2979 1770 3031 1822
rect 3043 1771 3095 1823
rect 3107 1772 3159 1824
rect 3171 1772 3223 1824
rect 2403 1700 2455 1752
rect 2467 1701 2519 1753
rect 2531 1700 2583 1752
rect 2595 1699 2647 1751
rect 2659 1700 2711 1752
rect 2723 1701 2775 1753
rect 2787 1702 2839 1754
rect 2851 1703 2903 1755
rect 2915 1704 2967 1756
rect 2979 1705 3031 1757
rect 3043 1706 3095 1758
rect 3107 1707 3159 1759
rect 3171 1707 3223 1759
rect 2403 1634 2455 1686
rect 2467 1636 2519 1688
rect 2531 1635 2583 1687
rect 2595 1634 2647 1686
rect 2659 1635 2711 1687
rect 2723 1636 2775 1688
rect 2787 1637 2839 1689
rect 2851 1638 2903 1690
rect 2915 1639 2967 1691
rect 2979 1640 3031 1692
rect 3043 1641 3095 1693
rect 3107 1642 3159 1694
rect 3171 1642 3223 1694
rect 2403 1568 2455 1620
rect 2467 1570 2519 1622
rect 2531 1570 2583 1622
rect 2595 1569 2647 1621
rect 2659 1570 2711 1622
rect 2723 1571 2775 1623
rect 2787 1572 2839 1624
rect 2851 1573 2903 1625
rect 2915 1574 2967 1626
rect 2979 1575 3031 1627
rect 3043 1576 3095 1628
rect 3107 1577 3159 1629
rect 3171 1577 3223 1629
rect 2403 1502 2455 1554
rect 2467 1504 2519 1556
rect 2531 1505 2583 1557
rect 2595 1504 2647 1556
rect 2659 1505 2711 1557
rect 2723 1506 2775 1558
rect 2787 1507 2839 1559
rect 2851 1508 2903 1560
rect 2915 1509 2967 1561
rect 2979 1510 3031 1562
rect 3043 1511 3095 1563
rect 3107 1512 3159 1564
rect 3171 1512 3223 1564
rect 1939 1436 1991 1488
rect 2006 1436 2058 1488
rect 2073 1436 2125 1488
rect 2139 1436 2191 1488
rect 2205 1436 2257 1488
rect 2271 1436 2323 1488
rect 2337 1436 2389 1488
rect 2403 1436 2455 1488
rect 2467 1438 2519 1490
rect 2531 1440 2583 1492
rect 2595 1439 2647 1491
rect 2659 1440 2711 1492
rect 2723 1441 2775 1493
rect 2787 1442 2839 1494
rect 2851 1443 2903 1495
rect 2915 1444 2967 1496
rect 2979 1445 3031 1497
rect 3043 1446 3095 1498
rect 3107 1447 3159 1499
rect 3171 1447 3223 1499
rect 1939 1372 1991 1424
rect 2005 1372 2057 1424
rect 2071 1372 2123 1424
rect 2137 1372 2189 1424
rect 2203 1372 2255 1424
rect 2269 1372 2321 1424
rect 2335 1372 2387 1424
rect 2401 1372 2453 1424
rect 2467 1372 2519 1424
rect 2531 1374 2583 1426
rect 2595 1374 2647 1426
rect 2659 1375 2711 1427
rect 2723 1376 2775 1428
rect 2787 1377 2839 1429
rect 2851 1378 2903 1430
rect 2915 1379 2967 1431
rect 2979 1380 3031 1432
rect 3043 1381 3095 1433
rect 3107 1382 3159 1434
rect 3171 1382 3223 1434
rect 1939 1308 1991 1360
rect 2005 1308 2057 1360
rect 2071 1308 2123 1360
rect 2137 1308 2189 1360
rect 2203 1308 2255 1360
rect 2269 1308 2321 1360
rect 2335 1308 2387 1360
rect 2401 1308 2453 1360
rect 2466 1308 2518 1360
rect 2531 1308 2583 1360
rect 2595 1309 2647 1361
rect 2659 1310 2711 1362
rect 2723 1311 2775 1363
rect 2787 1312 2839 1364
rect 2851 1313 2903 1365
rect 2915 1314 2967 1366
rect 2979 1315 3031 1367
rect 3043 1316 3095 1368
rect 3107 1317 3159 1369
rect 3171 1317 3223 1369
rect 1939 1244 1991 1296
rect 2005 1244 2057 1296
rect 2071 1244 2123 1296
rect 2137 1244 2189 1296
rect 2203 1244 2255 1296
rect 2269 1244 2321 1296
rect 2335 1244 2387 1296
rect 2400 1244 2452 1296
rect 2465 1244 2517 1296
rect 2530 1244 2582 1296
rect 2595 1244 2647 1296
rect 2659 1245 2711 1297
rect 2723 1246 2775 1298
rect 2787 1247 2839 1299
rect 2851 1248 2903 1300
rect 2915 1249 2967 1301
rect 2979 1250 3031 1302
rect 3043 1251 3095 1303
rect 3107 1252 3159 1304
rect 3171 1252 3223 1304
rect 1939 1180 1991 1232
rect 2005 1180 2057 1232
rect 2071 1180 2123 1232
rect 2137 1180 2189 1232
rect 2203 1180 2255 1232
rect 2269 1180 2321 1232
rect 2334 1180 2386 1232
rect 2399 1180 2451 1232
rect 2464 1180 2516 1232
rect 2529 1180 2581 1232
rect 2594 1180 2646 1232
rect 2659 1180 2711 1232
rect 2723 1181 2775 1233
rect 2787 1182 2839 1234
rect 2851 1183 2903 1235
rect 2915 1184 2967 1236
rect 2979 1185 3031 1237
rect 3043 1186 3095 1238
rect 3107 1187 3159 1239
rect 3171 1187 3223 1239
rect 1939 1116 1991 1168
rect 2005 1116 2057 1168
rect 2071 1116 2123 1168
rect 2137 1116 2189 1168
rect 2203 1116 2255 1168
rect 2268 1116 2320 1168
rect 2333 1116 2385 1168
rect 2398 1116 2450 1168
rect 2463 1116 2515 1168
rect 2528 1116 2580 1168
rect 2593 1116 2645 1168
rect 2658 1116 2710 1168
rect 2723 1116 2775 1168
rect 2787 1117 2839 1169
rect 2851 1118 2903 1170
rect 2915 1119 2967 1171
rect 2979 1120 3031 1172
rect 3043 1121 3095 1173
rect 3107 1122 3159 1174
rect 3171 1122 3223 1174
rect 1939 1052 1991 1104
rect 2005 1052 2057 1104
rect 2071 1052 2123 1104
rect 2137 1052 2189 1104
rect 2202 1052 2254 1104
rect 2267 1052 2319 1104
rect 2332 1052 2384 1104
rect 2397 1052 2449 1104
rect 2462 1052 2514 1104
rect 2527 1052 2579 1104
rect 2592 1052 2644 1104
rect 2657 1052 2709 1104
rect 2722 1052 2774 1104
rect 2787 1052 2839 1104
rect 2851 1053 2903 1105
rect 2915 1054 2967 1106
rect 2979 1055 3031 1107
rect 3043 1056 3095 1108
rect 3107 1057 3159 1109
rect 3171 1057 3223 1109
rect 1939 988 1991 1040
rect 2005 988 2057 1040
rect 2071 988 2123 1040
rect 2136 988 2188 1040
rect 2201 988 2253 1040
rect 2266 988 2318 1040
rect 2331 988 2383 1040
rect 2396 988 2448 1040
rect 2461 988 2513 1040
rect 2526 988 2578 1040
rect 2591 988 2643 1040
rect 2656 988 2708 1040
rect 2721 988 2773 1040
rect 2786 988 2838 1040
rect 2851 988 2903 1040
rect 2915 989 2967 1041
rect 2979 990 3031 1042
rect 3043 991 3095 1043
rect 3107 992 3159 1044
rect 3171 992 3223 1044
rect 3526 1850 3578 1902
rect 3608 1850 3660 1902
rect 3690 1850 3742 1902
rect 3772 1850 3824 1902
rect 3526 1782 3578 1834
rect 3608 1782 3660 1834
rect 3690 1782 3742 1834
rect 3772 1782 3824 1834
rect 3526 1714 3578 1766
rect 3608 1714 3660 1766
rect 3690 1714 3742 1766
rect 3772 1714 3824 1766
rect 3526 1646 3578 1698
rect 3608 1646 3660 1698
rect 3690 1646 3742 1698
rect 3772 1646 3824 1698
rect 3526 1578 3578 1630
rect 3608 1578 3660 1630
rect 3690 1578 3742 1630
rect 3772 1578 3824 1630
rect 3526 1510 3578 1562
rect 3608 1510 3660 1562
rect 3690 1510 3742 1562
rect 3772 1510 3824 1562
rect 3526 1442 3578 1494
rect 3608 1442 3660 1494
rect 3690 1442 3742 1494
rect 3772 1442 3824 1494
rect 3526 1374 3578 1426
rect 3608 1374 3660 1426
rect 3690 1374 3742 1426
rect 3772 1374 3824 1426
rect 3526 1306 3578 1358
rect 3608 1306 3660 1358
rect 3690 1306 3742 1358
rect 3772 1306 3824 1358
rect 3526 1237 3578 1289
rect 3608 1237 3660 1289
rect 3690 1237 3742 1289
rect 3772 1237 3824 1289
rect 3526 1168 3578 1220
rect 3608 1168 3660 1220
rect 3690 1168 3742 1220
rect 3772 1168 3824 1220
rect 3526 1099 3578 1151
rect 3608 1099 3660 1151
rect 3690 1099 3742 1151
rect 3772 1099 3824 1151
rect 3526 1030 3578 1082
rect 3608 1030 3660 1082
rect 3690 1030 3742 1082
rect 3772 1030 3824 1082
rect 4350 1850 4402 1902
rect 4432 1850 4484 1902
rect 4514 1850 4566 1902
rect 4596 1850 4648 1902
rect 4350 1786 4402 1838
rect 4432 1786 4484 1838
rect 4514 1786 4566 1838
rect 4596 1786 4648 1838
rect 4350 1722 4402 1774
rect 4432 1722 4484 1774
rect 4514 1722 4566 1774
rect 4596 1722 4648 1774
rect 4350 1658 4402 1710
rect 4432 1658 4484 1710
rect 4514 1658 4566 1710
rect 4596 1658 4648 1710
rect 4350 1594 4402 1646
rect 4432 1594 4484 1646
rect 4514 1594 4566 1646
rect 4596 1594 4648 1646
rect 4350 1530 4402 1582
rect 4432 1530 4484 1582
rect 4514 1530 4566 1582
rect 4596 1530 4648 1582
rect 4350 1466 4402 1518
rect 4432 1466 4484 1518
rect 4514 1466 4566 1518
rect 4596 1466 4648 1518
rect 4350 1402 4402 1454
rect 4432 1402 4484 1454
rect 4514 1402 4566 1454
rect 4596 1402 4648 1454
rect 4350 1338 4402 1390
rect 4432 1338 4484 1390
rect 4514 1338 4566 1390
rect 4596 1338 4648 1390
rect 4350 1274 4402 1326
rect 4432 1274 4484 1326
rect 4514 1274 4566 1326
rect 4596 1274 4648 1326
rect 4350 1210 4402 1262
rect 4432 1210 4484 1262
rect 4514 1210 4566 1262
rect 4596 1210 4648 1262
rect 4350 1146 4402 1198
rect 4432 1146 4484 1198
rect 4514 1146 4566 1198
rect 4596 1146 4648 1198
rect 4350 1082 4402 1134
rect 4432 1082 4484 1134
rect 4514 1082 4566 1134
rect 4596 1082 4648 1134
rect 4350 1018 4402 1070
rect 4432 1018 4484 1070
rect 4514 1018 4566 1070
rect 4596 1018 4648 1070
rect 1939 924 1991 976
rect 2005 924 2057 976
rect 2070 924 2122 976
rect 2135 924 2187 976
rect 2200 924 2252 976
rect 2265 924 2317 976
rect 2330 924 2382 976
rect 2395 924 2447 976
rect 2460 924 2512 976
rect 2525 924 2577 976
rect 2590 924 2642 976
rect 2655 924 2707 976
rect 2720 924 2772 976
rect 2785 924 2837 976
rect 2850 924 2902 976
rect 2915 924 2967 976
rect 2979 925 3031 977
rect 3043 926 3095 978
rect 3107 927 3159 979
rect 3171 927 3223 979
rect 3590 966 3642 1018
rect 3678 966 3730 1018
rect 3766 966 3818 1018
rect 4350 954 4402 1006
rect 4432 954 4484 1006
rect 4514 954 4566 1006
rect 4596 954 4648 1006
rect 1939 860 1991 912
rect 2004 860 2056 912
rect 2069 860 2121 912
rect 2134 860 2186 912
rect 2199 860 2251 912
rect 2264 860 2316 912
rect 2329 860 2381 912
rect 2394 860 2446 912
rect 2459 860 2511 912
rect 2524 860 2576 912
rect 2589 860 2641 912
rect 2654 860 2706 912
rect 2719 860 2771 912
rect 2784 860 2836 912
rect 2849 860 2901 912
rect 2914 860 2966 912
rect 2979 860 3031 912
rect 3043 861 3095 913
rect 3107 862 3159 914
rect 3171 862 3223 914
rect 3660 901 3712 953
rect 3766 901 3818 953
rect 4350 890 4402 942
rect 4432 890 4484 942
rect 4514 890 4566 942
rect 4596 890 4648 942
rect 1939 796 1991 848
rect 2004 796 2056 848
rect 2069 796 2121 848
rect 2134 796 2186 848
rect 2199 796 2251 848
rect 2264 796 2316 848
rect 2329 796 2381 848
rect 2394 796 2446 848
rect 2459 796 2511 848
rect 2524 796 2576 848
rect 2589 796 2641 848
rect 2654 796 2706 848
rect 2719 796 2771 848
rect 2784 796 2836 848
rect 2849 796 2901 848
rect 2914 796 2966 848
rect 2979 784 3095 848
rect 3107 797 3159 849
rect 3171 797 3223 849
rect 3753 815 3805 867
rect 4350 826 4402 878
rect 4432 826 4484 878
rect 4514 826 4566 878
rect 4596 826 4648 878
rect 1939 732 1991 784
rect 2004 732 2056 784
rect 2069 732 2121 784
rect 2134 732 2186 784
rect 2199 732 2251 784
rect 2264 732 2316 784
rect 2329 732 2381 784
rect 2394 732 2446 784
rect 2459 732 2511 784
rect 2524 732 2576 784
rect 2589 732 2641 784
rect 2654 732 2706 784
rect 2719 732 2771 784
rect 2784 732 2836 784
rect 2849 732 2901 784
rect 2914 732 2966 784
rect 1939 668 1991 720
rect 2004 668 2056 720
rect 2069 668 2121 720
rect 2134 668 2186 720
rect 2199 668 2251 720
rect 2264 668 2316 720
rect 2329 668 2381 720
rect 2394 668 2446 720
rect 2459 668 2511 720
rect 2524 668 2576 720
rect 2589 668 2641 720
rect 2654 668 2706 720
rect 2719 668 2771 720
rect 2784 668 2836 720
rect 2849 668 2901 720
rect 2914 668 2966 720
rect 2979 668 3159 784
rect 3171 732 3223 784
rect 4350 762 4402 814
rect 4432 762 4484 814
rect 4514 762 4566 814
rect 4596 762 4648 814
rect 4350 698 4402 750
rect 4432 698 4484 750
rect 4514 698 4566 750
rect 4596 698 4648 750
rect 4350 633 4402 685
rect 4432 633 4484 685
rect 4514 633 4566 685
rect 4596 633 4648 685
rect 4350 568 4402 620
rect 4432 568 4484 620
rect 4514 568 4566 620
rect 4596 568 4648 620
rect 4350 503 4402 555
rect 4432 503 4484 555
rect 4514 503 4566 555
rect 4596 503 4648 555
rect 4350 438 4402 490
rect 4432 438 4484 490
rect 4514 438 4566 490
rect 4596 438 4648 490
rect 4350 373 4402 425
rect 4432 373 4484 425
rect 4514 373 4566 425
rect 4596 373 4648 425
rect 5174 1850 5226 1902
rect 5256 1850 5308 1902
rect 5338 1850 5390 1902
rect 5420 1850 5472 1902
rect 5174 1786 5226 1838
rect 5256 1786 5308 1838
rect 5338 1786 5390 1838
rect 5420 1786 5472 1838
rect 5174 1722 5226 1774
rect 5256 1722 5308 1774
rect 5338 1722 5390 1774
rect 5420 1722 5472 1774
rect 5174 1658 5226 1710
rect 5256 1658 5308 1710
rect 5338 1658 5390 1710
rect 5420 1658 5472 1710
rect 5174 1594 5226 1646
rect 5256 1594 5308 1646
rect 5338 1594 5390 1646
rect 5420 1594 5472 1646
rect 5174 1530 5226 1582
rect 5256 1530 5308 1582
rect 5338 1530 5390 1582
rect 5420 1530 5472 1582
rect 5174 1466 5226 1518
rect 5256 1466 5308 1518
rect 5338 1466 5390 1518
rect 5420 1466 5472 1518
rect 5174 1402 5226 1454
rect 5256 1402 5308 1454
rect 5338 1402 5390 1454
rect 5420 1402 5472 1454
rect 5174 1338 5226 1390
rect 5256 1338 5308 1390
rect 5338 1338 5390 1390
rect 5420 1338 5472 1390
rect 5174 1274 5226 1326
rect 5256 1274 5308 1326
rect 5338 1274 5390 1326
rect 5420 1274 5472 1326
rect 5174 1210 5226 1262
rect 5256 1210 5308 1262
rect 5338 1210 5390 1262
rect 5420 1210 5472 1262
rect 5174 1146 5226 1198
rect 5256 1146 5308 1198
rect 5338 1146 5390 1198
rect 5420 1146 5472 1198
rect 5174 1082 5226 1134
rect 5256 1082 5308 1134
rect 5338 1082 5390 1134
rect 5420 1082 5472 1134
rect 5174 1018 5226 1070
rect 5256 1018 5308 1070
rect 5338 1018 5390 1070
rect 5420 1018 5472 1070
rect 5174 954 5226 1006
rect 5256 954 5308 1006
rect 5338 954 5390 1006
rect 5420 954 5472 1006
rect 5174 890 5226 942
rect 5256 890 5308 942
rect 5338 890 5390 942
rect 5420 890 5472 942
rect 5174 826 5226 878
rect 5256 826 5308 878
rect 5338 826 5390 878
rect 5420 826 5472 878
rect 5174 762 5226 814
rect 5256 762 5308 814
rect 5338 762 5390 814
rect 5420 762 5472 814
rect 5174 698 5226 750
rect 5256 698 5308 750
rect 5338 698 5390 750
rect 5420 698 5472 750
rect 5174 633 5226 685
rect 5256 633 5308 685
rect 5338 633 5390 685
rect 5420 633 5472 685
rect 5174 568 5226 620
rect 5256 568 5308 620
rect 5338 568 5390 620
rect 5420 568 5472 620
rect 5174 503 5226 555
rect 5256 503 5308 555
rect 5338 503 5390 555
rect 5420 503 5472 555
rect 5174 438 5226 490
rect 5256 438 5308 490
rect 5338 438 5390 490
rect 5420 438 5472 490
rect 5174 373 5226 425
rect 5256 373 5308 425
rect 5338 373 5390 425
rect 5420 373 5472 425
rect 5998 1850 6050 1902
rect 6080 1850 6132 1902
rect 6162 1850 6214 1902
rect 6244 1850 6296 1902
rect 5998 1786 6050 1838
rect 6080 1786 6132 1838
rect 6162 1786 6214 1838
rect 6244 1786 6296 1838
rect 5998 1722 6050 1774
rect 6080 1722 6132 1774
rect 6162 1722 6214 1774
rect 6244 1722 6296 1774
rect 5998 1658 6050 1710
rect 6080 1658 6132 1710
rect 6162 1658 6214 1710
rect 6244 1658 6296 1710
rect 5998 1594 6050 1646
rect 6080 1594 6132 1646
rect 6162 1594 6214 1646
rect 6244 1594 6296 1646
rect 5998 1530 6050 1582
rect 6080 1530 6132 1582
rect 6162 1530 6214 1582
rect 6244 1530 6296 1582
rect 5998 1466 6050 1518
rect 6080 1466 6132 1518
rect 6162 1466 6214 1518
rect 6244 1466 6296 1518
rect 5998 1402 6050 1454
rect 6080 1402 6132 1454
rect 6162 1402 6214 1454
rect 6244 1402 6296 1454
rect 5998 1338 6050 1390
rect 6080 1338 6132 1390
rect 6162 1338 6214 1390
rect 6244 1338 6296 1390
rect 5998 1274 6050 1326
rect 6080 1274 6132 1326
rect 6162 1274 6214 1326
rect 6244 1274 6296 1326
rect 5998 1210 6050 1262
rect 6080 1210 6132 1262
rect 6162 1210 6214 1262
rect 6244 1210 6296 1262
rect 5998 1146 6050 1198
rect 6080 1146 6132 1198
rect 6162 1146 6214 1198
rect 6244 1146 6296 1198
rect 5998 1082 6050 1134
rect 6080 1082 6132 1134
rect 6162 1082 6214 1134
rect 6244 1082 6296 1134
rect 5998 1018 6050 1070
rect 6080 1018 6132 1070
rect 6162 1018 6214 1070
rect 6244 1018 6296 1070
rect 5998 954 6050 1006
rect 6080 954 6132 1006
rect 6162 954 6214 1006
rect 6244 954 6296 1006
rect 5998 890 6050 942
rect 6080 890 6132 942
rect 6162 890 6214 942
rect 6244 890 6296 942
rect 5998 826 6050 878
rect 6080 826 6132 878
rect 6162 826 6214 878
rect 6244 826 6296 878
rect 5998 762 6050 814
rect 6080 762 6132 814
rect 6162 762 6214 814
rect 6244 762 6296 814
rect 5998 698 6050 750
rect 6080 698 6132 750
rect 6162 698 6214 750
rect 6244 698 6296 750
rect 5998 633 6050 685
rect 6080 633 6132 685
rect 6162 633 6214 685
rect 6244 633 6296 685
rect 5998 568 6050 620
rect 6080 568 6132 620
rect 6162 568 6214 620
rect 6244 568 6296 620
rect 5998 503 6050 555
rect 6080 503 6132 555
rect 6162 503 6214 555
rect 6244 503 6296 555
rect 5998 438 6050 490
rect 6080 438 6132 490
rect 6162 438 6214 490
rect 6244 438 6296 490
rect 5998 373 6050 425
rect 6080 373 6132 425
rect 6162 373 6214 425
rect 6244 373 6296 425
rect 6822 1850 6874 1902
rect 6904 1850 6956 1902
rect 6986 1850 7038 1902
rect 7068 1850 7120 1902
rect 6822 1786 6874 1838
rect 6904 1786 6956 1838
rect 6986 1786 7038 1838
rect 7068 1786 7120 1838
rect 6822 1722 6874 1774
rect 6904 1722 6956 1774
rect 6986 1722 7038 1774
rect 7068 1722 7120 1774
rect 6822 1658 6874 1710
rect 6904 1658 6956 1710
rect 6986 1658 7038 1710
rect 7068 1658 7120 1710
rect 6822 1594 6874 1646
rect 6904 1594 6956 1646
rect 6986 1594 7038 1646
rect 7068 1594 7120 1646
rect 6822 1530 6874 1582
rect 6904 1530 6956 1582
rect 6986 1530 7038 1582
rect 7068 1530 7120 1582
rect 6822 1466 6874 1518
rect 6904 1466 6956 1518
rect 6986 1466 7038 1518
rect 7068 1466 7120 1518
rect 6822 1402 6874 1454
rect 6904 1402 6956 1454
rect 6986 1402 7038 1454
rect 7068 1402 7120 1454
rect 6822 1338 6874 1390
rect 6904 1338 6956 1390
rect 6986 1338 7038 1390
rect 7068 1338 7120 1390
rect 6822 1274 6874 1326
rect 6904 1274 6956 1326
rect 6986 1274 7038 1326
rect 7068 1274 7120 1326
rect 6822 1210 6874 1262
rect 6904 1210 6956 1262
rect 6986 1210 7038 1262
rect 7068 1210 7120 1262
rect 6822 1146 6874 1198
rect 6904 1146 6956 1198
rect 6986 1146 7038 1198
rect 7068 1146 7120 1198
rect 6822 1082 6874 1134
rect 6904 1082 6956 1134
rect 6986 1082 7038 1134
rect 7068 1082 7120 1134
rect 6822 1018 6874 1070
rect 6904 1018 6956 1070
rect 6986 1018 7038 1070
rect 7068 1018 7120 1070
rect 6822 954 6874 1006
rect 6904 954 6956 1006
rect 6986 954 7038 1006
rect 7068 954 7120 1006
rect 6822 890 6874 942
rect 6904 890 6956 942
rect 6986 890 7038 942
rect 7068 890 7120 942
rect 6822 826 6874 878
rect 6904 826 6956 878
rect 6986 826 7038 878
rect 7068 826 7120 878
rect 6822 762 6874 814
rect 6904 762 6956 814
rect 6986 762 7038 814
rect 7068 762 7120 814
rect 6822 698 6874 750
rect 6904 698 6956 750
rect 6986 698 7038 750
rect 7068 698 7120 750
rect 6822 633 6874 685
rect 6904 633 6956 685
rect 6986 633 7038 685
rect 7068 633 7120 685
rect 6822 568 6874 620
rect 6904 568 6956 620
rect 6986 568 7038 620
rect 7068 568 7120 620
rect 6822 503 6874 555
rect 6904 503 6956 555
rect 6986 503 7038 555
rect 7068 503 7120 555
rect 6822 438 6874 490
rect 6904 438 6956 490
rect 6986 438 7038 490
rect 7068 438 7120 490
rect 6822 373 6874 425
rect 6904 373 6956 425
rect 6986 373 7038 425
rect 7068 373 7120 425
rect 7936 1850 7988 1902
rect 8018 1850 8070 1902
rect 8100 1850 8152 1902
rect 8182 1850 8234 1902
rect 7936 1786 7988 1838
rect 8018 1786 8070 1838
rect 8100 1786 8152 1838
rect 8182 1786 8234 1838
rect 7936 1722 7988 1774
rect 8018 1722 8070 1774
rect 8100 1722 8152 1774
rect 8182 1722 8234 1774
rect 7936 1658 7988 1710
rect 8018 1658 8070 1710
rect 8100 1658 8152 1710
rect 8182 1658 8234 1710
rect 7936 1594 7988 1646
rect 8018 1594 8070 1646
rect 8100 1594 8152 1646
rect 8182 1594 8234 1646
rect 7936 1530 7988 1582
rect 8018 1530 8070 1582
rect 8100 1530 8152 1582
rect 8182 1530 8234 1582
rect 7936 1466 7988 1518
rect 8018 1466 8070 1518
rect 8100 1466 8152 1518
rect 8182 1466 8234 1518
rect 7936 1402 7988 1454
rect 8018 1402 8070 1454
rect 8100 1402 8152 1454
rect 8182 1402 8234 1454
rect 7936 1338 7988 1390
rect 8018 1338 8070 1390
rect 8100 1338 8152 1390
rect 8182 1338 8234 1390
rect 7936 1274 7988 1326
rect 8018 1274 8070 1326
rect 8100 1274 8152 1326
rect 8182 1274 8234 1326
rect 7936 1210 7988 1262
rect 8018 1210 8070 1262
rect 8100 1210 8152 1262
rect 8182 1210 8234 1262
rect 7936 1146 7988 1198
rect 8018 1146 8070 1198
rect 8100 1146 8152 1198
rect 8182 1146 8234 1198
rect 7936 1082 7988 1134
rect 8018 1082 8070 1134
rect 8100 1082 8152 1134
rect 8182 1082 8234 1134
rect 7936 1018 7988 1070
rect 8018 1018 8070 1070
rect 8100 1018 8152 1070
rect 8182 1018 8234 1070
rect 7936 954 7988 1006
rect 8018 954 8070 1006
rect 8100 954 8152 1006
rect 8182 954 8234 1006
rect 7936 890 7988 942
rect 8018 890 8070 942
rect 8100 890 8152 942
rect 8182 890 8234 942
rect 7936 826 7988 878
rect 8018 826 8070 878
rect 8100 826 8152 878
rect 8182 826 8234 878
rect 7936 762 7988 814
rect 8018 762 8070 814
rect 8100 762 8152 814
rect 8182 762 8234 814
rect 7936 698 7988 750
rect 8018 698 8070 750
rect 8100 698 8152 750
rect 8182 698 8234 750
rect 7936 633 7988 685
rect 8018 633 8070 685
rect 8100 633 8152 685
rect 8182 633 8234 685
rect 7936 568 7988 620
rect 8018 568 8070 620
rect 8100 568 8152 620
rect 8182 568 8234 620
rect 7936 503 7988 555
rect 8018 503 8070 555
rect 8100 503 8152 555
rect 8182 503 8234 555
rect 7936 438 7988 490
rect 8018 438 8070 490
rect 8100 438 8152 490
rect 8182 438 8234 490
rect 7936 373 7988 425
rect 8018 373 8070 425
rect 8100 373 8152 425
rect 8182 373 8234 425
rect 8760 1850 8812 1902
rect 8842 1850 8894 1902
rect 8924 1850 8976 1902
rect 9006 1850 9058 1902
rect 8760 1786 8812 1838
rect 8842 1786 8894 1838
rect 8924 1786 8976 1838
rect 9006 1786 9058 1838
rect 8760 1722 8812 1774
rect 8842 1722 8894 1774
rect 8924 1722 8976 1774
rect 9006 1722 9058 1774
rect 8760 1658 8812 1710
rect 8842 1658 8894 1710
rect 8924 1658 8976 1710
rect 9006 1658 9058 1710
rect 8760 1594 8812 1646
rect 8842 1594 8894 1646
rect 8924 1594 8976 1646
rect 9006 1594 9058 1646
rect 8760 1530 8812 1582
rect 8842 1530 8894 1582
rect 8924 1530 8976 1582
rect 9006 1530 9058 1582
rect 8760 1466 8812 1518
rect 8842 1466 8894 1518
rect 8924 1466 8976 1518
rect 9006 1466 9058 1518
rect 8760 1402 8812 1454
rect 8842 1402 8894 1454
rect 8924 1402 8976 1454
rect 9006 1402 9058 1454
rect 8760 1338 8812 1390
rect 8842 1338 8894 1390
rect 8924 1338 8976 1390
rect 9006 1338 9058 1390
rect 8760 1274 8812 1326
rect 8842 1274 8894 1326
rect 8924 1274 8976 1326
rect 9006 1274 9058 1326
rect 8760 1210 8812 1262
rect 8842 1210 8894 1262
rect 8924 1210 8976 1262
rect 9006 1210 9058 1262
rect 8760 1146 8812 1198
rect 8842 1146 8894 1198
rect 8924 1146 8976 1198
rect 9006 1146 9058 1198
rect 8760 1082 8812 1134
rect 8842 1082 8894 1134
rect 8924 1082 8976 1134
rect 9006 1082 9058 1134
rect 8760 1018 8812 1070
rect 8842 1018 8894 1070
rect 8924 1018 8976 1070
rect 9006 1018 9058 1070
rect 8760 954 8812 1006
rect 8842 954 8894 1006
rect 8924 954 8976 1006
rect 9006 954 9058 1006
rect 8760 890 8812 942
rect 8842 890 8894 942
rect 8924 890 8976 942
rect 9006 890 9058 942
rect 8760 826 8812 878
rect 8842 826 8894 878
rect 8924 826 8976 878
rect 9006 826 9058 878
rect 8760 762 8812 814
rect 8842 762 8894 814
rect 8924 762 8976 814
rect 9006 762 9058 814
rect 8760 698 8812 750
rect 8842 698 8894 750
rect 8924 698 8976 750
rect 9006 698 9058 750
rect 8760 633 8812 685
rect 8842 633 8894 685
rect 8924 633 8976 685
rect 9006 633 9058 685
rect 8760 568 8812 620
rect 8842 568 8894 620
rect 8924 568 8976 620
rect 9006 568 9058 620
rect 8760 503 8812 555
rect 8842 503 8894 555
rect 8924 503 8976 555
rect 9006 503 9058 555
rect 8760 438 8812 490
rect 8842 438 8894 490
rect 8924 438 8976 490
rect 9006 438 9058 490
rect 8760 373 8812 425
rect 8842 373 8894 425
rect 8924 373 8976 425
rect 9006 373 9058 425
rect 9584 1850 9636 1902
rect 9666 1850 9718 1902
rect 9748 1850 9800 1902
rect 9830 1850 9882 1902
rect 9584 1786 9636 1838
rect 9666 1786 9718 1838
rect 9748 1786 9800 1838
rect 9830 1786 9882 1838
rect 9584 1722 9636 1774
rect 9666 1722 9718 1774
rect 9748 1722 9800 1774
rect 9830 1722 9882 1774
rect 9584 1658 9636 1710
rect 9666 1658 9718 1710
rect 9748 1658 9800 1710
rect 9830 1658 9882 1710
rect 9584 1594 9636 1646
rect 9666 1594 9718 1646
rect 9748 1594 9800 1646
rect 9830 1594 9882 1646
rect 9584 1530 9636 1582
rect 9666 1530 9718 1582
rect 9748 1530 9800 1582
rect 9830 1530 9882 1582
rect 9584 1466 9636 1518
rect 9666 1466 9718 1518
rect 9748 1466 9800 1518
rect 9830 1466 9882 1518
rect 9584 1402 9636 1454
rect 9666 1402 9718 1454
rect 9748 1402 9800 1454
rect 9830 1402 9882 1454
rect 9584 1338 9636 1390
rect 9666 1338 9718 1390
rect 9748 1338 9800 1390
rect 9830 1338 9882 1390
rect 9584 1274 9636 1326
rect 9666 1274 9718 1326
rect 9748 1274 9800 1326
rect 9830 1274 9882 1326
rect 9584 1210 9636 1262
rect 9666 1210 9718 1262
rect 9748 1210 9800 1262
rect 9830 1210 9882 1262
rect 9584 1146 9636 1198
rect 9666 1146 9718 1198
rect 9748 1146 9800 1198
rect 9830 1146 9882 1198
rect 9584 1082 9636 1134
rect 9666 1082 9718 1134
rect 9748 1082 9800 1134
rect 9830 1082 9882 1134
rect 9584 1018 9636 1070
rect 9666 1018 9718 1070
rect 9748 1018 9800 1070
rect 9830 1018 9882 1070
rect 9584 954 9636 1006
rect 9666 954 9718 1006
rect 9748 954 9800 1006
rect 9830 954 9882 1006
rect 9584 890 9636 942
rect 9666 890 9718 942
rect 9748 890 9800 942
rect 9830 890 9882 942
rect 9584 826 9636 878
rect 9666 826 9718 878
rect 9748 826 9800 878
rect 9830 826 9882 878
rect 9584 762 9636 814
rect 9666 762 9718 814
rect 9748 762 9800 814
rect 9830 762 9882 814
rect 9584 698 9636 750
rect 9666 698 9718 750
rect 9748 698 9800 750
rect 9830 698 9882 750
rect 9584 633 9636 685
rect 9666 633 9718 685
rect 9748 633 9800 685
rect 9830 633 9882 685
rect 9584 568 9636 620
rect 9666 568 9718 620
rect 9748 568 9800 620
rect 9830 568 9882 620
rect 9584 503 9636 555
rect 9666 503 9718 555
rect 9748 503 9800 555
rect 9830 503 9882 555
rect 9584 438 9636 490
rect 9666 438 9718 490
rect 9748 438 9800 490
rect 9830 438 9882 490
rect 9584 373 9636 425
rect 9666 373 9718 425
rect 9748 373 9800 425
rect 9830 373 9882 425
rect 10408 1850 10460 1902
rect 10490 1850 10542 1902
rect 10572 1850 10624 1902
rect 10654 1850 10706 1902
rect 10408 1786 10460 1838
rect 10490 1786 10542 1838
rect 10572 1786 10624 1838
rect 10654 1786 10706 1838
rect 10408 1722 10460 1774
rect 10490 1722 10542 1774
rect 10572 1722 10624 1774
rect 10654 1722 10706 1774
rect 10408 1658 10460 1710
rect 10490 1658 10542 1710
rect 10572 1658 10624 1710
rect 10654 1658 10706 1710
rect 10408 1594 10460 1646
rect 10490 1594 10542 1646
rect 10572 1594 10624 1646
rect 10654 1594 10706 1646
rect 10408 1530 10460 1582
rect 10490 1530 10542 1582
rect 10572 1530 10624 1582
rect 10654 1530 10706 1582
rect 10408 1466 10460 1518
rect 10490 1466 10542 1518
rect 10572 1466 10624 1518
rect 10654 1466 10706 1518
rect 10408 1402 10460 1454
rect 10490 1402 10542 1454
rect 10572 1402 10624 1454
rect 10654 1402 10706 1454
rect 10408 1338 10460 1390
rect 10490 1338 10542 1390
rect 10572 1338 10624 1390
rect 10654 1338 10706 1390
rect 10408 1274 10460 1326
rect 10490 1274 10542 1326
rect 10572 1274 10624 1326
rect 10654 1274 10706 1326
rect 10408 1210 10460 1262
rect 10490 1210 10542 1262
rect 10572 1210 10624 1262
rect 10654 1210 10706 1262
rect 10408 1146 10460 1198
rect 10490 1146 10542 1198
rect 10572 1146 10624 1198
rect 10654 1146 10706 1198
rect 10408 1082 10460 1134
rect 10490 1082 10542 1134
rect 10572 1082 10624 1134
rect 10654 1082 10706 1134
rect 10408 1018 10460 1070
rect 10490 1018 10542 1070
rect 10572 1018 10624 1070
rect 10654 1018 10706 1070
rect 10408 954 10460 1006
rect 10490 954 10542 1006
rect 10572 954 10624 1006
rect 10654 954 10706 1006
rect 10408 890 10460 942
rect 10490 890 10542 942
rect 10572 890 10624 942
rect 10654 890 10706 942
rect 10408 826 10460 878
rect 10490 826 10542 878
rect 10572 826 10624 878
rect 10654 826 10706 878
rect 10408 762 10460 814
rect 10490 762 10542 814
rect 10572 762 10624 814
rect 10654 762 10706 814
rect 10408 698 10460 750
rect 10490 698 10542 750
rect 10572 698 10624 750
rect 10654 698 10706 750
rect 10408 633 10460 685
rect 10490 633 10542 685
rect 10572 633 10624 685
rect 10654 633 10706 685
rect 10408 568 10460 620
rect 10490 568 10542 620
rect 10572 568 10624 620
rect 10654 568 10706 620
rect 10408 503 10460 555
rect 10490 503 10542 555
rect 10572 503 10624 555
rect 10654 503 10706 555
rect 10408 438 10460 490
rect 10490 438 10542 490
rect 10572 438 10624 490
rect 10654 438 10706 490
rect 10408 373 10460 425
rect 10490 373 10542 425
rect 10572 373 10624 425
rect 10654 373 10706 425
rect 4191 304 4243 356
rect 4259 304 4311 356
rect 4327 304 4379 356
rect 4395 304 4447 356
rect 4463 304 4515 356
rect 4531 304 4583 356
rect 4599 304 4651 356
rect 4666 304 4718 356
rect 4733 304 4785 356
rect 4800 304 4852 356
rect 4867 304 4919 356
rect 4934 304 4986 356
rect 5001 304 5053 356
rect 5068 304 5120 356
rect 5149 305 5201 357
rect 5221 305 5273 357
rect 5293 305 5345 357
rect 5365 305 5417 357
rect 5436 305 5488 357
rect 5507 305 5559 357
rect 5578 305 5630 357
rect 5659 304 5711 356
rect 5724 304 5776 356
rect 5789 304 5841 356
rect 5854 304 5906 356
rect 5919 304 5971 356
rect 5984 304 6036 356
rect 6049 304 6101 356
rect 6114 304 6166 356
rect 6179 304 6231 356
rect 6244 304 6296 356
rect 6309 304 6361 356
rect 6374 304 6426 356
rect 6439 304 6491 356
rect 6504 304 6556 356
rect 6569 304 6621 356
rect 6634 304 6686 356
rect 6699 304 6751 356
rect 6764 304 6816 356
rect 6829 304 6881 356
rect 6894 304 6946 356
rect 6959 304 7011 356
rect 7024 304 7076 356
rect 7089 304 7141 356
rect 7154 304 7206 356
rect 7219 304 7271 356
rect 7284 304 7336 356
rect 7349 304 7401 356
rect 7414 304 7466 356
rect 7479 304 7531 356
rect 7544 304 7596 356
rect 7609 304 7661 356
rect 7674 304 7726 356
rect 7739 304 7791 356
rect 7804 304 7856 356
rect 7869 304 7921 356
rect 7934 304 7986 356
rect 7999 304 8051 356
rect 8064 304 8116 356
rect 8129 304 8181 356
rect 8194 304 8246 356
rect 8259 304 8311 356
rect 8324 304 8376 356
rect 8389 304 8441 356
rect 8454 304 8506 356
rect 8519 304 8571 356
rect 8584 304 8636 356
rect 8649 304 8701 356
rect 8714 304 8766 356
rect 8779 304 8831 356
rect 8844 304 8896 356
rect 8909 304 8961 356
rect 8974 304 9026 356
rect 9039 304 9091 356
rect 9104 304 9156 356
rect 9169 304 9221 356
rect 9234 304 9286 356
rect 9299 304 9351 356
rect 9364 304 9416 356
rect 9429 304 9481 356
rect 9494 304 9546 356
rect 9559 304 9611 356
rect 9624 304 9676 356
rect 9689 304 9741 356
rect 9753 304 9805 356
rect 9817 304 9869 356
rect 9881 304 9933 356
rect 9945 304 9997 356
rect 10009 304 10061 356
rect 10073 304 10125 356
rect 10137 304 10189 356
rect 10201 304 10253 356
rect 10265 304 10317 356
rect 10329 304 10381 356
rect 10393 304 10445 356
rect 10457 304 10509 356
rect 10521 304 10573 356
rect 10585 304 10637 356
rect 10649 304 10701 356
rect 4191 230 4243 282
rect 4259 230 4311 282
rect 4327 230 4379 282
rect 4395 230 4447 282
rect 4463 230 4515 282
rect 4531 230 4583 282
rect 4599 230 4651 282
rect 4666 230 4718 282
rect 4733 230 4785 282
rect 4800 230 4852 282
rect 4867 230 4919 282
rect 4934 230 4986 282
rect 5001 230 5053 282
rect 5068 230 5120 282
rect 5149 225 5201 277
rect 5221 225 5273 277
rect 5293 225 5345 277
rect 5365 225 5417 277
rect 5436 225 5488 277
rect 5507 225 5559 277
rect 5578 225 5630 277
rect 5659 230 5711 282
rect 5724 230 5776 282
rect 5789 230 5841 282
rect 5854 230 5906 282
rect 5919 230 5971 282
rect 5984 230 6036 282
rect 6049 230 6101 282
rect 6114 230 6166 282
rect 6179 230 6231 282
rect 6244 230 6296 282
rect 6309 230 6361 282
rect 6374 230 6426 282
rect 6439 230 6491 282
rect 6504 230 6556 282
rect 6569 230 6621 282
rect 6634 230 6686 282
rect 6699 230 6751 282
rect 6764 230 6816 282
rect 6829 230 6881 282
rect 6894 230 6946 282
rect 6959 230 7011 282
rect 7024 230 7076 282
rect 7089 230 7141 282
rect 7154 230 7206 282
rect 7219 230 7271 282
rect 7284 230 7336 282
rect 7349 230 7401 282
rect 7414 230 7466 282
rect 7479 230 7531 282
rect 7544 230 7596 282
rect 7609 230 7661 282
rect 7674 230 7726 282
rect 7739 230 7791 282
rect 7804 230 7856 282
rect 7869 230 7921 282
rect 7934 230 7986 282
rect 7999 230 8051 282
rect 8064 230 8116 282
rect 8129 230 8181 282
rect 8194 230 8246 282
rect 8259 230 8311 282
rect 8324 230 8376 282
rect 8389 230 8441 282
rect 8454 230 8506 282
rect 8519 230 8571 282
rect 8584 230 8636 282
rect 8649 230 8701 282
rect 8714 230 8766 282
rect 8779 230 8831 282
rect 8844 230 8896 282
rect 8909 230 8961 282
rect 8974 230 9026 282
rect 9039 230 9091 282
rect 9104 230 9156 282
rect 9169 230 9221 282
rect 9234 230 9286 282
rect 9299 230 9351 282
rect 9364 230 9416 282
rect 9429 230 9481 282
rect 9494 230 9546 282
rect 9559 230 9611 282
rect 9624 230 9676 282
rect 9689 230 9741 282
rect 9753 230 9805 282
rect 9817 230 9869 282
rect 9881 230 9933 282
rect 9945 230 9997 282
rect 10009 230 10061 282
rect 10073 230 10125 282
rect 10137 230 10189 282
rect 10201 230 10253 282
rect 10265 230 10317 282
rect 10329 230 10381 282
rect 10393 230 10445 282
rect 10457 230 10509 282
rect 10521 230 10573 282
rect 10585 230 10637 282
rect 10649 230 10701 282
rect 4191 156 4243 208
rect 4259 156 4311 208
rect 4327 156 4379 208
rect 4395 156 4447 208
rect 4463 156 4515 208
rect 4531 156 4583 208
rect 4599 156 4651 208
rect 4666 156 4718 208
rect 4733 156 4785 208
rect 4800 156 4852 208
rect 4867 156 4919 208
rect 4934 156 4986 208
rect 5001 156 5053 208
rect 5068 156 5120 208
rect 5149 145 5201 197
rect 5221 145 5273 197
rect 5293 145 5345 197
rect 5365 145 5417 197
rect 5436 145 5488 197
rect 5507 145 5559 197
rect 5578 145 5630 197
rect 5659 156 5711 208
rect 5724 156 5776 208
rect 5789 156 5841 208
rect 5854 156 5906 208
rect 5919 156 5971 208
rect 5984 156 6036 208
rect 6049 156 6101 208
rect 6114 156 6166 208
rect 6179 156 6231 208
rect 6244 156 6296 208
rect 6309 156 6361 208
rect 6374 156 6426 208
rect 6439 156 6491 208
rect 6504 156 6556 208
rect 6569 156 6621 208
rect 6634 156 6686 208
rect 6699 156 6751 208
rect 6764 156 6816 208
rect 6829 156 6881 208
rect 6894 156 6946 208
rect 6959 156 7011 208
rect 7024 156 7076 208
rect 7089 156 7141 208
rect 7154 156 7206 208
rect 7219 156 7271 208
rect 7284 156 7336 208
rect 7349 156 7401 208
rect 7414 156 7466 208
rect 7479 156 7531 208
rect 7544 156 7596 208
rect 7609 156 7661 208
rect 7674 156 7726 208
rect 7739 156 7791 208
rect 7804 156 7856 208
rect 7869 156 7921 208
rect 7934 156 7986 208
rect 7999 156 8051 208
rect 8064 156 8116 208
rect 8129 156 8181 208
rect 8194 156 8246 208
rect 8259 156 8311 208
rect 8324 156 8376 208
rect 8389 156 8441 208
rect 8454 156 8506 208
rect 8519 156 8571 208
rect 8584 156 8636 208
rect 8649 156 8701 208
rect 8714 156 8766 208
rect 8779 156 8831 208
rect 8844 156 8896 208
rect 8909 156 8961 208
rect 8974 156 9026 208
rect 9039 156 9091 208
rect 9104 156 9156 208
rect 9169 156 9221 208
rect 9234 156 9286 208
rect 9299 156 9351 208
rect 9364 156 9416 208
rect 9429 156 9481 208
rect 9494 156 9546 208
rect 9559 156 9611 208
rect 9624 156 9676 208
rect 9689 156 9741 208
rect 9753 156 9805 208
rect 9817 156 9869 208
rect 9881 156 9933 208
rect 9945 156 9997 208
rect 10009 156 10061 208
rect 10073 156 10125 208
rect 10137 156 10189 208
rect 10201 156 10253 208
rect 10265 156 10317 208
rect 10329 156 10381 208
rect 10393 156 10445 208
rect 10457 156 10509 208
rect 10521 156 10573 208
rect 10585 156 10637 208
rect 10649 156 10701 208
rect 4191 82 4243 134
rect 4259 82 4311 134
rect 4327 82 4379 134
rect 4395 82 4447 134
rect 4463 82 4515 134
rect 4531 82 4583 134
rect 4599 82 4651 134
rect 4666 82 4718 134
rect 4733 82 4785 134
rect 4800 82 4852 134
rect 4867 82 4919 134
rect 4934 82 4986 134
rect 5001 82 5053 134
rect 5068 82 5120 134
rect 5149 65 5201 117
rect 5221 65 5273 117
rect 5293 65 5345 117
rect 5365 65 5417 117
rect 5436 65 5488 117
rect 5507 65 5559 117
rect 5578 65 5630 117
rect 5659 82 5711 134
rect 5724 82 5776 134
rect 5789 82 5841 134
rect 5854 82 5906 134
rect 5919 82 5971 134
rect 5984 82 6036 134
rect 6049 82 6101 134
rect 6114 82 6166 134
rect 6179 82 6231 134
rect 6244 82 6296 134
rect 6309 82 6361 134
rect 6374 82 6426 134
rect 6439 82 6491 134
rect 6504 82 6556 134
rect 6569 82 6621 134
rect 6634 82 6686 134
rect 6699 82 6751 134
rect 6764 82 6816 134
rect 6829 82 6881 134
rect 6894 82 6946 134
rect 6959 82 7011 134
rect 7024 82 7076 134
rect 7089 82 7141 134
rect 7154 82 7206 134
rect 7219 82 7271 134
rect 7284 82 7336 134
rect 7349 82 7401 134
rect 7414 82 7466 134
rect 7479 82 7531 134
rect 7544 82 7596 134
rect 7609 82 7661 134
rect 7674 82 7726 134
rect 7739 82 7791 134
rect 7804 82 7856 134
rect 7869 82 7921 134
rect 7934 82 7986 134
rect 7999 82 8051 134
rect 8064 82 8116 134
rect 8129 82 8181 134
rect 8194 82 8246 134
rect 8259 82 8311 134
rect 8324 82 8376 134
rect 8389 82 8441 134
rect 8454 82 8506 134
rect 8519 82 8571 134
rect 8584 82 8636 134
rect 8649 82 8701 134
rect 8714 82 8766 134
rect 8779 82 8831 134
rect 8844 82 8896 134
rect 8909 82 8961 134
rect 8974 82 9026 134
rect 9039 82 9091 134
rect 9104 82 9156 134
rect 9169 82 9221 134
rect 9234 82 9286 134
rect 9299 82 9351 134
rect 9364 82 9416 134
rect 9429 82 9481 134
rect 9494 82 9546 134
rect 9559 82 9611 134
rect 9624 82 9676 134
rect 9689 82 9741 134
rect 9753 82 9805 134
rect 9817 82 9869 134
rect 9881 82 9933 134
rect 9945 82 9997 134
rect 10009 82 10061 134
rect 10073 82 10125 134
rect 10137 82 10189 134
rect 10201 82 10253 134
rect 10265 82 10317 134
rect 10329 82 10381 134
rect 10393 82 10445 134
rect 10457 82 10509 134
rect 10521 82 10573 134
rect 10585 82 10637 134
rect 10649 82 10701 134
rect 4191 8 4243 60
rect 4259 8 4311 60
rect 4327 8 4379 60
rect 4395 8 4447 60
rect 4463 8 4515 60
rect 4531 8 4583 60
rect 4599 8 4651 60
rect 4666 8 4718 60
rect 4733 8 4785 60
rect 4800 8 4852 60
rect 4867 8 4919 60
rect 4934 8 4986 60
rect 5001 8 5053 60
rect 5068 8 5120 60
rect 5659 8 5711 60
rect 5724 8 5776 60
rect 5789 8 5841 60
rect 5854 8 5906 60
rect 5919 8 5971 60
rect 5984 8 6036 60
rect 6049 8 6101 60
rect 6114 8 6166 60
rect 6179 8 6231 60
rect 6244 8 6296 60
rect 6309 8 6361 60
rect 6374 8 6426 60
rect 6439 8 6491 60
rect 6504 8 6556 60
rect 6569 8 6621 60
rect 6634 8 6686 60
rect 6699 8 6751 60
rect 6764 8 6816 60
rect 6829 8 6881 60
rect 6894 8 6946 60
rect 6959 8 7011 60
rect 7024 8 7076 60
rect 7089 8 7141 60
rect 7154 8 7206 60
rect 7219 8 7271 60
rect 7284 8 7336 60
rect 7349 8 7401 60
rect 7414 8 7466 60
rect 7479 8 7531 60
rect 7544 8 7596 60
rect 7609 8 7661 60
rect 7674 8 7726 60
rect 7739 8 7791 60
rect 7804 8 7856 60
rect 7869 8 7921 60
rect 7934 8 7986 60
rect 7999 8 8051 60
rect 8064 8 8116 60
rect 8129 8 8181 60
rect 8194 8 8246 60
rect 8259 8 8311 60
rect 8324 8 8376 60
rect 8389 8 8441 60
rect 8454 8 8506 60
rect 8519 8 8571 60
rect 8584 8 8636 60
rect 8649 8 8701 60
rect 8714 8 8766 60
rect 8779 8 8831 60
rect 8844 8 8896 60
rect 8909 8 8961 60
rect 8974 8 9026 60
rect 9039 8 9091 60
rect 9104 8 9156 60
rect 9169 8 9221 60
rect 9234 8 9286 60
rect 9299 8 9351 60
rect 9364 8 9416 60
rect 9429 8 9481 60
rect 9494 8 9546 60
rect 9559 8 9611 60
rect 9624 8 9676 60
rect 9689 8 9741 60
rect 9753 8 9805 60
rect 9817 8 9869 60
rect 9881 8 9933 60
rect 9945 8 9997 60
rect 10009 8 10061 60
rect 10073 8 10125 60
rect 10137 8 10189 60
rect 10201 8 10253 60
rect 10265 8 10317 60
rect 10329 8 10381 60
rect 10393 8 10445 60
rect 10457 8 10509 60
rect 10521 8 10573 60
rect 10585 8 10637 60
rect 10649 8 10701 60
<< metal2 >>
rect 2872 38834 2878 38886
rect 2930 38834 2943 38886
rect 2995 38834 3008 38886
rect 3060 38834 3073 38886
rect 3125 38834 3138 38886
rect 3190 38834 3203 38886
rect 3255 38834 3268 38886
rect 3320 38834 3332 38886
rect 3384 38834 3396 38886
rect 3448 38834 3460 38886
rect 3512 38834 3524 38886
rect 3576 38834 3588 38886
rect 3640 38834 3652 38886
rect 3704 38834 3716 38886
rect 3768 38834 3780 38886
rect 3832 38834 3844 38886
rect 3896 38834 3908 38886
rect 3960 38834 3972 38886
rect 4024 38834 4036 38886
rect 4088 38834 4100 38886
rect 4152 38834 4164 38886
rect 4216 38834 4228 38886
rect 4280 38834 4292 38886
rect 4344 38834 4356 38886
rect 4408 38834 4420 38886
rect 4472 38834 4484 38886
rect 4536 38834 4548 38886
rect 4600 38834 4612 38886
rect 4664 38834 4676 38886
rect 4728 38834 4740 38886
rect 4792 38834 4804 38886
rect 4856 38834 4868 38886
rect 4920 38834 4932 38886
rect 4984 38834 4996 38886
rect 5048 38834 5060 38886
rect 5112 38834 5124 38886
rect 5176 38834 5188 38886
rect 5240 38834 5252 38886
rect 5304 38834 5316 38886
rect 5368 38834 5380 38886
rect 5432 38834 5444 38886
rect 5496 38834 5508 38886
rect 5560 38834 5572 38886
rect 5624 38834 5636 38886
rect 5688 38834 5700 38886
rect 5752 38834 5764 38886
rect 5816 38834 5828 38886
rect 5880 38834 5892 38886
rect 5944 38834 5956 38886
rect 6008 38834 6020 38886
rect 6072 38834 6084 38886
rect 6136 38834 6148 38886
rect 6200 38834 6212 38886
rect 6264 38834 6276 38886
rect 6328 38834 6340 38886
rect 6392 38834 6404 38886
rect 6456 38834 6468 38886
rect 6520 38834 6532 38886
rect 6584 38834 6596 38886
rect 6648 38834 6660 38886
rect 6712 38834 6724 38886
rect 6776 38834 6788 38886
rect 6840 38834 6852 38886
rect 6904 38834 6916 38886
rect 6968 38834 6980 38886
rect 7032 38834 7044 38886
rect 7096 38834 7108 38886
rect 7160 38834 7172 38886
rect 7224 38834 7236 38886
rect 7288 38834 7300 38886
rect 7352 38834 7364 38886
rect 7416 38834 7428 38886
rect 7480 38834 7492 38886
rect 7544 38834 7556 38886
rect 7608 38834 7620 38886
rect 7672 38834 7684 38886
rect 7736 38834 7748 38886
rect 7800 38834 7812 38886
rect 7864 38834 7876 38886
rect 7928 38834 7940 38886
rect 7992 38834 8004 38886
rect 8056 38834 8068 38886
rect 8120 38834 8132 38886
rect 8184 38834 8196 38886
rect 8248 38834 8260 38886
rect 8312 38834 8324 38886
rect 8376 38834 8388 38886
rect 8440 38834 8452 38886
rect 8504 38834 8516 38886
rect 8568 38834 8580 38886
rect 8632 38834 8644 38886
rect 8696 38834 8708 38886
rect 8760 38834 8772 38886
rect 8824 38834 8836 38886
rect 8888 38834 8900 38886
rect 8952 38834 8964 38886
rect 9016 38834 9028 38886
rect 9080 38834 9092 38886
rect 9144 38834 9156 38886
rect 9208 38834 9220 38886
rect 9272 38834 9284 38886
rect 9336 38834 9348 38886
rect 9400 38834 9412 38886
rect 9464 38834 9476 38886
rect 9528 38834 9540 38886
rect 9592 38834 9604 38886
rect 9656 38834 9668 38886
rect 9720 38834 9732 38886
rect 9784 38834 9796 38886
rect 9848 38834 9860 38886
rect 9912 38834 9924 38886
rect 9976 38834 9988 38886
rect 10040 38834 10052 38886
rect 10104 38834 10116 38886
rect 10168 38834 10180 38886
rect 10232 38834 10244 38886
rect 10296 38834 10308 38886
rect 10360 38834 10372 38886
rect 10424 38834 10436 38886
rect 10488 38834 10500 38886
rect 10552 38834 10564 38886
rect 10616 38834 10628 38886
rect 10680 38834 10692 38886
rect 10744 38834 10756 38886
rect 10808 38834 10820 38886
rect 10872 38834 10884 38886
rect 10936 38834 10948 38886
rect 11000 38834 11012 38886
rect 11064 38834 11076 38886
rect 11128 38834 11140 38886
rect 11192 38834 11204 38886
rect 11256 38834 11268 38886
rect 11320 38834 11332 38886
rect 11384 38834 11396 38886
rect 11448 38834 11460 38886
rect 11512 38834 11524 38886
rect 11576 38834 11588 38886
rect 11640 38834 11652 38886
rect 11704 38834 11716 38886
rect 11768 38834 11780 38886
rect 11832 38834 11844 38886
rect 11896 38834 11908 38886
rect 11960 38834 11972 38886
rect 12024 38834 12036 38886
rect 12088 38834 12100 38886
rect 12152 38834 12164 38886
rect 12216 38834 12228 38886
rect 12280 38834 12292 38886
rect 12344 38834 12356 38886
rect 12408 38834 12420 38886
rect 12472 38834 12484 38886
rect 12536 38834 12548 38886
rect 12600 38834 12612 38886
rect 12664 38834 12676 38886
rect 12728 38834 12740 38886
rect 12792 38834 12804 38886
rect 12856 38834 12868 38886
rect 12920 38834 12932 38886
rect 12984 38834 12996 38886
rect 13048 38834 13060 38886
rect 13112 38834 13118 38886
rect 100 38720 13602 38726
rect 100 38668 2249 38720
rect 2301 38668 2315 38720
rect 2367 38668 2673 38720
rect 2725 38668 2739 38720
rect 2791 38668 3227 38720
rect 3279 38668 3293 38720
rect 3345 38668 3781 38720
rect 3833 38668 3847 38720
rect 3899 38668 4335 38720
rect 4387 38668 4401 38720
rect 4453 38668 4889 38720
rect 4941 38668 4955 38720
rect 5007 38668 5443 38720
rect 5495 38668 5509 38720
rect 5561 38668 5997 38720
rect 6049 38668 6063 38720
rect 6115 38668 6551 38720
rect 6603 38668 6617 38720
rect 6669 38668 7105 38720
rect 7157 38668 7171 38720
rect 7223 38668 7659 38720
rect 7711 38668 7725 38720
rect 7777 38668 8213 38720
rect 8265 38668 8279 38720
rect 8331 38668 8767 38720
rect 8819 38668 8833 38720
rect 8885 38668 9321 38720
rect 9373 38668 9387 38720
rect 9439 38668 9875 38720
rect 9927 38668 9941 38720
rect 9993 38668 10429 38720
rect 10481 38668 10495 38720
rect 10547 38668 10983 38720
rect 11035 38668 11049 38720
rect 11101 38668 11537 38720
rect 11589 38668 11603 38720
rect 11655 38668 12091 38720
rect 12143 38668 12157 38720
rect 12209 38668 12645 38720
rect 12697 38668 12711 38720
rect 12763 38668 13200 38720
rect 13252 38668 13270 38720
rect 13322 38668 13340 38720
rect 13392 38668 13410 38720
rect 13462 38668 13480 38720
rect 13532 38668 13550 38720
rect 100 38656 13602 38668
rect 100 38604 2249 38656
rect 2301 38604 2315 38656
rect 2367 38604 2673 38656
rect 2725 38604 2739 38656
rect 2791 38654 13602 38656
rect 2791 38604 3227 38654
rect 100 38602 3227 38604
rect 3279 38602 3293 38654
rect 3345 38602 3781 38654
rect 3833 38602 3847 38654
rect 3899 38602 4335 38654
rect 4387 38602 4401 38654
rect 4453 38602 4889 38654
rect 4941 38602 4955 38654
rect 5007 38602 5443 38654
rect 5495 38602 5509 38654
rect 5561 38602 5997 38654
rect 6049 38602 6063 38654
rect 6115 38602 6551 38654
rect 6603 38602 6617 38654
rect 6669 38602 7105 38654
rect 7157 38602 7171 38654
rect 7223 38602 7659 38654
rect 7711 38602 7725 38654
rect 7777 38602 8213 38654
rect 8265 38602 8279 38654
rect 8331 38602 8767 38654
rect 8819 38602 8833 38654
rect 8885 38602 9321 38654
rect 9373 38602 9387 38654
rect 9439 38602 9875 38654
rect 9927 38602 9941 38654
rect 9993 38602 10429 38654
rect 10481 38602 10495 38654
rect 10547 38602 10983 38654
rect 11035 38602 11049 38654
rect 11101 38602 11537 38654
rect 11589 38602 11603 38654
rect 11655 38602 12091 38654
rect 12143 38602 12157 38654
rect 12209 38602 12645 38654
rect 12697 38602 12711 38654
rect 12763 38602 13200 38654
rect 13252 38602 13270 38654
rect 13322 38602 13340 38654
rect 13392 38602 13410 38654
rect 13462 38602 13480 38654
rect 13532 38602 13550 38654
rect 100 38592 13602 38602
rect 100 38540 2249 38592
rect 2301 38540 2315 38592
rect 2367 38540 2673 38592
rect 2725 38540 2739 38592
rect 2791 38588 13602 38592
rect 2791 38540 3227 38588
rect 100 38536 3227 38540
rect 3279 38536 3293 38588
rect 3345 38536 3781 38588
rect 3833 38536 3847 38588
rect 3899 38536 4335 38588
rect 4387 38536 4401 38588
rect 4453 38536 4889 38588
rect 4941 38536 4955 38588
rect 5007 38536 5443 38588
rect 5495 38536 5509 38588
rect 5561 38536 5997 38588
rect 6049 38536 6063 38588
rect 6115 38536 6551 38588
rect 6603 38536 6617 38588
rect 6669 38536 7105 38588
rect 7157 38536 7171 38588
rect 7223 38536 7659 38588
rect 7711 38536 7725 38588
rect 7777 38536 8213 38588
rect 8265 38536 8279 38588
rect 8331 38536 8767 38588
rect 8819 38536 8833 38588
rect 8885 38536 9321 38588
rect 9373 38536 9387 38588
rect 9439 38536 9875 38588
rect 9927 38536 9941 38588
rect 9993 38536 10429 38588
rect 10481 38536 10495 38588
rect 10547 38536 10983 38588
rect 11035 38536 11049 38588
rect 11101 38536 11537 38588
rect 11589 38536 11603 38588
rect 11655 38536 12091 38588
rect 12143 38536 12157 38588
rect 12209 38536 12645 38588
rect 12697 38536 12711 38588
rect 12763 38536 13200 38588
rect 13252 38536 13270 38588
rect 13322 38536 13340 38588
rect 13392 38536 13410 38588
rect 13462 38536 13480 38588
rect 13532 38536 13550 38588
rect 100 38528 13602 38536
rect 100 38476 2249 38528
rect 2301 38476 2315 38528
rect 2367 38476 2673 38528
rect 2725 38476 2739 38528
rect 2791 38522 13602 38528
rect 2791 38476 3227 38522
rect 100 38470 3227 38476
rect 3279 38470 3293 38522
rect 3345 38470 3781 38522
rect 3833 38470 3847 38522
rect 3899 38470 4335 38522
rect 4387 38470 4401 38522
rect 4453 38470 4889 38522
rect 4941 38470 4955 38522
rect 5007 38470 5443 38522
rect 5495 38470 5509 38522
rect 5561 38470 5997 38522
rect 6049 38470 6063 38522
rect 6115 38470 6551 38522
rect 6603 38470 6617 38522
rect 6669 38470 7105 38522
rect 7157 38470 7171 38522
rect 7223 38470 7659 38522
rect 7711 38470 7725 38522
rect 7777 38470 8213 38522
rect 8265 38470 8279 38522
rect 8331 38470 8767 38522
rect 8819 38470 8833 38522
rect 8885 38470 9321 38522
rect 9373 38470 9387 38522
rect 9439 38470 9875 38522
rect 9927 38470 9941 38522
rect 9993 38470 10429 38522
rect 10481 38470 10495 38522
rect 10547 38470 10983 38522
rect 11035 38470 11049 38522
rect 11101 38470 11537 38522
rect 11589 38470 11603 38522
rect 11655 38470 12091 38522
rect 12143 38470 12157 38522
rect 12209 38470 12645 38522
rect 12697 38470 12711 38522
rect 12763 38470 13200 38522
rect 13252 38470 13270 38522
rect 13322 38470 13340 38522
rect 13392 38470 13410 38522
rect 13462 38470 13480 38522
rect 13532 38470 13550 38522
rect 100 38464 13602 38470
rect 100 38412 2249 38464
rect 2301 38412 2315 38464
rect 2367 38412 2673 38464
rect 2725 38412 2739 38464
rect 2791 38456 13602 38464
rect 2791 38412 3227 38456
rect 100 38404 3227 38412
rect 3279 38404 3293 38456
rect 3345 38404 3781 38456
rect 3833 38404 3847 38456
rect 3899 38404 4335 38456
rect 4387 38404 4401 38456
rect 4453 38404 4889 38456
rect 4941 38404 4955 38456
rect 5007 38404 5443 38456
rect 5495 38404 5509 38456
rect 5561 38404 5997 38456
rect 6049 38404 6063 38456
rect 6115 38404 6551 38456
rect 6603 38404 6617 38456
rect 6669 38404 7105 38456
rect 7157 38404 7171 38456
rect 7223 38404 7659 38456
rect 7711 38404 7725 38456
rect 7777 38404 8213 38456
rect 8265 38404 8279 38456
rect 8331 38404 8767 38456
rect 8819 38404 8833 38456
rect 8885 38404 9321 38456
rect 9373 38404 9387 38456
rect 9439 38404 9875 38456
rect 9927 38404 9941 38456
rect 9993 38404 10429 38456
rect 10481 38404 10495 38456
rect 10547 38404 10983 38456
rect 11035 38404 11049 38456
rect 11101 38404 11537 38456
rect 11589 38404 11603 38456
rect 11655 38404 12091 38456
rect 12143 38404 12157 38456
rect 12209 38404 12645 38456
rect 12697 38404 12711 38456
rect 12763 38404 13200 38456
rect 13252 38404 13270 38456
rect 13322 38404 13340 38456
rect 13392 38404 13410 38456
rect 13462 38404 13480 38456
rect 13532 38404 13550 38456
rect 100 38400 13602 38404
rect 100 38348 2249 38400
rect 2301 38348 2315 38400
rect 2367 38348 2673 38400
rect 2725 38348 2739 38400
rect 2791 38390 13602 38400
rect 2791 38348 3227 38390
rect 100 38338 3227 38348
rect 3279 38338 3293 38390
rect 3345 38338 3781 38390
rect 3833 38338 3847 38390
rect 3899 38338 4335 38390
rect 4387 38338 4401 38390
rect 4453 38338 4889 38390
rect 4941 38338 4955 38390
rect 5007 38338 5443 38390
rect 5495 38338 5509 38390
rect 5561 38338 5997 38390
rect 6049 38338 6063 38390
rect 6115 38338 6551 38390
rect 6603 38338 6617 38390
rect 6669 38338 7105 38390
rect 7157 38338 7171 38390
rect 7223 38338 7659 38390
rect 7711 38338 7725 38390
rect 7777 38338 8213 38390
rect 8265 38338 8279 38390
rect 8331 38338 8767 38390
rect 8819 38338 8833 38390
rect 8885 38338 9321 38390
rect 9373 38338 9387 38390
rect 9439 38338 9875 38390
rect 9927 38338 9941 38390
rect 9993 38338 10429 38390
rect 10481 38338 10495 38390
rect 10547 38338 10983 38390
rect 11035 38338 11049 38390
rect 11101 38338 11537 38390
rect 11589 38338 11603 38390
rect 11655 38338 12091 38390
rect 12143 38338 12157 38390
rect 12209 38338 12645 38390
rect 12697 38338 12711 38390
rect 12763 38338 13200 38390
rect 13252 38338 13270 38390
rect 13322 38338 13340 38390
rect 13392 38338 13410 38390
rect 13462 38338 13480 38390
rect 13532 38338 13550 38390
rect 100 38336 13602 38338
rect 100 38284 2249 38336
rect 2301 38284 2315 38336
rect 2367 38284 2673 38336
rect 2725 38284 2739 38336
rect 2791 38323 13602 38336
rect 2791 38284 3227 38323
rect 100 38272 3227 38284
rect 100 38220 2249 38272
rect 2301 38220 2315 38272
rect 2367 38271 3227 38272
rect 3279 38271 3293 38323
rect 3345 38271 3781 38323
rect 3833 38271 3847 38323
rect 3899 38271 4335 38323
rect 4387 38271 4401 38323
rect 4453 38271 4889 38323
rect 4941 38271 4955 38323
rect 5007 38271 5443 38323
rect 5495 38271 5509 38323
rect 5561 38271 5997 38323
rect 6049 38271 6063 38323
rect 6115 38271 6551 38323
rect 6603 38271 6617 38323
rect 6669 38271 7105 38323
rect 7157 38271 7171 38323
rect 7223 38271 7659 38323
rect 7711 38271 7725 38323
rect 7777 38271 8213 38323
rect 8265 38271 8279 38323
rect 8331 38271 8767 38323
rect 8819 38271 8833 38323
rect 8885 38271 9321 38323
rect 9373 38271 9387 38323
rect 9439 38271 9875 38323
rect 9927 38271 9941 38323
rect 9993 38271 10429 38323
rect 10481 38271 10495 38323
rect 10547 38271 10983 38323
rect 11035 38271 11049 38323
rect 11101 38271 11537 38323
rect 11589 38271 11603 38323
rect 11655 38271 12091 38323
rect 12143 38271 12157 38323
rect 12209 38271 12645 38323
rect 12697 38271 12711 38323
rect 12763 38271 13200 38323
rect 13252 38271 13270 38323
rect 13322 38271 13340 38323
rect 13392 38271 13410 38323
rect 13462 38271 13480 38323
rect 13532 38271 13550 38323
rect 2367 38220 2673 38271
rect 100 38219 2673 38220
rect 2725 38219 2739 38271
rect 2791 38256 13602 38271
rect 2791 38219 3227 38256
rect 100 38208 3227 38219
rect 100 38156 2249 38208
rect 2301 38156 2315 38208
rect 2367 38206 3227 38208
rect 2367 38156 2673 38206
rect 100 38154 2673 38156
rect 2725 38154 2739 38206
rect 2791 38204 3227 38206
rect 3279 38204 3293 38256
rect 3345 38204 3781 38256
rect 3833 38204 3847 38256
rect 3899 38204 4335 38256
rect 4387 38204 4401 38256
rect 4453 38204 4889 38256
rect 4941 38204 4955 38256
rect 5007 38204 5443 38256
rect 5495 38204 5509 38256
rect 5561 38204 5997 38256
rect 6049 38204 6063 38256
rect 6115 38204 6551 38256
rect 6603 38204 6617 38256
rect 6669 38204 7105 38256
rect 7157 38204 7171 38256
rect 7223 38204 7659 38256
rect 7711 38204 7725 38256
rect 7777 38204 8213 38256
rect 8265 38204 8279 38256
rect 8331 38204 8767 38256
rect 8819 38204 8833 38256
rect 8885 38204 9321 38256
rect 9373 38204 9387 38256
rect 9439 38204 9875 38256
rect 9927 38204 9941 38256
rect 9993 38204 10429 38256
rect 10481 38204 10495 38256
rect 10547 38204 10983 38256
rect 11035 38204 11049 38256
rect 11101 38204 11537 38256
rect 11589 38204 11603 38256
rect 11655 38204 12091 38256
rect 12143 38204 12157 38256
rect 12209 38204 12645 38256
rect 12697 38204 12711 38256
rect 12763 38204 13200 38256
rect 13252 38204 13270 38256
rect 13322 38204 13340 38256
rect 13392 38204 13410 38256
rect 13462 38204 13480 38256
rect 13532 38204 13550 38256
rect 2791 38198 13602 38204
rect 2791 38154 2792 38198
rect 100 38144 2792 38154
rect 100 38092 2249 38144
rect 2301 38092 2315 38144
rect 2367 38141 2792 38144
rect 2367 38092 2673 38141
rect 100 38089 2673 38092
rect 2725 38089 2739 38141
rect 2791 38089 2792 38141
rect 100 38080 2792 38089
rect 100 38028 2249 38080
rect 2301 38028 2315 38080
rect 2367 38076 2792 38080
rect 2367 38028 2673 38076
rect 100 38024 2673 38028
rect 2725 38024 2739 38076
rect 2791 38024 2792 38076
rect 100 38016 2792 38024
rect 100 37964 2249 38016
rect 2301 37964 2315 38016
rect 2367 38011 2792 38016
rect 2367 37964 2673 38011
rect 100 37959 2673 37964
rect 2725 37959 2739 38011
rect 2791 37959 2792 38011
tri 2792 37988 3002 38198 nw
rect 100 37952 2792 37959
rect 100 37900 2249 37952
rect 2301 37900 2315 37952
rect 2367 37946 2792 37952
rect 2367 37900 2673 37946
rect 100 37894 2673 37900
rect 2725 37894 2739 37946
rect 2791 37894 2792 37946
rect 100 37888 2792 37894
rect 100 37836 2249 37888
rect 2301 37836 2315 37888
rect 2367 37881 2792 37888
rect 2367 37836 2673 37881
rect 100 37829 2673 37836
rect 2725 37829 2739 37881
rect 2791 37829 2792 37881
rect 100 37824 2792 37829
rect 100 37772 2249 37824
rect 2301 37772 2315 37824
rect 2367 37816 2792 37824
rect 2367 37772 2673 37816
rect 100 37764 2673 37772
rect 2725 37764 2739 37816
rect 2791 37764 2792 37816
rect 100 37760 2792 37764
rect 100 37708 2249 37760
rect 2301 37708 2315 37760
rect 2367 37751 2792 37760
rect 2367 37708 2673 37751
rect 100 37699 2673 37708
rect 2725 37699 2739 37751
rect 2791 37699 2792 37751
rect 100 37696 2792 37699
rect 100 37644 2249 37696
rect 2301 37644 2315 37696
rect 2367 37686 2792 37696
rect 2367 37644 2673 37686
rect 100 37634 2673 37644
rect 2725 37634 2739 37686
rect 2791 37634 2792 37686
rect 100 37632 2792 37634
rect 100 37580 2249 37632
rect 2301 37580 2315 37632
rect 2367 37621 2792 37632
rect 2367 37580 2673 37621
rect 100 37569 2673 37580
rect 2725 37569 2739 37621
rect 2791 37569 2792 37621
rect 100 37568 2792 37569
rect 100 37516 2249 37568
rect 2301 37516 2315 37568
rect 2367 37556 2792 37568
rect 2367 37516 2673 37556
rect 100 37504 2673 37516
rect 2725 37504 2739 37556
rect 2791 37504 2792 37556
rect 100 37452 2249 37504
rect 2301 37452 2315 37504
rect 2367 37491 2792 37504
rect 2367 37452 2673 37491
rect 100 37440 2673 37452
rect 100 37388 2249 37440
rect 2301 37388 2315 37440
rect 2367 37439 2673 37440
rect 2725 37439 2739 37491
rect 2791 37439 2792 37491
rect 2367 37426 2792 37439
rect 2367 37388 2673 37426
rect 100 37376 2673 37388
rect 100 37324 2249 37376
rect 2301 37324 2315 37376
rect 2367 37374 2673 37376
rect 2725 37374 2739 37426
rect 2791 37374 2792 37426
rect 2367 37324 2792 37374
rect 100 37312 2792 37324
rect 100 37260 2249 37312
rect 2301 37260 2315 37312
rect 2367 37260 2792 37312
rect 100 37248 2792 37260
rect 100 37196 2249 37248
rect 2301 37196 2315 37248
rect 2367 37196 2792 37248
rect 100 37184 2792 37196
rect 100 37132 2249 37184
rect 2301 37132 2315 37184
rect 2367 37132 2792 37184
rect 100 37120 2792 37132
rect 100 37068 2249 37120
rect 2301 37068 2315 37120
rect 2367 37068 2792 37120
rect 100 37056 2792 37068
rect 100 37004 2249 37056
rect 2301 37004 2315 37056
rect 2367 37004 2792 37056
rect 2950 37892 13317 37898
rect 3002 37840 3016 37892
rect 3068 37840 3504 37892
rect 3569 37840 3570 37892
rect 2950 37836 3513 37840
rect 3569 37836 3594 37840
rect 3650 37836 3675 37892
rect 3731 37836 3756 37892
rect 3812 37836 3837 37892
rect 3893 37836 3918 37892
rect 5014 37840 5166 37892
rect 5284 37840 5297 37892
rect 2950 37825 3918 37836
rect 5014 37836 5216 37840
rect 5272 37836 5297 37840
rect 5353 37836 5378 37892
rect 5434 37836 5459 37892
rect 5515 37836 5540 37892
rect 5596 37836 5621 37892
rect 5677 37836 5702 37892
rect 5772 37840 5783 37892
rect 5758 37836 5783 37840
rect 5839 37836 5864 37892
rect 5920 37836 5945 37892
rect 6001 37836 6026 37892
rect 6082 37836 6107 37892
rect 6163 37836 6188 37892
rect 6244 37836 6269 37892
rect 6326 37840 6340 37892
rect 6325 37836 6350 37840
rect 6406 37836 6431 37892
rect 6487 37836 6512 37892
rect 6568 37836 6593 37892
rect 6649 37836 6674 37892
rect 6730 37836 6755 37892
rect 6811 37840 6828 37892
rect 6892 37840 6894 37892
rect 6811 37836 6836 37840
rect 6892 37836 6917 37840
rect 6973 37836 6998 37892
rect 7054 37836 7079 37892
rect 7135 37836 7160 37892
rect 5014 37825 7160 37836
rect 3002 37773 3016 37825
rect 3068 37773 3504 37825
rect 3556 37812 3570 37825
rect 3622 37812 3918 37825
rect 3569 37773 3570 37812
rect 2950 37758 3513 37773
rect 3569 37758 3594 37773
rect 3002 37706 3016 37758
rect 3068 37706 3504 37758
rect 3569 37756 3570 37758
rect 3650 37756 3675 37812
rect 3731 37756 3756 37812
rect 3812 37756 3837 37812
rect 3893 37756 3918 37812
rect 5014 37773 5166 37825
rect 5218 37812 5232 37825
rect 5284 37812 5720 37825
rect 5772 37812 5786 37825
rect 5838 37812 6274 37825
rect 5284 37773 5297 37812
rect 5014 37758 5216 37773
rect 5272 37758 5297 37773
rect 3556 37732 3570 37756
rect 3622 37732 3918 37756
rect 3569 37706 3570 37732
rect 2950 37691 3513 37706
rect 3569 37691 3594 37706
rect 3002 37639 3016 37691
rect 3068 37639 3504 37691
rect 3569 37676 3570 37691
rect 3650 37676 3675 37732
rect 3731 37676 3756 37732
rect 3812 37676 3837 37732
rect 3893 37676 3918 37732
rect 5014 37706 5166 37758
rect 5284 37756 5297 37758
rect 5353 37756 5378 37812
rect 5434 37756 5459 37812
rect 5515 37756 5540 37812
rect 5596 37756 5621 37812
rect 5677 37756 5702 37812
rect 5772 37773 5783 37812
rect 5758 37758 5783 37773
rect 5772 37756 5783 37758
rect 5839 37756 5864 37812
rect 5920 37756 5945 37812
rect 6001 37756 6026 37812
rect 6082 37756 6107 37812
rect 6163 37756 6188 37812
rect 6244 37756 6269 37812
rect 6326 37773 6340 37825
rect 6392 37812 6828 37825
rect 6880 37812 6894 37825
rect 6946 37812 7160 37825
rect 6325 37758 6350 37773
rect 5218 37732 5232 37756
rect 5284 37732 5720 37756
rect 5772 37732 5786 37756
rect 5838 37732 6274 37756
rect 5284 37706 5297 37732
rect 5014 37691 5216 37706
rect 5272 37691 5297 37706
rect 3556 37652 3570 37676
rect 3622 37652 3918 37676
rect 3569 37639 3570 37652
rect 2950 37624 3513 37639
rect 3569 37624 3594 37639
rect 3002 37572 3016 37624
rect 3068 37572 3504 37624
rect 3569 37596 3570 37624
rect 3650 37596 3675 37652
rect 3731 37596 3756 37652
rect 3812 37596 3837 37652
rect 3893 37596 3918 37652
rect 5014 37639 5166 37691
rect 5284 37676 5297 37691
rect 5353 37676 5378 37732
rect 5434 37676 5459 37732
rect 5515 37676 5540 37732
rect 5596 37676 5621 37732
rect 5677 37676 5702 37732
rect 5772 37706 5783 37732
rect 5758 37691 5783 37706
rect 5772 37676 5783 37691
rect 5839 37676 5864 37732
rect 5920 37676 5945 37732
rect 6001 37676 6026 37732
rect 6082 37676 6107 37732
rect 6163 37676 6188 37732
rect 6244 37676 6269 37732
rect 6326 37706 6340 37758
rect 6406 37756 6431 37812
rect 6487 37756 6512 37812
rect 6568 37756 6593 37812
rect 6649 37756 6674 37812
rect 6730 37756 6755 37812
rect 6811 37773 6828 37812
rect 6892 37773 6894 37812
rect 6811 37758 6836 37773
rect 6892 37758 6917 37773
rect 6811 37756 6828 37758
rect 6892 37756 6894 37758
rect 6973 37756 6998 37812
rect 7054 37756 7079 37812
rect 7135 37756 7160 37812
rect 6392 37732 6828 37756
rect 6880 37732 6894 37756
rect 6946 37732 7160 37756
rect 6325 37691 6350 37706
rect 5218 37652 5232 37676
rect 5284 37652 5720 37676
rect 5772 37652 5786 37676
rect 5838 37652 6274 37676
rect 5284 37639 5297 37652
rect 5014 37624 5216 37639
rect 5272 37624 5297 37639
rect 3556 37572 3570 37596
rect 3622 37572 3918 37596
rect 5014 37572 5166 37624
rect 5284 37596 5297 37624
rect 5353 37596 5378 37652
rect 5434 37596 5459 37652
rect 5515 37596 5540 37652
rect 5596 37596 5621 37652
rect 5677 37596 5702 37652
rect 5772 37639 5783 37652
rect 5758 37624 5783 37639
rect 5772 37596 5783 37624
rect 5839 37596 5864 37652
rect 5920 37596 5945 37652
rect 6001 37596 6026 37652
rect 6082 37596 6107 37652
rect 6163 37596 6188 37652
rect 6244 37596 6269 37652
rect 6326 37639 6340 37691
rect 6406 37676 6431 37732
rect 6487 37676 6512 37732
rect 6568 37676 6593 37732
rect 6649 37676 6674 37732
rect 6730 37676 6755 37732
rect 6811 37706 6828 37732
rect 6892 37706 6894 37732
rect 6811 37691 6836 37706
rect 6892 37691 6917 37706
rect 6811 37676 6828 37691
rect 6892 37676 6894 37691
rect 6973 37676 6998 37732
rect 7054 37676 7079 37732
rect 7135 37676 7160 37732
rect 6392 37652 6828 37676
rect 6880 37652 6894 37676
rect 6946 37652 7160 37676
rect 6325 37624 6350 37639
rect 5218 37572 5232 37596
rect 5284 37572 5720 37596
rect 5772 37572 5786 37596
rect 5838 37572 6274 37596
rect 6326 37572 6340 37624
rect 6406 37596 6431 37652
rect 6487 37596 6512 37652
rect 6568 37596 6593 37652
rect 6649 37596 6674 37652
rect 6730 37596 6755 37652
rect 6811 37639 6828 37652
rect 6892 37639 6894 37652
rect 6811 37624 6836 37639
rect 6892 37624 6917 37639
rect 6811 37596 6828 37624
rect 6892 37596 6894 37624
rect 6973 37596 6998 37652
rect 7054 37596 7079 37652
rect 7135 37596 7160 37652
rect 6392 37572 6828 37596
rect 6880 37572 6894 37596
rect 6946 37572 7160 37596
rect 2950 37557 3513 37572
rect 3569 37557 3594 37572
rect 3002 37505 3016 37557
rect 3068 37505 3504 37557
rect 3569 37516 3570 37557
rect 3650 37516 3675 37572
rect 3731 37516 3756 37572
rect 3812 37516 3837 37572
rect 3893 37516 3918 37572
rect 5014 37557 5216 37572
rect 5272 37557 5297 37572
rect 3556 37505 3570 37516
rect 3622 37505 3918 37516
rect 5014 37505 5166 37557
rect 5284 37516 5297 37557
rect 5353 37516 5378 37572
rect 5434 37516 5459 37572
rect 5515 37516 5540 37572
rect 5596 37516 5621 37572
rect 5677 37516 5702 37572
rect 5758 37557 5783 37572
rect 5772 37516 5783 37557
rect 5839 37516 5864 37572
rect 5920 37516 5945 37572
rect 6001 37516 6026 37572
rect 6082 37516 6107 37572
rect 6163 37516 6188 37572
rect 6244 37516 6269 37572
rect 6325 37557 6350 37572
rect 5218 37505 5232 37516
rect 5284 37505 5720 37516
rect 5772 37505 5786 37516
rect 5838 37505 6274 37516
rect 6326 37505 6340 37557
rect 6406 37516 6431 37572
rect 6487 37516 6512 37572
rect 6568 37516 6593 37572
rect 6649 37516 6674 37572
rect 6730 37516 6755 37572
rect 6811 37557 6836 37572
rect 6892 37557 6917 37572
rect 6811 37516 6828 37557
rect 6892 37516 6894 37557
rect 6973 37516 6998 37572
rect 7054 37516 7079 37572
rect 7135 37516 7160 37572
rect 6392 37505 6828 37516
rect 6880 37505 6894 37516
rect 6946 37505 7160 37516
rect 2950 37492 3918 37505
rect 2950 37490 3513 37492
rect 3569 37490 3594 37492
rect 3002 37438 3016 37490
rect 3068 37438 3504 37490
rect 3569 37438 3570 37490
rect 2950 37436 3513 37438
rect 3569 37436 3594 37438
rect 3650 37436 3675 37492
rect 3731 37436 3756 37492
rect 3812 37436 3837 37492
rect 3893 37436 3918 37492
rect 5014 37492 7160 37505
rect 5014 37490 5216 37492
rect 5272 37490 5297 37492
rect 5014 37438 5166 37490
rect 5284 37438 5297 37490
rect 2950 37423 3918 37436
rect 5014 37436 5216 37438
rect 5272 37436 5297 37438
rect 5353 37436 5378 37492
rect 5434 37436 5459 37492
rect 5515 37436 5540 37492
rect 5596 37436 5621 37492
rect 5677 37436 5702 37492
rect 5758 37490 5783 37492
rect 5772 37438 5783 37490
rect 5758 37436 5783 37438
rect 5839 37436 5864 37492
rect 5920 37436 5945 37492
rect 6001 37436 6026 37492
rect 6082 37436 6107 37492
rect 6163 37436 6188 37492
rect 6244 37436 6269 37492
rect 6325 37490 6350 37492
rect 6326 37438 6340 37490
rect 6325 37436 6350 37438
rect 6406 37436 6431 37492
rect 6487 37436 6512 37492
rect 6568 37436 6593 37492
rect 6649 37436 6674 37492
rect 6730 37436 6755 37492
rect 6811 37490 6836 37492
rect 6892 37490 6917 37492
rect 6811 37438 6828 37490
rect 6892 37438 6894 37490
rect 6811 37436 6836 37438
rect 6892 37436 6917 37438
rect 6973 37436 6998 37492
rect 7054 37436 7079 37492
rect 7135 37436 7160 37492
rect 5014 37423 7160 37436
rect 3002 37371 3016 37423
rect 3068 37371 3504 37423
rect 3556 37412 3570 37423
rect 3622 37412 3918 37423
rect 3569 37371 3570 37412
rect 2950 37356 3513 37371
rect 3569 37356 3594 37371
rect 3650 37356 3675 37412
rect 3731 37356 3756 37412
rect 3812 37356 3837 37412
rect 3893 37356 3918 37412
rect 5014 37371 5166 37423
rect 5218 37412 5232 37423
rect 5284 37412 5720 37423
rect 5772 37412 5786 37423
rect 5838 37412 6274 37423
rect 5284 37371 5297 37412
rect 5014 37356 5216 37371
rect 5272 37356 5297 37371
rect 5353 37356 5378 37412
rect 5434 37356 5459 37412
rect 5515 37356 5540 37412
rect 5596 37356 5621 37412
rect 5677 37356 5702 37412
rect 5772 37371 5783 37412
rect 5758 37356 5783 37371
rect 5839 37356 5864 37412
rect 5920 37356 5945 37412
rect 6001 37356 6026 37412
rect 6082 37356 6107 37412
rect 6163 37356 6188 37412
rect 6244 37356 6269 37412
rect 6326 37371 6340 37423
rect 6392 37412 6828 37423
rect 6880 37412 6894 37423
rect 6946 37412 7160 37423
rect 6325 37356 6350 37371
rect 6406 37356 6431 37412
rect 6487 37356 6512 37412
rect 6568 37356 6593 37412
rect 6649 37356 6674 37412
rect 6730 37356 6755 37412
rect 6811 37371 6828 37412
rect 6892 37371 6894 37412
rect 6811 37356 6836 37371
rect 6892 37356 6917 37371
rect 6973 37356 6998 37412
rect 7054 37356 7079 37412
rect 7135 37356 7160 37412
rect 3002 37304 3016 37356
rect 3068 37304 3504 37356
rect 3556 37332 3570 37356
rect 3622 37332 3918 37356
rect 3569 37304 3570 37332
rect 2950 37289 3513 37304
rect 3569 37289 3594 37304
rect 3002 37237 3016 37289
rect 3068 37237 3504 37289
rect 3569 37276 3570 37289
rect 3650 37276 3675 37332
rect 3731 37276 3756 37332
rect 3812 37276 3837 37332
rect 3893 37276 3918 37332
rect 5014 37304 5166 37356
rect 5218 37332 5232 37356
rect 5284 37332 5720 37356
rect 5772 37332 5786 37356
rect 5838 37332 6274 37356
rect 5284 37304 5297 37332
rect 5014 37289 5216 37304
rect 5272 37289 5297 37304
rect 3556 37252 3570 37276
rect 3622 37252 3918 37276
rect 3569 37237 3570 37252
rect 2950 37222 3513 37237
rect 3569 37222 3594 37237
rect 3002 37170 3016 37222
rect 3068 37170 3504 37222
rect 3569 37196 3570 37222
rect 3650 37196 3675 37252
rect 3731 37196 3756 37252
rect 3812 37196 3837 37252
rect 3893 37196 3918 37252
rect 5014 37237 5166 37289
rect 5284 37276 5297 37289
rect 5353 37276 5378 37332
rect 5434 37276 5459 37332
rect 5515 37276 5540 37332
rect 5596 37276 5621 37332
rect 5677 37276 5702 37332
rect 5772 37304 5783 37332
rect 5758 37289 5783 37304
rect 5772 37276 5783 37289
rect 5839 37276 5864 37332
rect 5920 37276 5945 37332
rect 6001 37276 6026 37332
rect 6082 37276 6107 37332
rect 6163 37276 6188 37332
rect 6244 37276 6269 37332
rect 6326 37304 6340 37356
rect 6392 37332 6828 37356
rect 6880 37332 6894 37356
rect 6946 37332 7160 37356
rect 6325 37289 6350 37304
rect 5218 37252 5232 37276
rect 5284 37252 5720 37276
rect 5772 37252 5786 37276
rect 5838 37252 6274 37276
rect 5284 37237 5297 37252
rect 5014 37222 5216 37237
rect 5272 37222 5297 37237
rect 3556 37172 3570 37196
rect 3622 37172 3918 37196
rect 3569 37170 3570 37172
rect 2950 37155 3513 37170
rect 3569 37155 3594 37170
rect 3002 37103 3016 37155
rect 3068 37103 3504 37155
rect 3569 37116 3570 37155
rect 3650 37116 3675 37172
rect 3731 37116 3756 37172
rect 3812 37116 3837 37172
rect 3893 37116 3918 37172
rect 5014 37170 5166 37222
rect 5284 37196 5297 37222
rect 5353 37196 5378 37252
rect 5434 37196 5459 37252
rect 5515 37196 5540 37252
rect 5596 37196 5621 37252
rect 5677 37196 5702 37252
rect 5772 37237 5783 37252
rect 5758 37222 5783 37237
rect 5772 37196 5783 37222
rect 5839 37196 5864 37252
rect 5920 37196 5945 37252
rect 6001 37196 6026 37252
rect 6082 37196 6107 37252
rect 6163 37196 6188 37252
rect 6244 37196 6269 37252
rect 6326 37237 6340 37289
rect 6406 37276 6431 37332
rect 6487 37276 6512 37332
rect 6568 37276 6593 37332
rect 6649 37276 6674 37332
rect 6730 37276 6755 37332
rect 6811 37304 6828 37332
rect 6892 37304 6894 37332
rect 6811 37289 6836 37304
rect 6892 37289 6917 37304
rect 6811 37276 6828 37289
rect 6892 37276 6894 37289
rect 6973 37276 6998 37332
rect 7054 37276 7079 37332
rect 7135 37276 7160 37332
rect 6392 37252 6828 37276
rect 6880 37252 6894 37276
rect 6946 37252 7160 37276
rect 6325 37222 6350 37237
rect 5218 37172 5232 37196
rect 5284 37172 5720 37196
rect 5772 37172 5786 37196
rect 5838 37172 6274 37196
rect 5284 37170 5297 37172
rect 5014 37155 5216 37170
rect 5272 37155 5297 37170
rect 3556 37103 3570 37116
rect 3622 37103 3918 37116
rect 5014 37103 5166 37155
rect 5284 37116 5297 37155
rect 5353 37116 5378 37172
rect 5434 37116 5459 37172
rect 5515 37116 5540 37172
rect 5596 37116 5621 37172
rect 5677 37116 5702 37172
rect 5772 37170 5783 37172
rect 5758 37155 5783 37170
rect 5772 37116 5783 37155
rect 5839 37116 5864 37172
rect 5920 37116 5945 37172
rect 6001 37116 6026 37172
rect 6082 37116 6107 37172
rect 6163 37116 6188 37172
rect 6244 37116 6269 37172
rect 6326 37170 6340 37222
rect 6406 37196 6431 37252
rect 6487 37196 6512 37252
rect 6568 37196 6593 37252
rect 6649 37196 6674 37252
rect 6730 37196 6755 37252
rect 6811 37237 6828 37252
rect 6892 37237 6894 37252
rect 6811 37222 6836 37237
rect 6892 37222 6917 37237
rect 6811 37196 6828 37222
rect 6892 37196 6894 37222
rect 6973 37196 6998 37252
rect 7054 37196 7079 37252
rect 7135 37196 7160 37252
rect 6392 37172 6828 37196
rect 6880 37172 6894 37196
rect 6946 37172 7160 37196
rect 6325 37155 6350 37170
rect 5218 37103 5232 37116
rect 5284 37103 5720 37116
rect 5772 37103 5786 37116
rect 5838 37103 6274 37116
rect 6326 37103 6340 37155
rect 6406 37116 6431 37172
rect 6487 37116 6512 37172
rect 6568 37116 6593 37172
rect 6649 37116 6674 37172
rect 6730 37116 6755 37172
rect 6811 37170 6828 37172
rect 6892 37170 6894 37172
rect 6811 37155 6836 37170
rect 6892 37155 6917 37170
rect 6811 37116 6828 37155
rect 6892 37116 6894 37155
rect 6973 37116 6998 37172
rect 7054 37116 7079 37172
rect 7135 37116 7160 37172
rect 6392 37103 6828 37116
rect 6880 37103 6894 37116
rect 6946 37103 7160 37116
rect 2950 37092 3918 37103
rect 2950 37088 3513 37092
rect 3569 37088 3594 37092
rect 3002 37036 3016 37088
rect 3068 37036 3504 37088
rect 3569 37036 3570 37088
rect 3650 37036 3675 37092
rect 3731 37036 3756 37092
rect 3812 37036 3837 37092
rect 3893 37036 3918 37092
rect 5014 37092 7160 37103
rect 5014 37088 5216 37092
rect 5272 37088 5297 37092
rect 5014 37036 5166 37088
rect 5284 37036 5297 37088
rect 5353 37036 5378 37092
rect 5434 37036 5459 37092
rect 5515 37036 5540 37092
rect 5596 37036 5621 37092
rect 5677 37036 5702 37092
rect 5758 37088 5783 37092
rect 5772 37036 5783 37088
rect 5839 37036 5864 37092
rect 5920 37036 5945 37092
rect 6001 37036 6026 37092
rect 6082 37036 6107 37092
rect 6163 37036 6188 37092
rect 6244 37036 6269 37092
rect 6325 37088 6350 37092
rect 6326 37036 6340 37088
rect 6406 37036 6431 37092
rect 6487 37036 6512 37092
rect 6568 37036 6593 37092
rect 6649 37036 6674 37092
rect 6730 37036 6755 37092
rect 6811 37088 6836 37092
rect 6892 37088 6917 37092
rect 6811 37036 6828 37088
rect 6892 37036 6894 37088
rect 6973 37036 6998 37092
rect 7054 37036 7079 37092
rect 7135 37036 7160 37092
rect 7376 37840 7382 37892
rect 7434 37840 7448 37892
rect 7500 37840 7598 37892
rect 7376 37836 7598 37840
rect 7654 37836 7679 37892
rect 7735 37836 7760 37892
rect 7816 37836 7841 37892
rect 7897 37836 7922 37892
rect 7988 37840 8002 37892
rect 7978 37836 8003 37840
rect 8059 37836 8084 37892
rect 8140 37836 8165 37892
rect 8221 37836 8246 37892
rect 8302 37836 8327 37892
rect 8383 37836 8408 37892
rect 8464 37836 8489 37892
rect 8545 37840 8556 37892
rect 8545 37836 8570 37840
rect 8626 37836 8651 37892
rect 8707 37836 8732 37892
rect 8788 37836 8813 37892
rect 8869 37836 8894 37892
rect 8950 37836 8975 37892
rect 9031 37840 9044 37892
rect 9031 37836 9056 37840
rect 9112 37836 9137 37840
rect 9193 37836 9218 37892
rect 9274 37836 9299 37892
rect 9355 37836 9380 37892
rect 9436 37836 9461 37892
rect 9517 37836 9542 37892
rect 7376 37825 9542 37836
rect 9758 37836 9983 37892
rect 10039 37836 10064 37892
rect 10120 37836 10145 37892
rect 10204 37840 10218 37892
rect 10201 37836 10226 37840
rect 10282 37836 10307 37892
rect 10363 37836 10388 37892
rect 10444 37836 10469 37892
rect 10525 37836 10550 37892
rect 10606 37836 10631 37892
rect 10687 37840 10706 37892
rect 10768 37840 10772 37892
rect 10687 37836 10712 37840
rect 10768 37836 10793 37840
rect 10849 37836 10874 37892
rect 10930 37836 10955 37892
rect 11011 37836 11036 37892
rect 11092 37836 11117 37892
rect 11173 37836 11198 37892
rect 11254 37840 11260 37892
rect 11254 37836 11279 37840
rect 11335 37836 11360 37840
rect 11416 37836 11441 37892
rect 12057 37840 12368 37892
rect 12420 37840 12434 37892
rect 12486 37840 12922 37892
rect 12974 37840 12988 37892
rect 13040 37840 13317 37892
rect 9758 37825 11441 37836
rect 12057 37825 13317 37840
rect 7376 37773 7382 37825
rect 7434 37773 7448 37825
rect 7500 37812 7936 37825
rect 7500 37773 7598 37812
rect 7376 37758 7598 37773
rect 7376 37706 7382 37758
rect 7434 37706 7448 37758
rect 7500 37756 7598 37758
rect 7654 37756 7679 37812
rect 7735 37756 7760 37812
rect 7816 37756 7841 37812
rect 7897 37756 7922 37812
rect 7988 37773 8002 37825
rect 8054 37812 8490 37825
rect 8542 37812 8556 37825
rect 8608 37812 9044 37825
rect 9096 37812 9110 37825
rect 9162 37812 9542 37825
rect 7978 37758 8003 37773
rect 7500 37732 7936 37756
rect 7500 37706 7598 37732
rect 7376 37691 7598 37706
rect 7376 37639 7382 37691
rect 7434 37639 7448 37691
rect 7500 37676 7598 37691
rect 7654 37676 7679 37732
rect 7735 37676 7760 37732
rect 7816 37676 7841 37732
rect 7897 37676 7922 37732
rect 7988 37706 8002 37758
rect 8059 37756 8084 37812
rect 8140 37756 8165 37812
rect 8221 37756 8246 37812
rect 8302 37756 8327 37812
rect 8383 37756 8408 37812
rect 8464 37756 8489 37812
rect 8545 37773 8556 37812
rect 8545 37758 8570 37773
rect 8545 37756 8556 37758
rect 8626 37756 8651 37812
rect 8707 37756 8732 37812
rect 8788 37756 8813 37812
rect 8869 37756 8894 37812
rect 8950 37756 8975 37812
rect 9031 37773 9044 37812
rect 9031 37758 9056 37773
rect 9112 37758 9137 37773
rect 9031 37756 9044 37758
rect 9193 37756 9218 37812
rect 9274 37756 9299 37812
rect 9355 37756 9380 37812
rect 9436 37756 9461 37812
rect 9517 37756 9542 37812
rect 9758 37812 10152 37825
rect 8054 37732 8490 37756
rect 8542 37732 8556 37756
rect 8608 37732 9044 37756
rect 9096 37732 9110 37756
rect 9162 37732 9542 37756
rect 7978 37691 8003 37706
rect 7500 37652 7936 37676
rect 7500 37639 7598 37652
rect 7376 37624 7598 37639
rect 7376 37572 7382 37624
rect 7434 37572 7448 37624
rect 7500 37596 7598 37624
rect 7654 37596 7679 37652
rect 7735 37596 7760 37652
rect 7816 37596 7841 37652
rect 7897 37596 7922 37652
rect 7988 37639 8002 37691
rect 8059 37676 8084 37732
rect 8140 37676 8165 37732
rect 8221 37676 8246 37732
rect 8302 37676 8327 37732
rect 8383 37676 8408 37732
rect 8464 37676 8489 37732
rect 8545 37706 8556 37732
rect 8545 37691 8570 37706
rect 8545 37676 8556 37691
rect 8626 37676 8651 37732
rect 8707 37676 8732 37732
rect 8788 37676 8813 37732
rect 8869 37676 8894 37732
rect 8950 37676 8975 37732
rect 9031 37706 9044 37732
rect 9031 37691 9056 37706
rect 9112 37691 9137 37706
rect 9031 37676 9044 37691
rect 9193 37676 9218 37732
rect 9274 37676 9299 37732
rect 9355 37676 9380 37732
rect 9436 37676 9461 37732
rect 9517 37676 9542 37732
rect 9758 37756 9983 37812
rect 10039 37756 10064 37812
rect 10120 37756 10145 37812
rect 10204 37773 10218 37825
rect 10270 37812 10706 37825
rect 10758 37812 10772 37825
rect 10824 37812 11260 37825
rect 11312 37812 11326 37825
rect 11378 37812 11441 37825
rect 10201 37758 10226 37773
rect 9758 37732 10152 37756
rect 8054 37652 8490 37676
rect 8542 37652 8556 37676
rect 8608 37652 9044 37676
rect 9096 37652 9110 37676
rect 9162 37652 9542 37676
rect 7978 37624 8003 37639
rect 7500 37572 7936 37596
rect 7988 37572 8002 37624
rect 8059 37596 8084 37652
rect 8140 37596 8165 37652
rect 8221 37596 8246 37652
rect 8302 37596 8327 37652
rect 8383 37596 8408 37652
rect 8464 37596 8489 37652
rect 8545 37639 8556 37652
rect 8545 37624 8570 37639
rect 8545 37596 8556 37624
rect 8626 37596 8651 37652
rect 8707 37596 8732 37652
rect 8788 37596 8813 37652
rect 8869 37596 8894 37652
rect 8950 37596 8975 37652
rect 9031 37639 9044 37652
rect 9031 37624 9056 37639
rect 9112 37624 9137 37639
rect 9031 37596 9044 37624
rect 9193 37596 9218 37652
rect 9274 37596 9299 37652
rect 9355 37596 9380 37652
rect 9436 37596 9461 37652
rect 9517 37596 9542 37652
rect 9758 37676 9983 37732
rect 10039 37676 10064 37732
rect 10120 37676 10145 37732
rect 10204 37706 10218 37758
rect 10282 37756 10307 37812
rect 10363 37756 10388 37812
rect 10444 37756 10469 37812
rect 10525 37756 10550 37812
rect 10606 37756 10631 37812
rect 10687 37773 10706 37812
rect 10768 37773 10772 37812
rect 10687 37758 10712 37773
rect 10768 37758 10793 37773
rect 10687 37756 10706 37758
rect 10768 37756 10772 37758
rect 10849 37756 10874 37812
rect 10930 37756 10955 37812
rect 11011 37756 11036 37812
rect 11092 37756 11117 37812
rect 11173 37756 11198 37812
rect 11254 37773 11260 37812
rect 11254 37758 11279 37773
rect 11335 37758 11360 37773
rect 11254 37756 11260 37758
rect 11416 37756 11441 37812
rect 12057 37773 12368 37825
rect 12420 37773 12434 37825
rect 12486 37773 12922 37825
rect 12974 37773 12988 37825
rect 13040 37773 13317 37825
rect 12057 37758 13317 37773
rect 10270 37732 10706 37756
rect 10758 37732 10772 37756
rect 10824 37732 11260 37756
rect 11312 37732 11326 37756
rect 11378 37732 11441 37756
rect 10201 37691 10226 37706
rect 9758 37652 10152 37676
rect 8054 37572 8490 37596
rect 8542 37572 8556 37596
rect 8608 37572 9044 37596
rect 9096 37572 9110 37596
rect 9162 37572 9542 37596
rect 9758 37596 9983 37652
rect 10039 37596 10064 37652
rect 10120 37596 10145 37652
rect 10204 37639 10218 37691
rect 10282 37676 10307 37732
rect 10363 37676 10388 37732
rect 10444 37676 10469 37732
rect 10525 37676 10550 37732
rect 10606 37676 10631 37732
rect 10687 37706 10706 37732
rect 10768 37706 10772 37732
rect 10687 37691 10712 37706
rect 10768 37691 10793 37706
rect 10687 37676 10706 37691
rect 10768 37676 10772 37691
rect 10849 37676 10874 37732
rect 10930 37676 10955 37732
rect 11011 37676 11036 37732
rect 11092 37676 11117 37732
rect 11173 37676 11198 37732
rect 11254 37706 11260 37732
rect 11254 37691 11279 37706
rect 11335 37691 11360 37706
rect 11254 37676 11260 37691
rect 11416 37676 11441 37732
rect 12057 37706 12368 37758
rect 12420 37706 12434 37758
rect 12486 37706 12922 37758
rect 12974 37706 12988 37758
rect 13040 37706 13317 37758
rect 12057 37691 13317 37706
rect 10270 37652 10706 37676
rect 10758 37652 10772 37676
rect 10824 37652 11260 37676
rect 11312 37652 11326 37676
rect 11378 37652 11441 37676
rect 10201 37624 10226 37639
rect 9758 37572 10152 37596
rect 10204 37572 10218 37624
rect 10282 37596 10307 37652
rect 10363 37596 10388 37652
rect 10444 37596 10469 37652
rect 10525 37596 10550 37652
rect 10606 37596 10631 37652
rect 10687 37639 10706 37652
rect 10768 37639 10772 37652
rect 10687 37624 10712 37639
rect 10768 37624 10793 37639
rect 10687 37596 10706 37624
rect 10768 37596 10772 37624
rect 10849 37596 10874 37652
rect 10930 37596 10955 37652
rect 11011 37596 11036 37652
rect 11092 37596 11117 37652
rect 11173 37596 11198 37652
rect 11254 37639 11260 37652
rect 11254 37624 11279 37639
rect 11335 37624 11360 37639
rect 11254 37596 11260 37624
rect 11416 37596 11441 37652
rect 12057 37639 12368 37691
rect 12420 37639 12434 37691
rect 12486 37639 12922 37691
rect 12974 37639 12988 37691
rect 13040 37639 13317 37691
rect 12057 37624 13317 37639
rect 10270 37572 10706 37596
rect 10758 37572 10772 37596
rect 10824 37572 11260 37596
rect 11312 37572 11326 37596
rect 11378 37572 11441 37596
rect 12057 37572 12368 37624
rect 12420 37572 12434 37624
rect 12486 37572 12922 37624
rect 12974 37572 12988 37624
rect 13040 37572 13317 37624
rect 7376 37557 7598 37572
rect 7376 37505 7382 37557
rect 7434 37505 7448 37557
rect 7500 37516 7598 37557
rect 7654 37516 7679 37572
rect 7735 37516 7760 37572
rect 7816 37516 7841 37572
rect 7897 37516 7922 37572
rect 7978 37557 8003 37572
rect 7500 37505 7936 37516
rect 7988 37505 8002 37557
rect 8059 37516 8084 37572
rect 8140 37516 8165 37572
rect 8221 37516 8246 37572
rect 8302 37516 8327 37572
rect 8383 37516 8408 37572
rect 8464 37516 8489 37572
rect 8545 37557 8570 37572
rect 8545 37516 8556 37557
rect 8626 37516 8651 37572
rect 8707 37516 8732 37572
rect 8788 37516 8813 37572
rect 8869 37516 8894 37572
rect 8950 37516 8975 37572
rect 9031 37557 9056 37572
rect 9112 37557 9137 37572
rect 9031 37516 9044 37557
rect 9193 37516 9218 37572
rect 9274 37516 9299 37572
rect 9355 37516 9380 37572
rect 9436 37516 9461 37572
rect 9517 37516 9542 37572
rect 8054 37505 8490 37516
rect 8542 37505 8556 37516
rect 8608 37505 9044 37516
rect 9096 37505 9110 37516
rect 9162 37505 9542 37516
rect 9758 37516 9983 37572
rect 10039 37516 10064 37572
rect 10120 37516 10145 37572
rect 10201 37557 10226 37572
rect 9758 37505 10152 37516
rect 10204 37505 10218 37557
rect 10282 37516 10307 37572
rect 10363 37516 10388 37572
rect 10444 37516 10469 37572
rect 10525 37516 10550 37572
rect 10606 37516 10631 37572
rect 10687 37557 10712 37572
rect 10768 37557 10793 37572
rect 10687 37516 10706 37557
rect 10768 37516 10772 37557
rect 10849 37516 10874 37572
rect 10930 37516 10955 37572
rect 11011 37516 11036 37572
rect 11092 37516 11117 37572
rect 11173 37516 11198 37572
rect 11254 37557 11279 37572
rect 11335 37557 11360 37572
rect 11254 37516 11260 37557
rect 11416 37516 11441 37572
rect 12057 37557 13317 37572
rect 10270 37505 10706 37516
rect 10758 37505 10772 37516
rect 10824 37505 11260 37516
rect 11312 37505 11326 37516
rect 11378 37505 11441 37516
rect 12057 37505 12368 37557
rect 12420 37505 12434 37557
rect 12486 37505 12922 37557
rect 12974 37505 12988 37557
rect 13040 37505 13317 37557
rect 7376 37492 9542 37505
rect 7376 37490 7598 37492
rect 7376 37438 7382 37490
rect 7434 37438 7448 37490
rect 7500 37438 7598 37490
rect 7376 37436 7598 37438
rect 7654 37436 7679 37492
rect 7735 37436 7760 37492
rect 7816 37436 7841 37492
rect 7897 37436 7922 37492
rect 7978 37490 8003 37492
rect 7988 37438 8002 37490
rect 7978 37436 8003 37438
rect 8059 37436 8084 37492
rect 8140 37436 8165 37492
rect 8221 37436 8246 37492
rect 8302 37436 8327 37492
rect 8383 37436 8408 37492
rect 8464 37436 8489 37492
rect 8545 37490 8570 37492
rect 8545 37438 8556 37490
rect 8545 37436 8570 37438
rect 8626 37436 8651 37492
rect 8707 37436 8732 37492
rect 8788 37436 8813 37492
rect 8869 37436 8894 37492
rect 8950 37436 8975 37492
rect 9031 37490 9056 37492
rect 9112 37490 9137 37492
rect 9031 37438 9044 37490
rect 9031 37436 9056 37438
rect 9112 37436 9137 37438
rect 9193 37436 9218 37492
rect 9274 37436 9299 37492
rect 9355 37436 9380 37492
rect 9436 37436 9461 37492
rect 9517 37436 9542 37492
rect 9758 37492 11441 37505
rect 7376 37423 9542 37436
rect 9758 37436 9983 37492
rect 10039 37436 10064 37492
rect 10120 37436 10145 37492
rect 10201 37490 10226 37492
rect 10204 37438 10218 37490
rect 10201 37436 10226 37438
rect 10282 37436 10307 37492
rect 10363 37436 10388 37492
rect 10444 37436 10469 37492
rect 10525 37436 10550 37492
rect 10606 37436 10631 37492
rect 10687 37490 10712 37492
rect 10768 37490 10793 37492
rect 10687 37438 10706 37490
rect 10768 37438 10772 37490
rect 10687 37436 10712 37438
rect 10768 37436 10793 37438
rect 10849 37436 10874 37492
rect 10930 37436 10955 37492
rect 11011 37436 11036 37492
rect 11092 37436 11117 37492
rect 11173 37436 11198 37492
rect 11254 37490 11279 37492
rect 11335 37490 11360 37492
rect 11254 37438 11260 37490
rect 11254 37436 11279 37438
rect 11335 37436 11360 37438
rect 11416 37436 11441 37492
rect 12057 37490 13317 37505
rect 12057 37438 12368 37490
rect 12420 37438 12434 37490
rect 12486 37438 12922 37490
rect 12974 37438 12988 37490
rect 13040 37438 13317 37490
rect 9758 37423 11441 37436
rect 12057 37423 13317 37438
rect 7376 37371 7382 37423
rect 7434 37371 7448 37423
rect 7500 37412 7936 37423
rect 7500 37371 7598 37412
rect 7376 37356 7598 37371
rect 7654 37356 7679 37412
rect 7735 37356 7760 37412
rect 7816 37356 7841 37412
rect 7897 37356 7922 37412
rect 7988 37371 8002 37423
rect 8054 37412 8490 37423
rect 8542 37412 8556 37423
rect 8608 37412 9044 37423
rect 9096 37412 9110 37423
rect 9162 37412 9542 37423
rect 7978 37356 8003 37371
rect 8059 37356 8084 37412
rect 8140 37356 8165 37412
rect 8221 37356 8246 37412
rect 8302 37356 8327 37412
rect 8383 37356 8408 37412
rect 8464 37356 8489 37412
rect 8545 37371 8556 37412
rect 8545 37356 8570 37371
rect 8626 37356 8651 37412
rect 8707 37356 8732 37412
rect 8788 37356 8813 37412
rect 8869 37356 8894 37412
rect 8950 37356 8975 37412
rect 9031 37371 9044 37412
rect 9031 37356 9056 37371
rect 9112 37356 9137 37371
rect 9193 37356 9218 37412
rect 9274 37356 9299 37412
rect 9355 37356 9380 37412
rect 9436 37356 9461 37412
rect 9517 37356 9542 37412
rect 9758 37412 10152 37423
rect 9758 37356 9983 37412
rect 10039 37356 10064 37412
rect 10120 37356 10145 37412
rect 10204 37371 10218 37423
rect 10270 37412 10706 37423
rect 10758 37412 10772 37423
rect 10824 37412 11260 37423
rect 11312 37412 11326 37423
rect 11378 37412 11441 37423
rect 10201 37356 10226 37371
rect 10282 37356 10307 37412
rect 10363 37356 10388 37412
rect 10444 37356 10469 37412
rect 10525 37356 10550 37412
rect 10606 37356 10631 37412
rect 10687 37371 10706 37412
rect 10768 37371 10772 37412
rect 10687 37356 10712 37371
rect 10768 37356 10793 37371
rect 10849 37356 10874 37412
rect 10930 37356 10955 37412
rect 11011 37356 11036 37412
rect 11092 37356 11117 37412
rect 11173 37356 11198 37412
rect 11254 37371 11260 37412
rect 11254 37356 11279 37371
rect 11335 37356 11360 37371
rect 11416 37356 11441 37412
rect 12057 37371 12368 37423
rect 12420 37371 12434 37423
rect 12486 37371 12922 37423
rect 12974 37371 12988 37423
rect 13040 37371 13317 37423
rect 12057 37356 13317 37371
rect 7376 37304 7382 37356
rect 7434 37304 7448 37356
rect 7500 37332 7936 37356
rect 7500 37304 7598 37332
rect 7376 37289 7598 37304
rect 7376 37237 7382 37289
rect 7434 37237 7448 37289
rect 7500 37276 7598 37289
rect 7654 37276 7679 37332
rect 7735 37276 7760 37332
rect 7816 37276 7841 37332
rect 7897 37276 7922 37332
rect 7988 37304 8002 37356
rect 8054 37332 8490 37356
rect 8542 37332 8556 37356
rect 8608 37332 9044 37356
rect 9096 37332 9110 37356
rect 9162 37332 9542 37356
rect 7978 37289 8003 37304
rect 7500 37252 7936 37276
rect 7500 37237 7598 37252
rect 7376 37222 7598 37237
rect 7376 37170 7382 37222
rect 7434 37170 7448 37222
rect 7500 37196 7598 37222
rect 7654 37196 7679 37252
rect 7735 37196 7760 37252
rect 7816 37196 7841 37252
rect 7897 37196 7922 37252
rect 7988 37237 8002 37289
rect 8059 37276 8084 37332
rect 8140 37276 8165 37332
rect 8221 37276 8246 37332
rect 8302 37276 8327 37332
rect 8383 37276 8408 37332
rect 8464 37276 8489 37332
rect 8545 37304 8556 37332
rect 8545 37289 8570 37304
rect 8545 37276 8556 37289
rect 8626 37276 8651 37332
rect 8707 37276 8732 37332
rect 8788 37276 8813 37332
rect 8869 37276 8894 37332
rect 8950 37276 8975 37332
rect 9031 37304 9044 37332
rect 9031 37289 9056 37304
rect 9112 37289 9137 37304
rect 9031 37276 9044 37289
rect 9193 37276 9218 37332
rect 9274 37276 9299 37332
rect 9355 37276 9380 37332
rect 9436 37276 9461 37332
rect 9517 37276 9542 37332
rect 9758 37332 10152 37356
rect 8054 37252 8490 37276
rect 8542 37252 8556 37276
rect 8608 37252 9044 37276
rect 9096 37252 9110 37276
rect 9162 37252 9542 37276
rect 7978 37222 8003 37237
rect 7500 37172 7936 37196
rect 7500 37170 7598 37172
rect 7376 37155 7598 37170
rect 7376 37103 7382 37155
rect 7434 37103 7448 37155
rect 7500 37116 7598 37155
rect 7654 37116 7679 37172
rect 7735 37116 7760 37172
rect 7816 37116 7841 37172
rect 7897 37116 7922 37172
rect 7988 37170 8002 37222
rect 8059 37196 8084 37252
rect 8140 37196 8165 37252
rect 8221 37196 8246 37252
rect 8302 37196 8327 37252
rect 8383 37196 8408 37252
rect 8464 37196 8489 37252
rect 8545 37237 8556 37252
rect 8545 37222 8570 37237
rect 8545 37196 8556 37222
rect 8626 37196 8651 37252
rect 8707 37196 8732 37252
rect 8788 37196 8813 37252
rect 8869 37196 8894 37252
rect 8950 37196 8975 37252
rect 9031 37237 9044 37252
rect 9031 37222 9056 37237
rect 9112 37222 9137 37237
rect 9031 37196 9044 37222
rect 9193 37196 9218 37252
rect 9274 37196 9299 37252
rect 9355 37196 9380 37252
rect 9436 37196 9461 37252
rect 9517 37196 9542 37252
rect 9758 37276 9983 37332
rect 10039 37276 10064 37332
rect 10120 37276 10145 37332
rect 10204 37304 10218 37356
rect 10270 37332 10706 37356
rect 10758 37332 10772 37356
rect 10824 37332 11260 37356
rect 11312 37332 11326 37356
rect 11378 37332 11441 37356
rect 10201 37289 10226 37304
rect 9758 37252 10152 37276
rect 8054 37172 8490 37196
rect 8542 37172 8556 37196
rect 8608 37172 9044 37196
rect 9096 37172 9110 37196
rect 9162 37172 9542 37196
rect 7978 37155 8003 37170
rect 7500 37103 7936 37116
rect 7988 37103 8002 37155
rect 8059 37116 8084 37172
rect 8140 37116 8165 37172
rect 8221 37116 8246 37172
rect 8302 37116 8327 37172
rect 8383 37116 8408 37172
rect 8464 37116 8489 37172
rect 8545 37170 8556 37172
rect 8545 37155 8570 37170
rect 8545 37116 8556 37155
rect 8626 37116 8651 37172
rect 8707 37116 8732 37172
rect 8788 37116 8813 37172
rect 8869 37116 8894 37172
rect 8950 37116 8975 37172
rect 9031 37170 9044 37172
rect 9031 37155 9056 37170
rect 9112 37155 9137 37170
rect 9031 37116 9044 37155
rect 9193 37116 9218 37172
rect 9274 37116 9299 37172
rect 9355 37116 9380 37172
rect 9436 37116 9461 37172
rect 9517 37116 9542 37172
rect 9758 37196 9983 37252
rect 10039 37196 10064 37252
rect 10120 37196 10145 37252
rect 10204 37237 10218 37289
rect 10282 37276 10307 37332
rect 10363 37276 10388 37332
rect 10444 37276 10469 37332
rect 10525 37276 10550 37332
rect 10606 37276 10631 37332
rect 10687 37304 10706 37332
rect 10768 37304 10772 37332
rect 10687 37289 10712 37304
rect 10768 37289 10793 37304
rect 10687 37276 10706 37289
rect 10768 37276 10772 37289
rect 10849 37276 10874 37332
rect 10930 37276 10955 37332
rect 11011 37276 11036 37332
rect 11092 37276 11117 37332
rect 11173 37276 11198 37332
rect 11254 37304 11260 37332
rect 11254 37289 11279 37304
rect 11335 37289 11360 37304
rect 11254 37276 11260 37289
rect 11416 37276 11441 37332
rect 12057 37304 12368 37356
rect 12420 37304 12434 37356
rect 12486 37304 12922 37356
rect 12974 37304 12988 37356
rect 13040 37304 13317 37356
rect 12057 37289 13317 37304
rect 10270 37252 10706 37276
rect 10758 37252 10772 37276
rect 10824 37252 11260 37276
rect 11312 37252 11326 37276
rect 11378 37252 11441 37276
rect 10201 37222 10226 37237
rect 9758 37172 10152 37196
rect 8054 37103 8490 37116
rect 8542 37103 8556 37116
rect 8608 37103 9044 37116
rect 9096 37103 9110 37116
rect 9162 37103 9542 37116
rect 9758 37116 9983 37172
rect 10039 37116 10064 37172
rect 10120 37116 10145 37172
rect 10204 37170 10218 37222
rect 10282 37196 10307 37252
rect 10363 37196 10388 37252
rect 10444 37196 10469 37252
rect 10525 37196 10550 37252
rect 10606 37196 10631 37252
rect 10687 37237 10706 37252
rect 10768 37237 10772 37252
rect 10687 37222 10712 37237
rect 10768 37222 10793 37237
rect 10687 37196 10706 37222
rect 10768 37196 10772 37222
rect 10849 37196 10874 37252
rect 10930 37196 10955 37252
rect 11011 37196 11036 37252
rect 11092 37196 11117 37252
rect 11173 37196 11198 37252
rect 11254 37237 11260 37252
rect 11254 37222 11279 37237
rect 11335 37222 11360 37237
rect 11254 37196 11260 37222
rect 11416 37196 11441 37252
rect 12057 37237 12368 37289
rect 12420 37237 12434 37289
rect 12486 37237 12922 37289
rect 12974 37237 12988 37289
rect 13040 37237 13317 37289
rect 12057 37222 13317 37237
rect 10270 37172 10706 37196
rect 10758 37172 10772 37196
rect 10824 37172 11260 37196
rect 11312 37172 11326 37196
rect 11378 37172 11441 37196
rect 10201 37155 10226 37170
rect 9758 37103 10152 37116
rect 10204 37103 10218 37155
rect 10282 37116 10307 37172
rect 10363 37116 10388 37172
rect 10444 37116 10469 37172
rect 10525 37116 10550 37172
rect 10606 37116 10631 37172
rect 10687 37170 10706 37172
rect 10768 37170 10772 37172
rect 10687 37155 10712 37170
rect 10768 37155 10793 37170
rect 10687 37116 10706 37155
rect 10768 37116 10772 37155
rect 10849 37116 10874 37172
rect 10930 37116 10955 37172
rect 11011 37116 11036 37172
rect 11092 37116 11117 37172
rect 11173 37116 11198 37172
rect 11254 37170 11260 37172
rect 11254 37155 11279 37170
rect 11335 37155 11360 37170
rect 11254 37116 11260 37155
rect 11416 37116 11441 37172
rect 12057 37170 12368 37222
rect 12420 37170 12434 37222
rect 12486 37170 12922 37222
rect 12974 37170 12988 37222
rect 13040 37170 13317 37222
rect 12057 37155 13317 37170
rect 10270 37103 10706 37116
rect 10758 37103 10772 37116
rect 10824 37103 11260 37116
rect 11312 37103 11326 37116
rect 11378 37103 11441 37116
rect 12057 37103 12368 37155
rect 12420 37103 12434 37155
rect 12486 37103 12922 37155
rect 12974 37103 12988 37155
rect 13040 37103 13317 37155
rect 7376 37092 9542 37103
rect 7376 37088 7598 37092
rect 7376 37036 7382 37088
rect 7434 37036 7448 37088
rect 7500 37036 7598 37088
rect 7654 37036 7679 37092
rect 7735 37036 7760 37092
rect 7816 37036 7841 37092
rect 7897 37036 7922 37092
rect 7978 37088 8003 37092
rect 7988 37036 8002 37088
rect 8059 37036 8084 37092
rect 8140 37036 8165 37092
rect 8221 37036 8246 37092
rect 8302 37036 8327 37092
rect 8383 37036 8408 37092
rect 8464 37036 8489 37092
rect 8545 37088 8570 37092
rect 8545 37036 8556 37088
rect 8626 37036 8651 37092
rect 8707 37036 8732 37092
rect 8788 37036 8813 37092
rect 8869 37036 8894 37092
rect 8950 37036 8975 37092
rect 9031 37088 9056 37092
rect 9112 37088 9137 37092
rect 9031 37036 9044 37088
rect 9193 37036 9218 37092
rect 9274 37036 9299 37092
rect 9355 37036 9380 37092
rect 9436 37036 9461 37092
rect 9517 37036 9542 37092
rect 9758 37092 11441 37103
rect 9758 37036 9983 37092
rect 10039 37036 10064 37092
rect 10120 37036 10145 37092
rect 10201 37088 10226 37092
rect 10204 37036 10218 37088
rect 10282 37036 10307 37092
rect 10363 37036 10388 37092
rect 10444 37036 10469 37092
rect 10525 37036 10550 37092
rect 10606 37036 10631 37092
rect 10687 37088 10712 37092
rect 10768 37088 10793 37092
rect 10687 37036 10706 37088
rect 10768 37036 10772 37088
rect 10849 37036 10874 37092
rect 10930 37036 10955 37092
rect 11011 37036 11036 37092
rect 11092 37036 11117 37092
rect 11173 37036 11198 37092
rect 11254 37088 11279 37092
rect 11335 37088 11360 37092
rect 11254 37036 11260 37088
rect 11416 37036 11441 37092
rect 12057 37088 13317 37103
rect 12057 37036 12368 37088
rect 12420 37036 12434 37088
rect 12486 37036 12922 37088
rect 12974 37036 12988 37088
rect 13040 37036 13317 37088
rect 2950 37030 13317 37036
rect 100 36992 2792 37004
rect 100 36940 2249 36992
rect 2301 36940 2315 36992
rect 2367 36940 2792 36992
rect 100 36928 2792 36940
rect 100 36876 2249 36928
rect 2301 36876 2315 36928
rect 2367 36876 2792 36928
rect 100 36864 2792 36876
rect 100 36812 2249 36864
rect 2301 36812 2315 36864
rect 2367 36812 2792 36864
rect 100 36800 2792 36812
rect 100 36748 2249 36800
rect 2301 36748 2315 36800
rect 2367 36748 2792 36800
rect 100 36736 2792 36748
rect 100 36684 2249 36736
rect 2301 36684 2315 36736
rect 2367 36726 2792 36736
tri 2792 36726 3002 36936 sw
rect 2367 36720 13602 36726
rect 2367 36684 3227 36720
rect 100 36672 3227 36684
rect 100 36620 2249 36672
rect 2301 36620 2315 36672
rect 2367 36668 3227 36672
rect 3279 36668 3293 36720
rect 3345 36668 3781 36720
rect 3833 36668 3847 36720
rect 3899 36668 4335 36720
rect 4387 36668 4401 36720
rect 4453 36668 4889 36720
rect 4941 36668 4955 36720
rect 5007 36668 5443 36720
rect 5495 36668 5509 36720
rect 5561 36668 5997 36720
rect 6049 36668 6063 36720
rect 6115 36668 6551 36720
rect 6603 36668 6617 36720
rect 6669 36668 7105 36720
rect 7157 36668 7171 36720
rect 7223 36668 7659 36720
rect 7711 36668 7725 36720
rect 7777 36668 8213 36720
rect 8265 36668 8279 36720
rect 8331 36668 8767 36720
rect 8819 36668 8833 36720
rect 8885 36668 9321 36720
rect 9373 36668 9387 36720
rect 9439 36668 9875 36720
rect 9927 36668 9941 36720
rect 9993 36668 10429 36720
rect 10481 36668 10495 36720
rect 10547 36668 10983 36720
rect 11035 36668 11049 36720
rect 11101 36668 11537 36720
rect 11589 36668 11603 36720
rect 11655 36668 12091 36720
rect 12143 36668 12157 36720
rect 12209 36668 12645 36720
rect 12697 36668 12711 36720
rect 12763 36668 13200 36720
rect 13252 36668 13270 36720
rect 13322 36668 13340 36720
rect 13392 36668 13410 36720
rect 13462 36668 13480 36720
rect 13532 36668 13550 36720
rect 2367 36654 13602 36668
rect 2367 36620 3227 36654
rect 100 36608 3227 36620
rect 100 36556 2249 36608
rect 2301 36556 2315 36608
rect 2367 36602 3227 36608
rect 3279 36602 3293 36654
rect 3345 36602 3781 36654
rect 3833 36602 3847 36654
rect 3899 36602 4335 36654
rect 4387 36602 4401 36654
rect 4453 36602 4889 36654
rect 4941 36602 4955 36654
rect 5007 36602 5443 36654
rect 5495 36602 5509 36654
rect 5561 36602 5997 36654
rect 6049 36602 6063 36654
rect 6115 36602 6551 36654
rect 6603 36602 6617 36654
rect 6669 36602 7105 36654
rect 7157 36602 7171 36654
rect 7223 36602 7659 36654
rect 7711 36602 7725 36654
rect 7777 36602 8213 36654
rect 8265 36602 8279 36654
rect 8331 36602 8767 36654
rect 8819 36602 8833 36654
rect 8885 36602 9321 36654
rect 9373 36602 9387 36654
rect 9439 36602 9875 36654
rect 9927 36602 9941 36654
rect 9993 36602 10429 36654
rect 10481 36602 10495 36654
rect 10547 36602 10983 36654
rect 11035 36602 11049 36654
rect 11101 36602 11537 36654
rect 11589 36602 11603 36654
rect 11655 36602 12091 36654
rect 12143 36602 12157 36654
rect 12209 36602 12645 36654
rect 12697 36602 12711 36654
rect 12763 36602 13200 36654
rect 13252 36602 13270 36654
rect 13322 36602 13340 36654
rect 13392 36602 13410 36654
rect 13462 36602 13480 36654
rect 13532 36602 13550 36654
rect 2367 36588 13602 36602
rect 2367 36556 3227 36588
rect 100 36544 3227 36556
rect 100 36492 2249 36544
rect 2301 36492 2315 36544
rect 2367 36536 3227 36544
rect 3279 36536 3293 36588
rect 3345 36536 3781 36588
rect 3833 36536 3847 36588
rect 3899 36536 4335 36588
rect 4387 36536 4401 36588
rect 4453 36536 4889 36588
rect 4941 36536 4955 36588
rect 5007 36536 5443 36588
rect 5495 36536 5509 36588
rect 5561 36536 5997 36588
rect 6049 36536 6063 36588
rect 6115 36536 6551 36588
rect 6603 36536 6617 36588
rect 6669 36536 7105 36588
rect 7157 36536 7171 36588
rect 7223 36536 7659 36588
rect 7711 36536 7725 36588
rect 7777 36536 8213 36588
rect 8265 36536 8279 36588
rect 8331 36536 8767 36588
rect 8819 36536 8833 36588
rect 8885 36536 9321 36588
rect 9373 36536 9387 36588
rect 9439 36536 9875 36588
rect 9927 36536 9941 36588
rect 9993 36536 10429 36588
rect 10481 36536 10495 36588
rect 10547 36536 10983 36588
rect 11035 36536 11049 36588
rect 11101 36536 11537 36588
rect 11589 36536 11603 36588
rect 11655 36536 12091 36588
rect 12143 36536 12157 36588
rect 12209 36536 12645 36588
rect 12697 36536 12711 36588
rect 12763 36536 13200 36588
rect 13252 36536 13270 36588
rect 13322 36536 13340 36588
rect 13392 36536 13410 36588
rect 13462 36536 13480 36588
rect 13532 36536 13550 36588
rect 2367 36522 13602 36536
rect 2367 36492 3227 36522
rect 100 36480 3227 36492
rect 100 36428 2249 36480
rect 2301 36428 2315 36480
rect 2367 36470 3227 36480
rect 3279 36470 3293 36522
rect 3345 36470 3781 36522
rect 3833 36470 3847 36522
rect 3899 36470 4335 36522
rect 4387 36470 4401 36522
rect 4453 36470 4889 36522
rect 4941 36470 4955 36522
rect 5007 36470 5443 36522
rect 5495 36470 5509 36522
rect 5561 36470 5997 36522
rect 6049 36470 6063 36522
rect 6115 36470 6551 36522
rect 6603 36470 6617 36522
rect 6669 36470 7105 36522
rect 7157 36470 7171 36522
rect 7223 36470 7659 36522
rect 7711 36470 7725 36522
rect 7777 36470 8213 36522
rect 8265 36470 8279 36522
rect 8331 36470 8767 36522
rect 8819 36470 8833 36522
rect 8885 36470 9321 36522
rect 9373 36470 9387 36522
rect 9439 36470 9875 36522
rect 9927 36470 9941 36522
rect 9993 36470 10429 36522
rect 10481 36470 10495 36522
rect 10547 36470 10983 36522
rect 11035 36470 11049 36522
rect 11101 36470 11537 36522
rect 11589 36470 11603 36522
rect 11655 36470 12091 36522
rect 12143 36470 12157 36522
rect 12209 36470 12645 36522
rect 12697 36470 12711 36522
rect 12763 36470 13200 36522
rect 13252 36470 13270 36522
rect 13322 36470 13340 36522
rect 13392 36470 13410 36522
rect 13462 36470 13480 36522
rect 13532 36470 13550 36522
rect 2367 36456 13602 36470
rect 2367 36428 3227 36456
rect 100 36416 3227 36428
rect 100 36364 2249 36416
rect 2301 36364 2315 36416
rect 2367 36404 3227 36416
rect 3279 36404 3293 36456
rect 3345 36404 3781 36456
rect 3833 36404 3847 36456
rect 3899 36404 4335 36456
rect 4387 36404 4401 36456
rect 4453 36404 4889 36456
rect 4941 36404 4955 36456
rect 5007 36404 5443 36456
rect 5495 36404 5509 36456
rect 5561 36404 5997 36456
rect 6049 36404 6063 36456
rect 6115 36404 6551 36456
rect 6603 36404 6617 36456
rect 6669 36404 7105 36456
rect 7157 36404 7171 36456
rect 7223 36404 7659 36456
rect 7711 36404 7725 36456
rect 7777 36404 8213 36456
rect 8265 36404 8279 36456
rect 8331 36404 8767 36456
rect 8819 36404 8833 36456
rect 8885 36404 9321 36456
rect 9373 36404 9387 36456
rect 9439 36404 9875 36456
rect 9927 36404 9941 36456
rect 9993 36404 10429 36456
rect 10481 36404 10495 36456
rect 10547 36404 10983 36456
rect 11035 36404 11049 36456
rect 11101 36404 11537 36456
rect 11589 36404 11603 36456
rect 11655 36404 12091 36456
rect 12143 36404 12157 36456
rect 12209 36404 12645 36456
rect 12697 36404 12711 36456
rect 12763 36404 13200 36456
rect 13252 36404 13270 36456
rect 13322 36404 13340 36456
rect 13392 36404 13410 36456
rect 13462 36404 13480 36456
rect 13532 36404 13550 36456
rect 2367 36390 13602 36404
rect 2367 36364 3227 36390
rect 100 36352 3227 36364
rect 100 36300 2249 36352
rect 2301 36300 2315 36352
rect 2367 36338 3227 36352
rect 3279 36338 3293 36390
rect 3345 36338 3781 36390
rect 3833 36338 3847 36390
rect 3899 36338 4335 36390
rect 4387 36338 4401 36390
rect 4453 36338 4889 36390
rect 4941 36338 4955 36390
rect 5007 36338 5443 36390
rect 5495 36338 5509 36390
rect 5561 36338 5997 36390
rect 6049 36338 6063 36390
rect 6115 36338 6551 36390
rect 6603 36338 6617 36390
rect 6669 36338 7105 36390
rect 7157 36338 7171 36390
rect 7223 36338 7659 36390
rect 7711 36338 7725 36390
rect 7777 36338 8213 36390
rect 8265 36338 8279 36390
rect 8331 36338 8767 36390
rect 8819 36338 8833 36390
rect 8885 36338 9321 36390
rect 9373 36338 9387 36390
rect 9439 36338 9875 36390
rect 9927 36338 9941 36390
rect 9993 36338 10429 36390
rect 10481 36338 10495 36390
rect 10547 36338 10983 36390
rect 11035 36338 11049 36390
rect 11101 36338 11537 36390
rect 11589 36338 11603 36390
rect 11655 36338 12091 36390
rect 12143 36338 12157 36390
rect 12209 36338 12645 36390
rect 12697 36338 12711 36390
rect 12763 36338 13200 36390
rect 13252 36338 13270 36390
rect 13322 36338 13340 36390
rect 13392 36338 13410 36390
rect 13462 36338 13480 36390
rect 13532 36338 13550 36390
rect 2367 36323 13602 36338
rect 2367 36300 3227 36323
rect 100 36288 3227 36300
rect 100 36236 2249 36288
rect 2301 36236 2315 36288
rect 2367 36271 3227 36288
rect 3279 36271 3293 36323
rect 3345 36271 3781 36323
rect 3833 36271 3847 36323
rect 3899 36271 4335 36323
rect 4387 36271 4401 36323
rect 4453 36271 4889 36323
rect 4941 36271 4955 36323
rect 5007 36271 5443 36323
rect 5495 36271 5509 36323
rect 5561 36271 5997 36323
rect 6049 36271 6063 36323
rect 6115 36271 6551 36323
rect 6603 36271 6617 36323
rect 6669 36271 7105 36323
rect 7157 36271 7171 36323
rect 7223 36271 7659 36323
rect 7711 36271 7725 36323
rect 7777 36271 8213 36323
rect 8265 36271 8279 36323
rect 8331 36271 8767 36323
rect 8819 36271 8833 36323
rect 8885 36271 9321 36323
rect 9373 36271 9387 36323
rect 9439 36271 9875 36323
rect 9927 36271 9941 36323
rect 9993 36271 10429 36323
rect 10481 36271 10495 36323
rect 10547 36271 10983 36323
rect 11035 36271 11049 36323
rect 11101 36271 11537 36323
rect 11589 36271 11603 36323
rect 11655 36271 12091 36323
rect 12143 36271 12157 36323
rect 12209 36271 12645 36323
rect 12697 36271 12711 36323
rect 12763 36271 13200 36323
rect 13252 36271 13270 36323
rect 13322 36271 13340 36323
rect 13392 36271 13410 36323
rect 13462 36271 13480 36323
rect 13532 36271 13550 36323
rect 2367 36256 13602 36271
rect 2367 36236 3227 36256
rect 100 36224 3227 36236
rect 100 36172 2249 36224
rect 2301 36172 2315 36224
rect 2367 36204 3227 36224
rect 3279 36204 3293 36256
rect 3345 36204 3781 36256
rect 3833 36204 3847 36256
rect 3899 36204 4335 36256
rect 4387 36204 4401 36256
rect 4453 36204 4889 36256
rect 4941 36204 4955 36256
rect 5007 36204 5443 36256
rect 5495 36204 5509 36256
rect 5561 36204 5997 36256
rect 6049 36204 6063 36256
rect 6115 36204 6551 36256
rect 6603 36204 6617 36256
rect 6669 36204 7105 36256
rect 7157 36204 7171 36256
rect 7223 36204 7659 36256
rect 7711 36204 7725 36256
rect 7777 36204 8213 36256
rect 8265 36204 8279 36256
rect 8331 36204 8767 36256
rect 8819 36204 8833 36256
rect 8885 36204 9321 36256
rect 9373 36204 9387 36256
rect 9439 36204 9875 36256
rect 9927 36204 9941 36256
rect 9993 36204 10429 36256
rect 10481 36204 10495 36256
rect 10547 36204 10983 36256
rect 11035 36204 11049 36256
rect 11101 36204 11537 36256
rect 11589 36204 11603 36256
rect 11655 36204 12091 36256
rect 12143 36204 12157 36256
rect 12209 36204 12645 36256
rect 12697 36204 12711 36256
rect 12763 36204 13200 36256
rect 13252 36204 13270 36256
rect 13322 36204 13340 36256
rect 13392 36204 13410 36256
rect 13462 36204 13480 36256
rect 13532 36204 13550 36256
rect 2367 36198 13602 36204
rect 2367 36172 2792 36198
rect 100 36160 2792 36172
rect 100 36108 2249 36160
rect 2301 36108 2315 36160
rect 2367 36108 2792 36160
rect 100 36096 2792 36108
rect 100 36044 2249 36096
rect 2301 36044 2315 36096
rect 2367 36044 2792 36096
rect 100 36032 2792 36044
rect 100 35980 2249 36032
rect 2301 35980 2315 36032
rect 2367 35980 2792 36032
tri 2792 35988 3002 36198 nw
rect 100 35968 2792 35980
rect 100 35916 2249 35968
rect 2301 35916 2315 35968
rect 2367 35916 2792 35968
rect 100 35904 2792 35916
rect 100 35852 2249 35904
rect 2301 35852 2315 35904
rect 2367 35852 2792 35904
rect 100 35840 2792 35852
rect 100 35788 2249 35840
rect 2301 35788 2315 35840
rect 2367 35788 2792 35840
rect 100 35776 2792 35788
rect 100 35724 2249 35776
rect 2301 35724 2315 35776
rect 2367 35724 2792 35776
rect 100 35712 2792 35724
rect 100 35660 2249 35712
rect 2301 35660 2315 35712
rect 2367 35660 2792 35712
rect 100 35648 2792 35660
rect 100 35596 2249 35648
rect 2301 35596 2315 35648
rect 2367 35596 2792 35648
rect 100 35584 2792 35596
rect 100 35532 2249 35584
rect 2301 35532 2315 35584
rect 2367 35532 2792 35584
rect 100 35520 2792 35532
rect 100 35468 2249 35520
rect 2301 35468 2315 35520
rect 2367 35468 2792 35520
rect 100 35456 2792 35468
rect 100 35404 2249 35456
rect 2301 35404 2315 35456
rect 2367 35404 2792 35456
rect 100 35392 2792 35404
rect 100 35340 2249 35392
rect 2301 35340 2315 35392
rect 2367 35340 2792 35392
rect 3504 35896 13317 35898
rect 3504 35892 3513 35896
rect 3569 35892 3593 35896
rect 3569 35840 3570 35892
rect 3649 35840 3673 35896
rect 3729 35840 3753 35896
rect 3809 35840 3833 35896
rect 3889 35840 3913 35896
rect 3969 35840 3993 35896
rect 4049 35892 4073 35896
rect 4129 35892 4153 35896
rect 4049 35840 4058 35892
rect 4209 35840 4233 35896
rect 4289 35840 4314 35896
rect 4370 35840 4395 35896
rect 4451 35840 4476 35896
rect 4532 35840 4557 35896
rect 4613 35892 4638 35896
rect 4694 35892 4719 35896
rect 4775 35840 4800 35896
rect 4856 35840 4881 35896
rect 4937 35840 4962 35896
rect 5018 35892 13317 35896
rect 5018 35840 5166 35892
rect 5218 35877 5232 35892
rect 5284 35877 5720 35892
rect 5772 35877 5786 35892
rect 5838 35877 6274 35892
rect 5284 35840 5296 35877
rect 3504 35826 5215 35840
rect 5271 35826 5296 35840
rect 3556 35802 3570 35826
rect 3622 35802 4058 35826
rect 4110 35802 4124 35826
rect 4176 35802 4612 35826
rect 4664 35802 4678 35826
rect 4730 35802 5166 35826
rect 5284 35821 5296 35826
rect 5352 35821 5377 35877
rect 5433 35821 5458 35877
rect 5514 35821 5539 35877
rect 5595 35821 5620 35877
rect 5676 35821 5701 35877
rect 5772 35840 5782 35877
rect 5757 35826 5782 35840
rect 5772 35821 5782 35826
rect 5838 35821 5863 35877
rect 5919 35821 5944 35877
rect 6000 35821 6025 35877
rect 6081 35821 6106 35877
rect 6162 35821 6187 35877
rect 6243 35821 6268 35877
rect 6326 35840 6340 35892
rect 6392 35877 6828 35892
rect 6880 35877 6894 35892
rect 6946 35877 7382 35892
rect 6324 35826 6349 35840
rect 3569 35774 3570 35802
rect 3504 35760 3513 35774
rect 3569 35760 3593 35774
rect 3569 35746 3570 35760
rect 3649 35746 3673 35802
rect 3729 35746 3753 35802
rect 3809 35746 3833 35802
rect 3889 35746 3913 35802
rect 3969 35746 3993 35802
rect 4049 35774 4058 35802
rect 4049 35760 4073 35774
rect 4129 35760 4153 35774
rect 4049 35746 4058 35760
rect 4209 35746 4233 35802
rect 4289 35746 4314 35802
rect 4370 35746 4395 35802
rect 4451 35746 4476 35802
rect 4532 35746 4557 35802
rect 4613 35760 4638 35774
rect 4694 35760 4719 35774
rect 4775 35746 4800 35802
rect 4856 35746 4881 35802
rect 4937 35746 4962 35802
rect 5018 35774 5166 35802
rect 5218 35789 5232 35821
rect 5284 35789 5720 35821
rect 5772 35789 5786 35821
rect 5838 35789 6274 35821
rect 5284 35774 5296 35789
rect 5018 35760 5215 35774
rect 5271 35760 5296 35774
rect 5018 35746 5166 35760
rect 3556 35708 3570 35746
rect 3622 35708 4058 35746
rect 4110 35708 4124 35746
rect 4176 35708 4612 35746
rect 4664 35708 4678 35746
rect 4730 35708 5166 35746
rect 5284 35733 5296 35760
rect 5352 35733 5377 35789
rect 5433 35733 5458 35789
rect 5514 35733 5539 35789
rect 5595 35733 5620 35789
rect 5676 35733 5701 35789
rect 5772 35774 5782 35789
rect 5757 35760 5782 35774
rect 5772 35733 5782 35760
rect 5838 35733 5863 35789
rect 5919 35733 5944 35789
rect 6000 35733 6025 35789
rect 6081 35733 6106 35789
rect 6162 35733 6187 35789
rect 6243 35733 6268 35789
rect 6326 35774 6340 35826
rect 6405 35821 6430 35877
rect 6486 35821 6511 35877
rect 6567 35821 6592 35877
rect 6648 35821 6673 35877
rect 6729 35821 6754 35877
rect 6810 35840 6828 35877
rect 6891 35840 6894 35877
rect 6810 35826 6835 35840
rect 6891 35826 6916 35840
rect 6810 35821 6828 35826
rect 6891 35821 6894 35826
rect 6972 35821 6997 35877
rect 7053 35821 7078 35877
rect 7134 35821 7159 35877
rect 7215 35821 7240 35877
rect 7296 35821 7320 35877
rect 7376 35840 7382 35877
rect 7434 35840 7448 35892
rect 7500 35877 7936 35892
rect 7500 35840 7598 35877
rect 7376 35826 7598 35840
rect 7376 35821 7382 35826
rect 6392 35789 6828 35821
rect 6880 35789 6894 35821
rect 6946 35789 7382 35821
rect 6324 35760 6349 35774
rect 5218 35708 5232 35733
rect 5284 35708 5720 35733
rect 5772 35708 5786 35733
rect 5838 35708 6274 35733
rect 6326 35708 6340 35760
rect 6405 35733 6430 35789
rect 6486 35733 6511 35789
rect 6567 35733 6592 35789
rect 6648 35733 6673 35789
rect 6729 35733 6754 35789
rect 6810 35774 6828 35789
rect 6891 35774 6894 35789
rect 6810 35760 6835 35774
rect 6891 35760 6916 35774
rect 6810 35733 6828 35760
rect 6891 35733 6894 35760
rect 6972 35733 6997 35789
rect 7053 35733 7078 35789
rect 7134 35733 7159 35789
rect 7215 35733 7240 35789
rect 7296 35733 7320 35789
rect 7376 35774 7382 35789
rect 7434 35774 7448 35826
rect 7500 35821 7598 35826
rect 7654 35821 7678 35877
rect 7734 35821 7759 35877
rect 7815 35821 7840 35877
rect 7896 35821 7921 35877
rect 7988 35840 8002 35892
rect 8054 35877 8490 35892
rect 8542 35877 8556 35892
rect 8608 35877 9044 35892
rect 9096 35877 9110 35892
rect 9162 35877 9598 35892
rect 9650 35877 9664 35892
rect 9716 35877 10152 35892
rect 7977 35826 8002 35840
rect 7500 35789 7936 35821
rect 7500 35774 7598 35789
rect 7376 35760 7598 35774
rect 7376 35733 7382 35760
rect 6392 35708 6828 35733
rect 6880 35708 6894 35733
rect 6946 35708 7382 35733
rect 7434 35708 7448 35760
rect 7500 35733 7598 35760
rect 7654 35733 7678 35789
rect 7734 35733 7759 35789
rect 7815 35733 7840 35789
rect 7896 35733 7921 35789
rect 7988 35774 8002 35826
rect 8058 35821 8083 35877
rect 8139 35821 8164 35877
rect 8220 35821 8245 35877
rect 8301 35821 8326 35877
rect 8382 35821 8407 35877
rect 8463 35821 8488 35877
rect 8544 35840 8556 35877
rect 8544 35826 8569 35840
rect 8544 35821 8556 35826
rect 8625 35821 8650 35877
rect 8706 35821 8731 35877
rect 8787 35821 8812 35877
rect 8868 35821 8893 35877
rect 8949 35821 8974 35877
rect 9030 35840 9044 35877
rect 9030 35826 9055 35840
rect 9111 35826 9136 35840
rect 9030 35821 9044 35826
rect 9192 35821 9217 35877
rect 9273 35821 9298 35877
rect 9354 35821 9379 35877
rect 9435 35821 9460 35877
rect 9516 35821 9541 35877
rect 9597 35840 9598 35877
rect 9597 35826 9622 35840
rect 9678 35826 9703 35840
rect 9597 35821 9598 35826
rect 9759 35821 9983 35877
rect 10039 35821 10063 35877
rect 10119 35821 10143 35877
rect 10204 35840 10218 35892
rect 10270 35877 10706 35892
rect 10758 35877 10772 35892
rect 10824 35877 11260 35892
rect 11312 35877 11326 35892
rect 11378 35877 11814 35892
rect 11866 35877 11880 35892
rect 11932 35877 12368 35892
rect 10199 35826 10223 35840
rect 8054 35789 8490 35821
rect 8542 35789 8556 35821
rect 8608 35789 9044 35821
rect 9096 35789 9110 35821
rect 9162 35789 9598 35821
rect 9650 35789 9664 35821
rect 9716 35789 10152 35821
rect 7977 35760 8002 35774
rect 7500 35708 7936 35733
rect 7988 35708 8002 35760
rect 8058 35733 8083 35789
rect 8139 35733 8164 35789
rect 8220 35733 8245 35789
rect 8301 35733 8326 35789
rect 8382 35733 8407 35789
rect 8463 35733 8488 35789
rect 8544 35774 8556 35789
rect 8544 35760 8569 35774
rect 8544 35733 8556 35760
rect 8625 35733 8650 35789
rect 8706 35733 8731 35789
rect 8787 35733 8812 35789
rect 8868 35733 8893 35789
rect 8949 35733 8974 35789
rect 9030 35774 9044 35789
rect 9030 35760 9055 35774
rect 9111 35760 9136 35774
rect 9030 35733 9044 35760
rect 9192 35733 9217 35789
rect 9273 35733 9298 35789
rect 9354 35733 9379 35789
rect 9435 35733 9460 35789
rect 9516 35733 9541 35789
rect 9597 35774 9598 35789
rect 9597 35760 9622 35774
rect 9678 35760 9703 35774
rect 9597 35733 9598 35760
rect 9759 35733 9983 35789
rect 10039 35733 10063 35789
rect 10119 35733 10143 35789
rect 10204 35774 10218 35826
rect 10279 35821 10303 35877
rect 10359 35821 10383 35877
rect 10439 35821 10463 35877
rect 10519 35821 10544 35877
rect 10600 35821 10625 35877
rect 10681 35821 10706 35877
rect 10762 35840 10772 35877
rect 10762 35826 10787 35840
rect 10762 35821 10772 35826
rect 10843 35821 10868 35877
rect 10924 35821 10949 35877
rect 11005 35821 11030 35877
rect 11086 35821 11111 35877
rect 11167 35821 11192 35877
rect 11248 35840 11260 35877
rect 11248 35826 11273 35840
rect 11329 35826 11354 35840
rect 11248 35821 11260 35826
rect 11410 35821 11435 35877
rect 11491 35821 11516 35877
rect 11572 35821 11597 35877
rect 11653 35821 11678 35877
rect 11734 35821 11759 35877
rect 11815 35826 11840 35840
rect 11896 35826 11921 35840
rect 11977 35821 12002 35877
rect 12058 35840 12368 35877
rect 12420 35840 12434 35892
rect 12486 35840 12922 35892
rect 12974 35840 12988 35892
rect 13040 35840 13317 35892
rect 12058 35826 13317 35840
rect 12058 35821 12368 35826
rect 10270 35789 10706 35821
rect 10758 35789 10772 35821
rect 10824 35789 11260 35821
rect 11312 35789 11326 35821
rect 11378 35789 11814 35821
rect 11866 35789 11880 35821
rect 11932 35789 12368 35821
rect 10199 35760 10223 35774
rect 8054 35708 8490 35733
rect 8542 35708 8556 35733
rect 8608 35708 9044 35733
rect 9096 35708 9110 35733
rect 9162 35708 9598 35733
rect 9650 35708 9664 35733
rect 9716 35708 10152 35733
rect 10204 35708 10218 35760
rect 10279 35733 10303 35789
rect 10359 35733 10383 35789
rect 10439 35733 10463 35789
rect 10519 35733 10544 35789
rect 10600 35733 10625 35789
rect 10681 35733 10706 35789
rect 10762 35774 10772 35789
rect 10762 35760 10787 35774
rect 10762 35733 10772 35760
rect 10843 35733 10868 35789
rect 10924 35733 10949 35789
rect 11005 35733 11030 35789
rect 11086 35733 11111 35789
rect 11167 35733 11192 35789
rect 11248 35774 11260 35789
rect 11248 35760 11273 35774
rect 11329 35760 11354 35774
rect 11248 35733 11260 35760
rect 11410 35733 11435 35789
rect 11491 35733 11516 35789
rect 11572 35733 11597 35789
rect 11653 35733 11678 35789
rect 11734 35733 11759 35789
rect 11815 35760 11840 35774
rect 11896 35760 11921 35774
rect 11977 35733 12002 35789
rect 12058 35774 12368 35789
rect 12420 35774 12434 35826
rect 12486 35774 12922 35826
rect 12974 35774 12988 35826
rect 13040 35774 13317 35826
rect 12058 35760 13317 35774
rect 12058 35733 12368 35760
rect 10270 35708 10706 35733
rect 10758 35708 10772 35733
rect 10824 35708 11260 35733
rect 11312 35708 11326 35733
rect 11378 35708 11814 35733
rect 11866 35708 11880 35733
rect 11932 35708 12368 35733
rect 12420 35708 12434 35760
rect 12486 35708 12922 35760
rect 12974 35708 12988 35760
rect 13040 35708 13317 35760
rect 3504 35694 3513 35708
rect 3569 35694 3593 35708
rect 3569 35652 3570 35694
rect 3649 35652 3673 35708
rect 3729 35652 3753 35708
rect 3809 35652 3833 35708
rect 3889 35652 3913 35708
rect 3969 35652 3993 35708
rect 4049 35694 4073 35708
rect 4129 35694 4153 35708
rect 4049 35652 4058 35694
rect 4209 35652 4233 35708
rect 4289 35652 4314 35708
rect 4370 35652 4395 35708
rect 4451 35652 4476 35708
rect 4532 35652 4557 35708
rect 4613 35694 4638 35708
rect 4694 35694 4719 35708
rect 4775 35652 4800 35708
rect 4856 35652 4881 35708
rect 4937 35652 4962 35708
rect 5018 35701 13317 35708
rect 5018 35694 5215 35701
rect 5271 35694 5296 35701
rect 5018 35652 5166 35694
rect 3556 35642 3570 35652
rect 3622 35642 4058 35652
rect 4110 35642 4124 35652
rect 4176 35642 4612 35652
rect 4664 35642 4678 35652
rect 4730 35642 5166 35652
rect 5284 35645 5296 35694
rect 5352 35645 5377 35701
rect 5433 35645 5458 35701
rect 5514 35645 5539 35701
rect 5595 35645 5620 35701
rect 5676 35645 5701 35701
rect 5757 35694 5782 35701
rect 5772 35645 5782 35694
rect 5838 35645 5863 35701
rect 5919 35645 5944 35701
rect 6000 35645 6025 35701
rect 6081 35645 6106 35701
rect 6162 35645 6187 35701
rect 6243 35645 6268 35701
rect 6324 35694 6349 35701
rect 5218 35642 5232 35645
rect 5284 35642 5720 35645
rect 5772 35642 5786 35645
rect 5838 35642 6274 35645
rect 6326 35642 6340 35694
rect 6405 35645 6430 35701
rect 6486 35645 6511 35701
rect 6567 35645 6592 35701
rect 6648 35645 6673 35701
rect 6729 35645 6754 35701
rect 6810 35694 6835 35701
rect 6891 35694 6916 35701
rect 6810 35645 6828 35694
rect 6891 35645 6894 35694
rect 6972 35645 6997 35701
rect 7053 35645 7078 35701
rect 7134 35645 7159 35701
rect 7215 35645 7240 35701
rect 7296 35645 7320 35701
rect 7376 35694 7598 35701
rect 7376 35645 7382 35694
rect 6392 35642 6828 35645
rect 6880 35642 6894 35645
rect 6946 35642 7382 35645
rect 7434 35642 7448 35694
rect 7500 35645 7598 35694
rect 7654 35645 7678 35701
rect 7734 35645 7759 35701
rect 7815 35645 7840 35701
rect 7896 35645 7921 35701
rect 7977 35694 8002 35701
rect 7500 35642 7936 35645
rect 7988 35642 8002 35694
rect 8058 35645 8083 35701
rect 8139 35645 8164 35701
rect 8220 35645 8245 35701
rect 8301 35645 8326 35701
rect 8382 35645 8407 35701
rect 8463 35645 8488 35701
rect 8544 35694 8569 35701
rect 8544 35645 8556 35694
rect 8625 35645 8650 35701
rect 8706 35645 8731 35701
rect 8787 35645 8812 35701
rect 8868 35645 8893 35701
rect 8949 35645 8974 35701
rect 9030 35694 9055 35701
rect 9111 35694 9136 35701
rect 9030 35645 9044 35694
rect 9192 35645 9217 35701
rect 9273 35645 9298 35701
rect 9354 35645 9379 35701
rect 9435 35645 9460 35701
rect 9516 35645 9541 35701
rect 9597 35694 9622 35701
rect 9678 35694 9703 35701
rect 9597 35645 9598 35694
rect 9759 35645 9983 35701
rect 10039 35645 10063 35701
rect 10119 35645 10143 35701
rect 10199 35694 10223 35701
rect 8054 35642 8490 35645
rect 8542 35642 8556 35645
rect 8608 35642 9044 35645
rect 9096 35642 9110 35645
rect 9162 35642 9598 35645
rect 9650 35642 9664 35645
rect 9716 35642 10152 35645
rect 10204 35642 10218 35694
rect 10279 35645 10303 35701
rect 10359 35645 10383 35701
rect 10439 35645 10463 35701
rect 10519 35645 10544 35701
rect 10600 35645 10625 35701
rect 10681 35645 10706 35701
rect 10762 35694 10787 35701
rect 10762 35645 10772 35694
rect 10843 35645 10868 35701
rect 10924 35645 10949 35701
rect 11005 35645 11030 35701
rect 11086 35645 11111 35701
rect 11167 35645 11192 35701
rect 11248 35694 11273 35701
rect 11329 35694 11354 35701
rect 11248 35645 11260 35694
rect 11410 35645 11435 35701
rect 11491 35645 11516 35701
rect 11572 35645 11597 35701
rect 11653 35645 11678 35701
rect 11734 35645 11759 35701
rect 11815 35694 11840 35701
rect 11896 35694 11921 35701
rect 11977 35645 12002 35701
rect 12058 35694 13317 35701
rect 12058 35645 12368 35694
rect 10270 35642 10706 35645
rect 10758 35642 10772 35645
rect 10824 35642 11260 35645
rect 11312 35642 11326 35645
rect 11378 35642 11814 35645
rect 11866 35642 11880 35645
rect 11932 35642 12368 35645
rect 12420 35642 12434 35694
rect 12486 35642 12922 35694
rect 12974 35642 12988 35694
rect 13040 35642 13317 35694
rect 3504 35627 13317 35642
rect 3556 35614 3570 35627
rect 3622 35614 4058 35627
rect 4110 35614 4124 35627
rect 4176 35614 4612 35627
rect 4664 35614 4678 35627
rect 4730 35614 5166 35627
rect 3569 35575 3570 35614
rect 3504 35560 3513 35575
rect 3569 35560 3593 35575
rect 3569 35558 3570 35560
rect 3649 35558 3673 35614
rect 3729 35558 3753 35614
rect 3809 35558 3833 35614
rect 3889 35558 3913 35614
rect 3969 35558 3993 35614
rect 4049 35575 4058 35614
rect 4049 35560 4073 35575
rect 4129 35560 4153 35575
rect 4049 35558 4058 35560
rect 4209 35558 4233 35614
rect 4289 35558 4314 35614
rect 4370 35558 4395 35614
rect 4451 35558 4476 35614
rect 4532 35558 4557 35614
rect 4613 35560 4638 35575
rect 4694 35560 4719 35575
rect 4775 35558 4800 35614
rect 4856 35558 4881 35614
rect 4937 35558 4962 35614
rect 5018 35575 5166 35614
rect 5218 35613 5232 35627
rect 5284 35613 5720 35627
rect 5772 35613 5786 35627
rect 5838 35613 6274 35627
rect 5284 35575 5296 35613
rect 5018 35560 5215 35575
rect 5271 35560 5296 35575
rect 5018 35558 5166 35560
rect 3556 35520 3570 35558
rect 3622 35520 4058 35558
rect 4110 35520 4124 35558
rect 4176 35520 4612 35558
rect 4664 35520 4678 35558
rect 4730 35520 5166 35558
rect 5284 35557 5296 35560
rect 5352 35557 5377 35613
rect 5433 35557 5458 35613
rect 5514 35557 5539 35613
rect 5595 35557 5620 35613
rect 5676 35557 5701 35613
rect 5772 35575 5782 35613
rect 5757 35560 5782 35575
rect 5772 35557 5782 35560
rect 5838 35557 5863 35613
rect 5919 35557 5944 35613
rect 6000 35557 6025 35613
rect 6081 35557 6106 35613
rect 6162 35557 6187 35613
rect 6243 35557 6268 35613
rect 6326 35575 6340 35627
rect 6392 35613 6828 35627
rect 6880 35613 6894 35627
rect 6946 35613 7382 35627
rect 6324 35560 6349 35575
rect 5218 35525 5232 35557
rect 5284 35525 5720 35557
rect 5772 35525 5786 35557
rect 5838 35525 6274 35557
rect 3569 35508 3570 35520
rect 3504 35493 3513 35508
rect 3569 35493 3593 35508
rect 3569 35464 3570 35493
rect 3649 35464 3673 35520
rect 3729 35464 3753 35520
rect 3809 35464 3833 35520
rect 3889 35464 3913 35520
rect 3969 35464 3993 35520
rect 4049 35508 4058 35520
rect 4049 35493 4073 35508
rect 4129 35493 4153 35508
rect 4049 35464 4058 35493
rect 4209 35464 4233 35520
rect 4289 35464 4314 35520
rect 4370 35464 4395 35520
rect 4451 35464 4476 35520
rect 4532 35464 4557 35520
rect 4613 35493 4638 35508
rect 4694 35493 4719 35508
rect 4775 35464 4800 35520
rect 4856 35464 4881 35520
rect 4937 35464 4962 35520
rect 5018 35508 5166 35520
rect 5284 35508 5296 35525
rect 5018 35493 5215 35508
rect 5271 35493 5296 35508
rect 5018 35464 5166 35493
rect 5284 35469 5296 35493
rect 5352 35469 5377 35525
rect 5433 35469 5458 35525
rect 5514 35469 5539 35525
rect 5595 35469 5620 35525
rect 5676 35469 5701 35525
rect 5772 35508 5782 35525
rect 5757 35493 5782 35508
rect 5772 35469 5782 35493
rect 5838 35469 5863 35525
rect 5919 35469 5944 35525
rect 6000 35469 6025 35525
rect 6081 35469 6106 35525
rect 6162 35469 6187 35525
rect 6243 35469 6268 35525
rect 6326 35508 6340 35560
rect 6405 35557 6430 35613
rect 6486 35557 6511 35613
rect 6567 35557 6592 35613
rect 6648 35557 6673 35613
rect 6729 35557 6754 35613
rect 6810 35575 6828 35613
rect 6891 35575 6894 35613
rect 6810 35560 6835 35575
rect 6891 35560 6916 35575
rect 6810 35557 6828 35560
rect 6891 35557 6894 35560
rect 6972 35557 6997 35613
rect 7053 35557 7078 35613
rect 7134 35557 7159 35613
rect 7215 35557 7240 35613
rect 7296 35557 7320 35613
rect 7376 35575 7382 35613
rect 7434 35575 7448 35627
rect 7500 35613 7936 35627
rect 7500 35575 7598 35613
rect 7376 35560 7598 35575
rect 7376 35557 7382 35560
rect 6392 35525 6828 35557
rect 6880 35525 6894 35557
rect 6946 35525 7382 35557
rect 6324 35493 6349 35508
rect 3556 35441 3570 35464
rect 3622 35441 4058 35464
rect 4110 35441 4124 35464
rect 4176 35441 4612 35464
rect 4664 35441 4678 35464
rect 4730 35441 5166 35464
rect 5218 35441 5232 35469
rect 5284 35441 5720 35469
rect 5772 35441 5786 35469
rect 5838 35441 6274 35469
rect 6326 35441 6340 35493
rect 6405 35469 6430 35525
rect 6486 35469 6511 35525
rect 6567 35469 6592 35525
rect 6648 35469 6673 35525
rect 6729 35469 6754 35525
rect 6810 35508 6828 35525
rect 6891 35508 6894 35525
rect 6810 35493 6835 35508
rect 6891 35493 6916 35508
rect 6810 35469 6828 35493
rect 6891 35469 6894 35493
rect 6972 35469 6997 35525
rect 7053 35469 7078 35525
rect 7134 35469 7159 35525
rect 7215 35469 7240 35525
rect 7296 35469 7320 35525
rect 7376 35508 7382 35525
rect 7434 35508 7448 35560
rect 7500 35557 7598 35560
rect 7654 35557 7678 35613
rect 7734 35557 7759 35613
rect 7815 35557 7840 35613
rect 7896 35557 7921 35613
rect 7988 35575 8002 35627
rect 8054 35613 8490 35627
rect 8542 35613 8556 35627
rect 8608 35613 9044 35627
rect 9096 35613 9110 35627
rect 9162 35613 9598 35627
rect 9650 35613 9664 35627
rect 9716 35613 10152 35627
rect 7977 35560 8002 35575
rect 7500 35525 7936 35557
rect 7500 35508 7598 35525
rect 7376 35493 7598 35508
rect 7376 35469 7382 35493
rect 6392 35441 6828 35469
rect 6880 35441 6894 35469
rect 6946 35441 7382 35469
rect 7434 35441 7448 35493
rect 7500 35469 7598 35493
rect 7654 35469 7678 35525
rect 7734 35469 7759 35525
rect 7815 35469 7840 35525
rect 7896 35469 7921 35525
rect 7988 35508 8002 35560
rect 8058 35557 8083 35613
rect 8139 35557 8164 35613
rect 8220 35557 8245 35613
rect 8301 35557 8326 35613
rect 8382 35557 8407 35613
rect 8463 35557 8488 35613
rect 8544 35575 8556 35613
rect 8544 35560 8569 35575
rect 8544 35557 8556 35560
rect 8625 35557 8650 35613
rect 8706 35557 8731 35613
rect 8787 35557 8812 35613
rect 8868 35557 8893 35613
rect 8949 35557 8974 35613
rect 9030 35575 9044 35613
rect 9030 35560 9055 35575
rect 9111 35560 9136 35575
rect 9030 35557 9044 35560
rect 9192 35557 9217 35613
rect 9273 35557 9298 35613
rect 9354 35557 9379 35613
rect 9435 35557 9460 35613
rect 9516 35557 9541 35613
rect 9597 35575 9598 35613
rect 9597 35560 9622 35575
rect 9678 35560 9703 35575
rect 9597 35557 9598 35560
rect 9759 35557 9983 35613
rect 10039 35557 10063 35613
rect 10119 35557 10143 35613
rect 10204 35575 10218 35627
rect 10270 35613 10706 35627
rect 10758 35613 10772 35627
rect 10824 35613 11260 35627
rect 11312 35613 11326 35627
rect 11378 35613 11814 35627
rect 11866 35613 11880 35627
rect 11932 35613 12368 35627
rect 10199 35560 10223 35575
rect 8054 35525 8490 35557
rect 8542 35525 8556 35557
rect 8608 35525 9044 35557
rect 9096 35525 9110 35557
rect 9162 35525 9598 35557
rect 9650 35525 9664 35557
rect 9716 35525 10152 35557
rect 7977 35493 8002 35508
rect 7500 35441 7936 35469
rect 7988 35441 8002 35493
rect 8058 35469 8083 35525
rect 8139 35469 8164 35525
rect 8220 35469 8245 35525
rect 8301 35469 8326 35525
rect 8382 35469 8407 35525
rect 8463 35469 8488 35525
rect 8544 35508 8556 35525
rect 8544 35493 8569 35508
rect 8544 35469 8556 35493
rect 8625 35469 8650 35525
rect 8706 35469 8731 35525
rect 8787 35469 8812 35525
rect 8868 35469 8893 35525
rect 8949 35469 8974 35525
rect 9030 35508 9044 35525
rect 9030 35493 9055 35508
rect 9111 35493 9136 35508
rect 9030 35469 9044 35493
rect 9192 35469 9217 35525
rect 9273 35469 9298 35525
rect 9354 35469 9379 35525
rect 9435 35469 9460 35525
rect 9516 35469 9541 35525
rect 9597 35508 9598 35525
rect 9597 35493 9622 35508
rect 9678 35493 9703 35508
rect 9597 35469 9598 35493
rect 9759 35469 9983 35525
rect 10039 35469 10063 35525
rect 10119 35469 10143 35525
rect 10204 35508 10218 35560
rect 10279 35557 10303 35613
rect 10359 35557 10383 35613
rect 10439 35557 10463 35613
rect 10519 35557 10544 35613
rect 10600 35557 10625 35613
rect 10681 35557 10706 35613
rect 10762 35575 10772 35613
rect 10762 35560 10787 35575
rect 10762 35557 10772 35560
rect 10843 35557 10868 35613
rect 10924 35557 10949 35613
rect 11005 35557 11030 35613
rect 11086 35557 11111 35613
rect 11167 35557 11192 35613
rect 11248 35575 11260 35613
rect 11248 35560 11273 35575
rect 11329 35560 11354 35575
rect 11248 35557 11260 35560
rect 11410 35557 11435 35613
rect 11491 35557 11516 35613
rect 11572 35557 11597 35613
rect 11653 35557 11678 35613
rect 11734 35557 11759 35613
rect 11815 35560 11840 35575
rect 11896 35560 11921 35575
rect 11977 35557 12002 35613
rect 12058 35575 12368 35613
rect 12420 35575 12434 35627
rect 12486 35575 12922 35627
rect 12974 35575 12988 35627
rect 13040 35575 13317 35627
rect 12058 35560 13317 35575
rect 12058 35557 12368 35560
rect 10270 35525 10706 35557
rect 10758 35525 10772 35557
rect 10824 35525 11260 35557
rect 11312 35525 11326 35557
rect 11378 35525 11814 35557
rect 11866 35525 11880 35557
rect 11932 35525 12368 35557
rect 10199 35493 10223 35508
rect 8054 35441 8490 35469
rect 8542 35441 8556 35469
rect 8608 35441 9044 35469
rect 9096 35441 9110 35469
rect 9162 35441 9598 35469
rect 9650 35441 9664 35469
rect 9716 35441 10152 35469
rect 10204 35441 10218 35493
rect 10279 35469 10303 35525
rect 10359 35469 10383 35525
rect 10439 35469 10463 35525
rect 10519 35469 10544 35525
rect 10600 35469 10625 35525
rect 10681 35469 10706 35525
rect 10762 35508 10772 35525
rect 10762 35493 10787 35508
rect 10762 35469 10772 35493
rect 10843 35469 10868 35525
rect 10924 35469 10949 35525
rect 11005 35469 11030 35525
rect 11086 35469 11111 35525
rect 11167 35469 11192 35525
rect 11248 35508 11260 35525
rect 11248 35493 11273 35508
rect 11329 35493 11354 35508
rect 11248 35469 11260 35493
rect 11410 35469 11435 35525
rect 11491 35469 11516 35525
rect 11572 35469 11597 35525
rect 11653 35469 11678 35525
rect 11734 35469 11759 35525
rect 11815 35493 11840 35508
rect 11896 35493 11921 35508
rect 11977 35469 12002 35525
rect 12058 35508 12368 35525
rect 12420 35508 12434 35560
rect 12486 35508 12922 35560
rect 12974 35508 12988 35560
rect 13040 35508 13317 35560
rect 12058 35493 13317 35508
rect 12058 35469 12368 35493
rect 10270 35441 10706 35469
rect 10758 35441 10772 35469
rect 10824 35441 11260 35469
rect 11312 35441 11326 35469
rect 11378 35441 11814 35469
rect 11866 35441 11880 35469
rect 11932 35441 12368 35469
rect 12420 35441 12434 35493
rect 12486 35441 12922 35493
rect 12974 35441 12988 35493
rect 13040 35441 13317 35493
rect 3504 35437 13317 35441
rect 3504 35426 5215 35437
rect 5271 35426 5296 35437
rect 3569 35374 3570 35426
rect 3504 35370 3513 35374
rect 3569 35370 3593 35374
rect 3649 35370 3673 35426
rect 3729 35370 3753 35426
rect 3809 35370 3833 35426
rect 3889 35370 3913 35426
rect 3969 35370 3993 35426
rect 4049 35374 4058 35426
rect 4049 35370 4073 35374
rect 4129 35370 4153 35374
rect 4209 35370 4233 35426
rect 4289 35370 4314 35426
rect 4370 35370 4395 35426
rect 4451 35370 4476 35426
rect 4532 35370 4557 35426
rect 4613 35370 4638 35374
rect 4694 35370 4719 35374
rect 4775 35370 4800 35426
rect 4856 35370 4881 35426
rect 4937 35370 4962 35426
rect 5018 35374 5166 35426
rect 5284 35381 5296 35426
rect 5352 35381 5377 35437
rect 5433 35381 5458 35437
rect 5514 35381 5539 35437
rect 5595 35381 5620 35437
rect 5676 35381 5701 35437
rect 5757 35426 5782 35437
rect 5772 35381 5782 35426
rect 5838 35381 5863 35437
rect 5919 35381 5944 35437
rect 6000 35381 6025 35437
rect 6081 35381 6106 35437
rect 6162 35381 6187 35437
rect 6243 35381 6268 35437
rect 6324 35426 6349 35437
rect 5218 35374 5232 35381
rect 5284 35374 5720 35381
rect 5772 35374 5786 35381
rect 5838 35374 6274 35381
rect 6326 35374 6340 35426
rect 6405 35381 6430 35437
rect 6486 35381 6511 35437
rect 6567 35381 6592 35437
rect 6648 35381 6673 35437
rect 6729 35381 6754 35437
rect 6810 35426 6835 35437
rect 6891 35426 6916 35437
rect 6810 35381 6828 35426
rect 6891 35381 6894 35426
rect 6972 35381 6997 35437
rect 7053 35381 7078 35437
rect 7134 35381 7159 35437
rect 7215 35381 7240 35437
rect 7296 35381 7320 35437
rect 7376 35426 7598 35437
rect 7376 35381 7382 35426
rect 6392 35374 6828 35381
rect 6880 35374 6894 35381
rect 6946 35374 7382 35381
rect 7434 35374 7448 35426
rect 7500 35381 7598 35426
rect 7654 35381 7678 35437
rect 7734 35381 7759 35437
rect 7815 35381 7840 35437
rect 7896 35381 7921 35437
rect 7977 35426 8002 35437
rect 7500 35374 7936 35381
rect 7988 35374 8002 35426
rect 8058 35381 8083 35437
rect 8139 35381 8164 35437
rect 8220 35381 8245 35437
rect 8301 35381 8326 35437
rect 8382 35381 8407 35437
rect 8463 35381 8488 35437
rect 8544 35426 8569 35437
rect 8544 35381 8556 35426
rect 8625 35381 8650 35437
rect 8706 35381 8731 35437
rect 8787 35381 8812 35437
rect 8868 35381 8893 35437
rect 8949 35381 8974 35437
rect 9030 35426 9055 35437
rect 9111 35426 9136 35437
rect 9030 35381 9044 35426
rect 9192 35381 9217 35437
rect 9273 35381 9298 35437
rect 9354 35381 9379 35437
rect 9435 35381 9460 35437
rect 9516 35381 9541 35437
rect 9597 35426 9622 35437
rect 9678 35426 9703 35437
rect 9597 35381 9598 35426
rect 9759 35381 9983 35437
rect 10039 35381 10063 35437
rect 10119 35381 10143 35437
rect 10199 35426 10223 35437
rect 8054 35374 8490 35381
rect 8542 35374 8556 35381
rect 8608 35374 9044 35381
rect 9096 35374 9110 35381
rect 9162 35374 9598 35381
rect 9650 35374 9664 35381
rect 9716 35374 10152 35381
rect 10204 35374 10218 35426
rect 10279 35381 10303 35437
rect 10359 35381 10383 35437
rect 10439 35381 10463 35437
rect 10519 35381 10544 35437
rect 10600 35381 10625 35437
rect 10681 35381 10706 35437
rect 10762 35426 10787 35437
rect 10762 35381 10772 35426
rect 10843 35381 10868 35437
rect 10924 35381 10949 35437
rect 11005 35381 11030 35437
rect 11086 35381 11111 35437
rect 11167 35381 11192 35437
rect 11248 35426 11273 35437
rect 11329 35426 11354 35437
rect 11248 35381 11260 35426
rect 11410 35381 11435 35437
rect 11491 35381 11516 35437
rect 11572 35381 11597 35437
rect 11653 35381 11678 35437
rect 11734 35381 11759 35437
rect 11815 35426 11840 35437
rect 11896 35426 11921 35437
rect 11977 35381 12002 35437
rect 12058 35426 13317 35437
rect 12058 35381 12368 35426
rect 10270 35374 10706 35381
rect 10758 35374 10772 35381
rect 10824 35374 11260 35381
rect 11312 35374 11326 35381
rect 11378 35374 11814 35381
rect 11866 35374 11880 35381
rect 11932 35374 12368 35381
rect 12420 35374 12434 35426
rect 12486 35374 12922 35426
rect 12974 35374 12988 35426
rect 13040 35374 13317 35426
rect 5018 35370 13317 35374
rect 3504 35368 13317 35370
rect 100 35328 2792 35340
rect 100 35276 2249 35328
rect 2301 35276 2315 35328
rect 2367 35276 2792 35328
rect 100 35264 2792 35276
rect 100 35212 2249 35264
rect 2301 35212 2315 35264
rect 2367 35212 2792 35264
rect 100 35200 2792 35212
rect 100 35148 2249 35200
rect 2301 35148 2315 35200
rect 2367 35148 2792 35200
rect 100 35136 2792 35148
rect 100 35084 2249 35136
rect 2301 35084 2315 35136
rect 2367 35084 2792 35136
rect 100 35072 2792 35084
rect 100 35020 2249 35072
rect 2301 35020 2315 35072
rect 2367 35020 2792 35072
rect 100 35008 2792 35020
rect 100 34956 2249 35008
rect 2301 34956 2315 35008
rect 2367 34956 2792 35008
rect 100 34944 2792 34956
rect 100 34892 2249 34944
rect 2301 34892 2315 34944
rect 2367 34892 2792 34944
rect 100 34880 2792 34892
rect 100 34828 2249 34880
rect 2301 34828 2315 34880
rect 2367 34828 2792 34880
rect 100 34816 2792 34828
rect 100 34764 2249 34816
rect 2301 34764 2315 34816
rect 2367 34764 2792 34816
rect 100 34752 2792 34764
rect 100 34700 2249 34752
rect 2301 34700 2315 34752
rect 2367 34726 2792 34752
tri 2792 34726 3002 34936 sw
rect 2367 34720 13602 34726
rect 2367 34700 3167 34720
rect 100 34688 3167 34700
rect 100 34636 2249 34688
rect 2301 34636 2315 34688
rect 2367 34668 3167 34688
rect 3219 34668 3233 34720
rect 3285 34668 4003 34720
rect 4055 34668 4069 34720
rect 4121 34668 4839 34720
rect 4891 34668 4905 34720
rect 4957 34668 5675 34720
rect 5727 34668 5741 34720
rect 5793 34668 6511 34720
rect 6563 34668 6577 34720
rect 6629 34668 7347 34720
rect 7399 34668 7413 34720
rect 7465 34668 8183 34720
rect 8235 34668 8249 34720
rect 8301 34668 9019 34720
rect 9071 34668 9085 34720
rect 9137 34668 9855 34720
rect 9907 34668 9921 34720
rect 9973 34668 10691 34720
rect 10743 34668 10757 34720
rect 10809 34668 11527 34720
rect 11579 34668 11593 34720
rect 11645 34668 12363 34720
rect 12415 34668 12429 34720
rect 12481 34668 13200 34720
rect 13252 34668 13270 34720
rect 13322 34668 13340 34720
rect 13392 34668 13410 34720
rect 13462 34668 13480 34720
rect 13532 34668 13550 34720
rect 2367 34654 13602 34668
rect 2367 34636 3167 34654
rect 100 34624 3167 34636
rect 100 34572 2249 34624
rect 2301 34572 2315 34624
rect 2367 34602 3167 34624
rect 3219 34602 3233 34654
rect 3285 34602 4003 34654
rect 4055 34602 4069 34654
rect 4121 34602 4839 34654
rect 4891 34602 4905 34654
rect 4957 34602 5675 34654
rect 5727 34602 5741 34654
rect 5793 34602 6511 34654
rect 6563 34602 6577 34654
rect 6629 34602 7347 34654
rect 7399 34602 7413 34654
rect 7465 34602 8183 34654
rect 8235 34602 8249 34654
rect 8301 34602 9019 34654
rect 9071 34602 9085 34654
rect 9137 34602 9855 34654
rect 9907 34602 9921 34654
rect 9973 34602 10691 34654
rect 10743 34602 10757 34654
rect 10809 34602 11527 34654
rect 11579 34602 11593 34654
rect 11645 34602 12363 34654
rect 12415 34602 12429 34654
rect 12481 34602 13200 34654
rect 13252 34602 13270 34654
rect 13322 34602 13340 34654
rect 13392 34602 13410 34654
rect 13462 34602 13480 34654
rect 13532 34602 13550 34654
rect 2367 34588 13602 34602
rect 2367 34572 3167 34588
rect 100 34560 3167 34572
rect 100 34508 2249 34560
rect 2301 34508 2315 34560
rect 2367 34536 3167 34560
rect 3219 34536 3233 34588
rect 3285 34536 4003 34588
rect 4055 34536 4069 34588
rect 4121 34536 4839 34588
rect 4891 34536 4905 34588
rect 4957 34536 5675 34588
rect 5727 34536 5741 34588
rect 5793 34536 6511 34588
rect 6563 34536 6577 34588
rect 6629 34536 7347 34588
rect 7399 34536 7413 34588
rect 7465 34536 8183 34588
rect 8235 34536 8249 34588
rect 8301 34536 9019 34588
rect 9071 34536 9085 34588
rect 9137 34536 9855 34588
rect 9907 34536 9921 34588
rect 9973 34536 10691 34588
rect 10743 34536 10757 34588
rect 10809 34536 11527 34588
rect 11579 34536 11593 34588
rect 11645 34536 12363 34588
rect 12415 34536 12429 34588
rect 12481 34536 13200 34588
rect 13252 34536 13270 34588
rect 13322 34536 13340 34588
rect 13392 34536 13410 34588
rect 13462 34536 13480 34588
rect 13532 34536 13550 34588
rect 2367 34522 13602 34536
rect 2367 34508 3167 34522
rect 100 34496 3167 34508
rect 100 34444 2249 34496
rect 2301 34444 2315 34496
rect 2367 34470 3167 34496
rect 3219 34470 3233 34522
rect 3285 34470 4003 34522
rect 4055 34470 4069 34522
rect 4121 34470 4839 34522
rect 4891 34470 4905 34522
rect 4957 34470 5675 34522
rect 5727 34470 5741 34522
rect 5793 34470 6511 34522
rect 6563 34470 6577 34522
rect 6629 34470 7347 34522
rect 7399 34470 7413 34522
rect 7465 34470 8183 34522
rect 8235 34470 8249 34522
rect 8301 34470 9019 34522
rect 9071 34470 9085 34522
rect 9137 34470 9855 34522
rect 9907 34470 9921 34522
rect 9973 34470 10691 34522
rect 10743 34470 10757 34522
rect 10809 34470 11527 34522
rect 11579 34470 11593 34522
rect 11645 34470 12363 34522
rect 12415 34470 12429 34522
rect 12481 34470 13200 34522
rect 13252 34470 13270 34522
rect 13322 34470 13340 34522
rect 13392 34470 13410 34522
rect 13462 34470 13480 34522
rect 13532 34470 13550 34522
rect 2367 34456 13602 34470
rect 2367 34444 3167 34456
rect 100 34432 3167 34444
rect 100 34380 2249 34432
rect 2301 34380 2315 34432
rect 2367 34404 3167 34432
rect 3219 34404 3233 34456
rect 3285 34404 4003 34456
rect 4055 34404 4069 34456
rect 4121 34404 4839 34456
rect 4891 34404 4905 34456
rect 4957 34404 5675 34456
rect 5727 34404 5741 34456
rect 5793 34404 6511 34456
rect 6563 34404 6577 34456
rect 6629 34404 7347 34456
rect 7399 34404 7413 34456
rect 7465 34404 8183 34456
rect 8235 34404 8249 34456
rect 8301 34404 9019 34456
rect 9071 34404 9085 34456
rect 9137 34404 9855 34456
rect 9907 34404 9921 34456
rect 9973 34404 10691 34456
rect 10743 34404 10757 34456
rect 10809 34404 11527 34456
rect 11579 34404 11593 34456
rect 11645 34404 12363 34456
rect 12415 34404 12429 34456
rect 12481 34404 13200 34456
rect 13252 34404 13270 34456
rect 13322 34404 13340 34456
rect 13392 34404 13410 34456
rect 13462 34404 13480 34456
rect 13532 34404 13550 34456
rect 2367 34390 13602 34404
rect 2367 34380 3167 34390
rect 100 34368 3167 34380
rect 100 34316 2249 34368
rect 2301 34316 2315 34368
rect 2367 34338 3167 34368
rect 3219 34338 3233 34390
rect 3285 34338 4003 34390
rect 4055 34338 4069 34390
rect 4121 34338 4839 34390
rect 4891 34338 4905 34390
rect 4957 34338 5675 34390
rect 5727 34338 5741 34390
rect 5793 34338 6511 34390
rect 6563 34338 6577 34390
rect 6629 34338 7347 34390
rect 7399 34338 7413 34390
rect 7465 34338 8183 34390
rect 8235 34338 8249 34390
rect 8301 34338 9019 34390
rect 9071 34338 9085 34390
rect 9137 34338 9855 34390
rect 9907 34338 9921 34390
rect 9973 34338 10691 34390
rect 10743 34338 10757 34390
rect 10809 34338 11527 34390
rect 11579 34338 11593 34390
rect 11645 34338 12363 34390
rect 12415 34338 12429 34390
rect 12481 34338 13200 34390
rect 13252 34338 13270 34390
rect 13322 34338 13340 34390
rect 13392 34338 13410 34390
rect 13462 34338 13480 34390
rect 13532 34338 13550 34390
rect 2367 34323 13602 34338
rect 2367 34316 3167 34323
rect 100 34304 3167 34316
rect 100 34252 2249 34304
rect 2301 34252 2315 34304
rect 2367 34271 3167 34304
rect 3219 34271 3233 34323
rect 3285 34271 4003 34323
rect 4055 34271 4069 34323
rect 4121 34271 4839 34323
rect 4891 34271 4905 34323
rect 4957 34271 5675 34323
rect 5727 34271 5741 34323
rect 5793 34271 6511 34323
rect 6563 34271 6577 34323
rect 6629 34271 7347 34323
rect 7399 34271 7413 34323
rect 7465 34271 8183 34323
rect 8235 34271 8249 34323
rect 8301 34271 9019 34323
rect 9071 34271 9085 34323
rect 9137 34271 9855 34323
rect 9907 34271 9921 34323
rect 9973 34271 10691 34323
rect 10743 34271 10757 34323
rect 10809 34271 11527 34323
rect 11579 34271 11593 34323
rect 11645 34271 12363 34323
rect 12415 34271 12429 34323
rect 12481 34271 13200 34323
rect 13252 34271 13270 34323
rect 13322 34271 13340 34323
rect 13392 34271 13410 34323
rect 13462 34271 13480 34323
rect 13532 34271 13550 34323
rect 2367 34256 13602 34271
rect 2367 34252 3167 34256
rect 100 34240 3167 34252
rect 100 34188 2249 34240
rect 2301 34188 2315 34240
rect 2367 34204 3167 34240
rect 3219 34204 3233 34256
rect 3285 34204 4003 34256
rect 4055 34204 4069 34256
rect 4121 34204 4839 34256
rect 4891 34204 4905 34256
rect 4957 34204 5675 34256
rect 5727 34204 5741 34256
rect 5793 34204 6511 34256
rect 6563 34204 6577 34256
rect 6629 34204 7347 34256
rect 7399 34204 7413 34256
rect 7465 34204 8183 34256
rect 8235 34204 8249 34256
rect 8301 34204 9019 34256
rect 9071 34204 9085 34256
rect 9137 34204 9855 34256
rect 9907 34204 9921 34256
rect 9973 34204 10691 34256
rect 10743 34204 10757 34256
rect 10809 34204 11527 34256
rect 11579 34204 11593 34256
rect 11645 34204 12363 34256
rect 12415 34204 12429 34256
rect 12481 34204 13200 34256
rect 13252 34204 13270 34256
rect 13322 34204 13340 34256
rect 13392 34204 13410 34256
rect 13462 34204 13480 34256
rect 13532 34204 13550 34256
rect 2367 34198 13602 34204
rect 2367 34188 2792 34198
rect 100 34176 2792 34188
rect 100 34124 2249 34176
rect 2301 34124 2315 34176
rect 2367 34124 2792 34176
rect 100 34112 2792 34124
rect 100 34060 2249 34112
rect 2301 34060 2315 34112
rect 2367 34060 2792 34112
rect 100 34048 2792 34060
rect 100 33996 2249 34048
rect 2301 33996 2315 34048
rect 2367 33996 2792 34048
rect 100 33984 2792 33996
tri 2792 33988 3002 34198 nw
rect 100 33932 2249 33984
rect 2301 33932 2315 33984
rect 2367 33932 2792 33984
rect 100 33920 2792 33932
rect 100 33868 2249 33920
rect 2301 33868 2315 33920
rect 2367 33868 2792 33920
rect 100 33856 2792 33868
rect 100 33804 2249 33856
rect 2301 33804 2315 33856
rect 2367 33804 2792 33856
rect 100 33792 2792 33804
rect 100 33740 2249 33792
rect 2301 33740 2315 33792
rect 2367 33740 2792 33792
rect 100 33728 2792 33740
rect 100 33676 2249 33728
rect 2301 33676 2315 33728
rect 2367 33676 2792 33728
rect 100 33664 2792 33676
rect 100 33612 2249 33664
rect 2301 33612 2315 33664
rect 2367 33612 2792 33664
rect 100 33600 2792 33612
rect 100 33548 2249 33600
rect 2301 33548 2315 33600
rect 2367 33548 2792 33600
rect 100 33536 2792 33548
rect 100 33484 2249 33536
rect 2301 33484 2315 33536
rect 2367 33484 2792 33536
rect 100 33472 2792 33484
rect 100 33420 2249 33472
rect 2301 33420 2315 33472
rect 2367 33420 2792 33472
rect 100 33408 2792 33420
rect 100 33356 2249 33408
rect 2301 33356 2315 33408
rect 2367 33356 2792 33408
rect 3504 33896 13317 33898
rect 3504 33840 3513 33896
rect 3569 33892 3594 33896
rect 3650 33892 3675 33896
rect 3569 33840 3585 33892
rect 3650 33840 3651 33892
rect 3731 33840 3757 33896
rect 3813 33840 3839 33896
rect 3895 33840 3921 33896
rect 3977 33840 4003 33896
rect 4059 33840 4085 33896
rect 4141 33840 4167 33896
rect 4223 33840 4249 33896
rect 4305 33892 13317 33896
rect 4305 33880 4421 33892
rect 4473 33880 4487 33892
rect 4539 33886 5257 33892
rect 4305 33840 4354 33880
rect 3504 33826 4354 33840
rect 3504 33802 3585 33826
rect 3637 33802 3651 33826
rect 3703 33824 4354 33826
rect 4410 33840 4421 33880
rect 4539 33840 4556 33886
rect 4410 33826 4446 33840
rect 4502 33830 4556 33840
rect 4612 33878 5257 33886
rect 5309 33878 5323 33892
rect 5375 33878 6093 33892
rect 6145 33878 6159 33892
rect 6211 33878 6929 33892
rect 6981 33878 6995 33892
rect 7047 33878 7765 33892
rect 4612 33830 5216 33878
rect 5375 33840 5382 33878
rect 4502 33826 5216 33830
rect 5272 33826 5299 33840
rect 5355 33826 5382 33840
rect 4410 33824 4421 33826
rect 3703 33802 4421 33824
rect 3504 33746 3513 33802
rect 3569 33774 3585 33802
rect 3650 33774 3651 33802
rect 3569 33760 3594 33774
rect 3650 33760 3675 33774
rect 3569 33746 3585 33760
rect 3650 33746 3651 33760
rect 3731 33746 3757 33802
rect 3813 33746 3839 33802
rect 3895 33746 3921 33802
rect 3977 33746 4003 33802
rect 4059 33746 4085 33802
rect 4141 33746 4167 33802
rect 4223 33746 4249 33802
rect 4305 33780 4421 33802
rect 4473 33780 4487 33824
rect 4539 33822 5216 33826
rect 5375 33822 5382 33826
rect 5438 33822 5465 33878
rect 5521 33822 5548 33878
rect 5604 33822 5631 33878
rect 5687 33822 5714 33878
rect 5770 33822 5797 33878
rect 5853 33822 5880 33878
rect 5936 33822 5963 33878
rect 6019 33822 6046 33878
rect 6102 33826 6129 33840
rect 6185 33826 6211 33840
rect 6267 33822 6293 33878
rect 6349 33822 6375 33878
rect 6431 33822 6457 33878
rect 6513 33822 6539 33878
rect 6595 33822 6621 33878
rect 6677 33822 6703 33878
rect 6759 33822 6785 33878
rect 6841 33822 6867 33878
rect 6923 33840 6929 33878
rect 6923 33826 6949 33840
rect 7005 33826 7031 33840
rect 6923 33822 6929 33826
rect 7087 33822 7113 33878
rect 7169 33822 7195 33878
rect 7251 33858 7765 33878
rect 7251 33822 7636 33858
rect 4539 33804 5257 33822
rect 4305 33746 4354 33780
rect 3504 33708 3585 33746
rect 3637 33708 3651 33746
rect 3703 33724 4354 33746
rect 4410 33774 4421 33780
rect 4539 33774 4556 33804
rect 4410 33760 4446 33774
rect 4502 33760 4556 33774
rect 4410 33724 4421 33760
rect 4539 33748 4556 33760
rect 4612 33790 5257 33804
rect 5309 33790 5323 33822
rect 5375 33790 6093 33822
rect 6145 33790 6159 33822
rect 6211 33790 6929 33822
rect 6981 33790 6995 33822
rect 7047 33802 7636 33822
rect 7692 33802 7716 33858
rect 7817 33840 7831 33892
rect 7883 33881 8601 33892
rect 7772 33826 7838 33840
rect 7047 33790 7765 33802
rect 4612 33748 5216 33790
rect 5375 33774 5382 33790
rect 5272 33760 5299 33774
rect 5355 33760 5382 33774
rect 4539 33734 5216 33748
rect 5375 33734 5382 33760
rect 5438 33734 5465 33790
rect 5521 33734 5548 33790
rect 5604 33734 5631 33790
rect 5687 33734 5714 33790
rect 5770 33734 5797 33790
rect 5853 33734 5880 33790
rect 5936 33734 5963 33790
rect 6019 33734 6046 33790
rect 6102 33760 6129 33774
rect 6185 33760 6211 33774
rect 6267 33734 6293 33790
rect 6349 33734 6375 33790
rect 6431 33734 6457 33790
rect 6513 33734 6539 33790
rect 6595 33734 6621 33790
rect 6677 33734 6703 33790
rect 6759 33734 6785 33790
rect 6841 33734 6867 33790
rect 6923 33774 6929 33790
rect 6923 33760 6949 33774
rect 7005 33760 7031 33774
rect 6923 33734 6929 33760
rect 7087 33734 7113 33790
rect 7169 33734 7195 33790
rect 7251 33774 7765 33790
rect 7817 33774 7831 33826
rect 7894 33825 7922 33881
rect 7978 33878 8601 33881
rect 8653 33878 8667 33892
rect 8719 33878 9437 33892
rect 9489 33878 9503 33892
rect 9555 33881 10273 33892
rect 10325 33881 10339 33892
rect 9555 33878 10202 33881
rect 7978 33825 8041 33878
rect 7883 33822 8041 33825
rect 8097 33822 8124 33878
rect 8180 33822 8207 33878
rect 8263 33822 8290 33878
rect 8346 33822 8373 33878
rect 8429 33822 8456 33878
rect 8512 33822 8539 33878
rect 8595 33840 8601 33878
rect 8595 33826 8622 33840
rect 8678 33826 8705 33840
rect 8595 33822 8601 33826
rect 8761 33822 8788 33878
rect 8844 33822 8871 33878
rect 8927 33822 8954 33878
rect 9010 33822 9037 33878
rect 9093 33822 9120 33878
rect 9176 33822 9203 33878
rect 9259 33822 9286 33878
rect 9342 33822 9369 33878
rect 9425 33840 9437 33878
rect 9425 33826 9452 33840
rect 9508 33826 9535 33840
rect 9425 33822 9437 33826
rect 9591 33822 9618 33878
rect 9674 33822 9702 33878
rect 9758 33858 10202 33878
rect 9758 33822 10000 33858
rect 7883 33790 8601 33822
rect 8653 33790 8667 33822
rect 8719 33790 9437 33822
rect 9489 33790 9503 33822
rect 9555 33802 10000 33822
rect 10056 33802 10080 33858
rect 10136 33825 10202 33858
rect 10258 33840 10273 33881
rect 10391 33878 11109 33892
rect 11161 33878 11175 33892
rect 11227 33878 11945 33892
rect 11997 33878 12011 33892
rect 10391 33840 10397 33878
rect 10258 33826 10286 33840
rect 10342 33826 10397 33840
rect 10258 33825 10273 33826
rect 10136 33802 10273 33825
rect 9555 33790 10273 33802
rect 7883 33774 8041 33790
rect 7251 33766 8041 33774
rect 7251 33760 7838 33766
rect 7251 33751 7765 33760
rect 7251 33734 7723 33751
rect 3703 33708 4421 33724
rect 4473 33708 4487 33724
rect 4539 33708 5257 33734
rect 5309 33708 5323 33734
rect 5375 33708 6093 33734
rect 6145 33708 6159 33734
rect 6211 33708 6929 33734
rect 6981 33708 6995 33734
rect 7047 33708 7723 33734
rect 7817 33708 7831 33760
rect 7894 33710 7922 33766
rect 7978 33734 8041 33766
rect 8097 33734 8124 33790
rect 8180 33734 8207 33790
rect 8263 33734 8290 33790
rect 8346 33734 8373 33790
rect 8429 33734 8456 33790
rect 8512 33734 8539 33790
rect 8595 33774 8601 33790
rect 8595 33760 8622 33774
rect 8678 33760 8705 33774
rect 8595 33734 8601 33760
rect 8761 33734 8788 33790
rect 8844 33734 8871 33790
rect 8927 33734 8954 33790
rect 9010 33734 9037 33790
rect 9093 33734 9120 33790
rect 9176 33734 9203 33790
rect 9259 33734 9286 33790
rect 9342 33734 9369 33790
rect 9425 33774 9437 33790
rect 9425 33760 9452 33774
rect 9508 33760 9535 33774
rect 9425 33734 9437 33760
rect 9591 33734 9618 33790
rect 9674 33734 9702 33790
rect 9758 33774 10273 33790
rect 10325 33774 10339 33825
rect 10391 33822 10397 33826
rect 10453 33822 10477 33878
rect 10533 33822 10557 33878
rect 10613 33822 10637 33878
rect 10693 33822 10717 33878
rect 10773 33822 10797 33878
rect 10853 33822 10877 33878
rect 10933 33822 10957 33878
rect 11013 33822 11037 33878
rect 11093 33840 11109 33878
rect 11173 33840 11175 33878
rect 11093 33826 11117 33840
rect 11173 33826 11197 33840
rect 11093 33822 11109 33826
rect 11173 33822 11175 33826
rect 11253 33822 11277 33878
rect 11333 33822 11357 33878
rect 11413 33822 11437 33878
rect 11493 33822 11517 33878
rect 11573 33822 11597 33878
rect 11653 33822 11677 33878
rect 11733 33822 11758 33878
rect 11814 33822 11839 33878
rect 11895 33822 11920 33878
rect 11997 33840 12001 33878
rect 12063 33840 12781 33892
rect 12833 33840 12847 33892
rect 12899 33840 13317 33892
rect 11976 33826 12001 33840
rect 12057 33826 13317 33840
rect 11997 33822 12001 33826
rect 10391 33790 11109 33822
rect 11161 33790 11175 33822
rect 11227 33790 11945 33822
rect 11997 33790 12011 33822
rect 10391 33774 10397 33790
rect 9758 33766 10397 33774
rect 9758 33751 10202 33766
rect 9758 33734 10087 33751
rect 7978 33710 8601 33734
rect 7883 33708 8601 33710
rect 8653 33708 8667 33734
rect 8719 33708 9437 33734
rect 9489 33708 9503 33734
rect 9555 33708 10087 33734
rect 3504 33652 3513 33708
rect 3569 33694 3594 33708
rect 3650 33694 3675 33708
rect 3569 33652 3585 33694
rect 3650 33652 3651 33694
rect 3731 33652 3757 33708
rect 3813 33652 3839 33708
rect 3895 33652 3921 33708
rect 3977 33652 4003 33708
rect 4059 33652 4085 33708
rect 4141 33652 4167 33708
rect 4223 33652 4249 33708
rect 4305 33702 7723 33708
rect 4305 33694 5216 33702
rect 5272 33694 5299 33702
rect 5355 33694 5382 33702
rect 4305 33679 4421 33694
rect 4473 33679 4487 33694
rect 4305 33652 4354 33679
rect 3504 33642 3585 33652
rect 3637 33642 3651 33652
rect 3703 33642 4354 33652
rect 3504 33627 4354 33642
rect 3504 33614 3585 33627
rect 3637 33614 3651 33627
rect 3703 33623 4354 33627
rect 4410 33642 4421 33679
rect 4539 33646 5216 33694
rect 5375 33646 5382 33694
rect 5438 33646 5465 33702
rect 5521 33646 5548 33702
rect 5604 33646 5631 33702
rect 5687 33646 5714 33702
rect 5770 33646 5797 33702
rect 5853 33646 5880 33702
rect 5936 33646 5963 33702
rect 6019 33646 6046 33702
rect 6102 33694 6129 33702
rect 6185 33694 6211 33702
rect 6267 33646 6293 33702
rect 6349 33646 6375 33702
rect 6431 33646 6457 33702
rect 6513 33646 6539 33702
rect 6595 33646 6621 33702
rect 6677 33646 6703 33702
rect 6759 33646 6785 33702
rect 6841 33646 6867 33702
rect 6923 33694 6949 33702
rect 7005 33694 7031 33702
rect 6923 33646 6929 33694
rect 7087 33646 7113 33702
rect 7169 33646 7195 33702
rect 7251 33695 7723 33702
rect 7779 33702 10087 33708
rect 7779 33695 8041 33702
rect 7251 33694 8041 33695
rect 7251 33646 7765 33694
rect 4539 33642 5257 33646
rect 5309 33642 5323 33646
rect 5375 33642 6093 33646
rect 6145 33642 6159 33646
rect 6211 33642 6929 33646
rect 6981 33642 6995 33646
rect 7047 33642 7765 33646
rect 7817 33642 7831 33694
rect 7883 33650 8041 33694
rect 4410 33627 4446 33642
rect 4502 33627 7838 33642
rect 4410 33623 4421 33627
rect 3703 33614 4421 33623
rect 3504 33558 3513 33614
rect 3569 33575 3585 33614
rect 3650 33575 3651 33614
rect 3569 33560 3594 33575
rect 3650 33560 3675 33575
rect 3569 33558 3585 33560
rect 3650 33558 3651 33560
rect 3731 33558 3757 33614
rect 3813 33558 3839 33614
rect 3895 33558 3921 33614
rect 3977 33558 4003 33614
rect 4059 33558 4085 33614
rect 4141 33558 4167 33614
rect 4223 33558 4249 33614
rect 4305 33575 4421 33614
rect 4473 33575 4487 33623
rect 4539 33614 5257 33627
rect 5309 33614 5323 33627
rect 5375 33614 6093 33627
rect 6145 33614 6159 33627
rect 6211 33614 6929 33627
rect 6981 33614 6995 33627
rect 7047 33614 7765 33627
rect 4539 33575 5216 33614
rect 5375 33575 5382 33614
rect 4305 33560 5216 33575
rect 5272 33560 5299 33575
rect 5355 33560 5382 33575
rect 4305 33558 4421 33560
rect 3504 33520 3585 33558
rect 3637 33520 3651 33558
rect 3703 33520 4421 33558
rect 3504 33464 3513 33520
rect 3569 33508 3585 33520
rect 3650 33508 3651 33520
rect 3569 33493 3594 33508
rect 3650 33493 3675 33508
rect 3569 33464 3585 33493
rect 3650 33464 3651 33493
rect 3731 33464 3757 33520
rect 3813 33464 3839 33520
rect 3895 33464 3921 33520
rect 3977 33464 4003 33520
rect 4059 33464 4085 33520
rect 4141 33464 4167 33520
rect 4223 33464 4249 33520
rect 4305 33508 4421 33520
rect 4473 33508 4487 33560
rect 4539 33558 5216 33560
rect 5375 33558 5382 33560
rect 5438 33558 5465 33614
rect 5521 33558 5548 33614
rect 5604 33558 5631 33614
rect 5687 33558 5714 33614
rect 5770 33558 5797 33614
rect 5853 33558 5880 33614
rect 5936 33558 5963 33614
rect 6019 33558 6046 33614
rect 6102 33560 6129 33575
rect 6185 33560 6211 33575
rect 6267 33558 6293 33614
rect 6349 33558 6375 33614
rect 6431 33558 6457 33614
rect 6513 33558 6539 33614
rect 6595 33558 6621 33614
rect 6677 33558 6703 33614
rect 6759 33558 6785 33614
rect 6841 33558 6867 33614
rect 6923 33575 6929 33614
rect 6923 33560 6949 33575
rect 7005 33560 7031 33575
rect 6923 33558 6929 33560
rect 7087 33558 7113 33614
rect 7169 33558 7195 33614
rect 7251 33575 7765 33614
rect 7817 33575 7831 33627
rect 7894 33594 7922 33650
rect 7978 33646 8041 33650
rect 8097 33646 8124 33702
rect 8180 33646 8207 33702
rect 8263 33646 8290 33702
rect 8346 33646 8373 33702
rect 8429 33646 8456 33702
rect 8512 33646 8539 33702
rect 8595 33694 8622 33702
rect 8678 33694 8705 33702
rect 8595 33646 8601 33694
rect 8761 33646 8788 33702
rect 8844 33646 8871 33702
rect 8927 33646 8954 33702
rect 9010 33646 9037 33702
rect 9093 33646 9120 33702
rect 9176 33646 9203 33702
rect 9259 33646 9286 33702
rect 9342 33646 9369 33702
rect 9425 33694 9452 33702
rect 9508 33694 9535 33702
rect 9425 33646 9437 33694
rect 9591 33646 9618 33702
rect 9674 33646 9702 33702
rect 9758 33695 10087 33702
rect 10143 33710 10202 33751
rect 10258 33760 10286 33766
rect 10342 33760 10397 33766
rect 10258 33710 10273 33760
rect 10391 33734 10397 33760
rect 10453 33734 10477 33790
rect 10533 33734 10557 33790
rect 10613 33734 10637 33790
rect 10693 33734 10717 33790
rect 10773 33734 10797 33790
rect 10853 33734 10877 33790
rect 10933 33734 10957 33790
rect 11013 33734 11037 33790
rect 11093 33774 11109 33790
rect 11173 33774 11175 33790
rect 11093 33760 11117 33774
rect 11173 33760 11197 33774
rect 11093 33734 11109 33760
rect 11173 33734 11175 33760
rect 11253 33734 11277 33790
rect 11333 33734 11357 33790
rect 11413 33734 11437 33790
rect 11493 33734 11517 33790
rect 11573 33734 11597 33790
rect 11653 33734 11677 33790
rect 11733 33734 11758 33790
rect 11814 33734 11839 33790
rect 11895 33734 11920 33790
rect 11997 33774 12001 33790
rect 12063 33774 12781 33826
rect 12833 33774 12847 33826
rect 12899 33774 13317 33826
rect 11976 33760 12001 33774
rect 12057 33760 13317 33774
rect 11997 33734 12001 33760
rect 10143 33708 10273 33710
rect 10325 33708 10339 33710
rect 10391 33708 11109 33734
rect 11161 33708 11175 33734
rect 11227 33708 11945 33734
rect 11997 33708 12011 33734
rect 12063 33708 12781 33760
rect 12833 33708 12847 33760
rect 12899 33708 13317 33760
rect 10143 33702 13317 33708
rect 10143 33695 10397 33702
rect 9758 33694 10397 33695
rect 9758 33650 10273 33694
rect 10325 33650 10339 33694
rect 9758 33646 10202 33650
rect 7978 33642 8601 33646
rect 8653 33642 8667 33646
rect 8719 33642 9437 33646
rect 9489 33642 9503 33646
rect 9555 33642 10202 33646
rect 7978 33627 10202 33642
rect 7978 33614 8601 33627
rect 8653 33614 8667 33627
rect 8719 33614 9437 33627
rect 9489 33614 9503 33627
rect 9555 33614 10202 33627
rect 7978 33594 8041 33614
rect 7883 33575 8041 33594
rect 7251 33560 8041 33575
rect 7251 33558 7765 33560
rect 4539 33526 5257 33558
rect 5309 33526 5323 33558
rect 5375 33526 6093 33558
rect 6145 33526 6159 33558
rect 6211 33526 6929 33558
rect 6981 33526 6995 33558
rect 7047 33526 7765 33558
rect 4539 33508 5216 33526
rect 5375 33508 5382 33526
rect 4305 33493 5216 33508
rect 5272 33493 5299 33508
rect 5355 33493 5382 33508
rect 4305 33464 4421 33493
rect 3504 33441 3585 33464
rect 3637 33441 3651 33464
rect 3703 33441 4421 33464
rect 4473 33441 4487 33493
rect 4539 33470 5216 33493
rect 5375 33470 5382 33493
rect 5438 33470 5465 33526
rect 5521 33470 5548 33526
rect 5604 33470 5631 33526
rect 5687 33470 5714 33526
rect 5770 33470 5797 33526
rect 5853 33470 5880 33526
rect 5936 33470 5963 33526
rect 6019 33470 6046 33526
rect 6102 33493 6129 33508
rect 6185 33493 6211 33508
rect 6267 33470 6293 33526
rect 6349 33470 6375 33526
rect 6431 33470 6457 33526
rect 6513 33470 6539 33526
rect 6595 33470 6621 33526
rect 6677 33470 6703 33526
rect 6759 33470 6785 33526
rect 6841 33470 6867 33526
rect 6923 33508 6929 33526
rect 6923 33493 6949 33508
rect 7005 33493 7031 33508
rect 6923 33470 6929 33493
rect 7087 33470 7113 33526
rect 7169 33470 7195 33526
rect 7251 33508 7765 33526
rect 7817 33508 7831 33560
rect 7883 33558 8041 33560
rect 8097 33558 8124 33614
rect 8180 33558 8207 33614
rect 8263 33558 8290 33614
rect 8346 33558 8373 33614
rect 8429 33558 8456 33614
rect 8512 33558 8539 33614
rect 8595 33575 8601 33614
rect 8595 33560 8622 33575
rect 8678 33560 8705 33575
rect 8595 33558 8601 33560
rect 8761 33558 8788 33614
rect 8844 33558 8871 33614
rect 8927 33558 8954 33614
rect 9010 33558 9037 33614
rect 9093 33558 9120 33614
rect 9176 33558 9203 33614
rect 9259 33558 9286 33614
rect 9342 33558 9369 33614
rect 9425 33575 9437 33614
rect 9425 33560 9452 33575
rect 9508 33560 9535 33575
rect 9425 33558 9437 33560
rect 9591 33558 9618 33614
rect 9674 33558 9702 33614
rect 9758 33594 10202 33614
rect 10258 33642 10273 33650
rect 10391 33646 10397 33694
rect 10453 33646 10477 33702
rect 10533 33646 10557 33702
rect 10613 33646 10637 33702
rect 10693 33646 10717 33702
rect 10773 33646 10797 33702
rect 10853 33646 10877 33702
rect 10933 33646 10957 33702
rect 11013 33646 11037 33702
rect 11093 33694 11117 33702
rect 11173 33694 11197 33702
rect 11093 33646 11109 33694
rect 11173 33646 11175 33694
rect 11253 33646 11277 33702
rect 11333 33646 11357 33702
rect 11413 33646 11437 33702
rect 11493 33646 11517 33702
rect 11573 33646 11597 33702
rect 11653 33646 11677 33702
rect 11733 33646 11758 33702
rect 11814 33646 11839 33702
rect 11895 33646 11920 33702
rect 11976 33694 12001 33702
rect 12057 33694 13317 33702
rect 11997 33646 12001 33694
rect 10391 33642 11109 33646
rect 11161 33642 11175 33646
rect 11227 33642 11945 33646
rect 11997 33642 12011 33646
rect 12063 33642 12781 33694
rect 12833 33642 12847 33694
rect 12899 33642 13317 33694
rect 10258 33627 10286 33642
rect 10342 33627 13317 33642
rect 10258 33594 10273 33627
rect 10391 33614 11109 33627
rect 11161 33614 11175 33627
rect 11227 33614 11945 33627
rect 11997 33614 12011 33627
rect 9758 33575 10273 33594
rect 10325 33575 10339 33594
rect 10391 33575 10397 33614
rect 9758 33560 10397 33575
rect 9758 33558 10273 33560
rect 7883 33535 8601 33558
rect 7883 33508 7943 33535
rect 7251 33493 7943 33508
rect 7251 33470 7765 33493
rect 4539 33441 5257 33470
rect 5309 33441 5323 33470
rect 5375 33441 6093 33470
rect 6145 33441 6159 33470
rect 6211 33441 6929 33470
rect 6981 33441 6995 33470
rect 7047 33441 7765 33470
rect 7817 33441 7831 33493
rect 7883 33479 7943 33493
rect 7999 33526 8601 33535
rect 8653 33526 8667 33558
rect 8719 33526 9437 33558
rect 9489 33526 9503 33558
rect 9555 33526 10273 33558
rect 10325 33535 10339 33560
rect 10391 33558 10397 33560
rect 10453 33558 10477 33614
rect 10533 33558 10557 33614
rect 10613 33558 10637 33614
rect 10693 33558 10717 33614
rect 10773 33558 10797 33614
rect 10853 33558 10877 33614
rect 10933 33558 10957 33614
rect 11013 33558 11037 33614
rect 11093 33575 11109 33614
rect 11173 33575 11175 33614
rect 11093 33560 11117 33575
rect 11173 33560 11197 33575
rect 11093 33558 11109 33560
rect 11173 33558 11175 33560
rect 11253 33558 11277 33614
rect 11333 33558 11357 33614
rect 11413 33558 11437 33614
rect 11493 33558 11517 33614
rect 11573 33558 11597 33614
rect 11653 33558 11677 33614
rect 11733 33558 11758 33614
rect 11814 33558 11839 33614
rect 11895 33558 11920 33614
rect 11997 33575 12001 33614
rect 12063 33575 12781 33627
rect 12833 33575 12847 33627
rect 12899 33575 13317 33627
rect 11976 33560 12001 33575
rect 12057 33560 13317 33575
rect 11997 33558 12001 33560
rect 7999 33479 8041 33526
rect 7883 33470 8041 33479
rect 8097 33470 8124 33526
rect 8180 33470 8207 33526
rect 8263 33470 8290 33526
rect 8346 33470 8373 33526
rect 8429 33470 8456 33526
rect 8512 33470 8539 33526
rect 8595 33508 8601 33526
rect 8595 33493 8622 33508
rect 8678 33493 8705 33508
rect 8595 33470 8601 33493
rect 8761 33470 8788 33526
rect 8844 33470 8871 33526
rect 8927 33470 8954 33526
rect 9010 33470 9037 33526
rect 9093 33470 9120 33526
rect 9176 33470 9203 33526
rect 9259 33470 9286 33526
rect 9342 33470 9369 33526
rect 9425 33508 9437 33526
rect 9425 33493 9452 33508
rect 9508 33493 9535 33508
rect 9425 33470 9437 33493
rect 9591 33470 9618 33526
rect 9674 33470 9702 33526
rect 9758 33508 10273 33526
rect 10391 33526 11109 33558
rect 11161 33526 11175 33558
rect 11227 33526 11945 33558
rect 11997 33526 12011 33558
rect 10391 33508 10397 33526
rect 9758 33493 10307 33508
rect 10363 33493 10397 33508
rect 9758 33470 10273 33493
rect 7883 33441 8601 33470
rect 8653 33441 8667 33470
rect 8719 33441 9437 33470
rect 9489 33441 9503 33470
rect 9555 33441 10273 33470
rect 10325 33441 10339 33479
rect 10391 33470 10397 33493
rect 10453 33470 10477 33526
rect 10533 33470 10557 33526
rect 10613 33470 10637 33526
rect 10693 33470 10717 33526
rect 10773 33470 10797 33526
rect 10853 33470 10877 33526
rect 10933 33470 10957 33526
rect 11013 33470 11037 33526
rect 11093 33508 11109 33526
rect 11173 33508 11175 33526
rect 11093 33493 11117 33508
rect 11173 33493 11197 33508
rect 11093 33470 11109 33493
rect 11173 33470 11175 33493
rect 11253 33470 11277 33526
rect 11333 33470 11357 33526
rect 11413 33470 11437 33526
rect 11493 33470 11517 33526
rect 11573 33470 11597 33526
rect 11653 33470 11677 33526
rect 11733 33470 11758 33526
rect 11814 33470 11839 33526
rect 11895 33470 11920 33526
rect 11997 33508 12001 33526
rect 12063 33508 12781 33560
rect 12833 33508 12847 33560
rect 12899 33508 13317 33560
rect 11976 33493 12001 33508
rect 12057 33493 13317 33508
rect 11997 33470 12001 33493
rect 10391 33441 11109 33470
rect 11161 33441 11175 33470
rect 11227 33441 11945 33470
rect 11997 33441 12011 33470
rect 12063 33441 12781 33493
rect 12833 33441 12847 33493
rect 12899 33441 13317 33493
rect 3504 33438 13317 33441
rect 3504 33426 5216 33438
rect 5272 33426 5299 33438
rect 5355 33426 5382 33438
rect 3504 33370 3513 33426
rect 3569 33374 3585 33426
rect 3650 33374 3651 33426
rect 3569 33370 3594 33374
rect 3650 33370 3675 33374
rect 3731 33370 3757 33426
rect 3813 33370 3839 33426
rect 3895 33370 3921 33426
rect 3977 33370 4003 33426
rect 4059 33370 4085 33426
rect 4141 33370 4167 33426
rect 4223 33370 4249 33426
rect 4305 33374 4421 33426
rect 4473 33374 4487 33426
rect 4539 33382 5216 33426
rect 5375 33382 5382 33426
rect 5438 33382 5465 33438
rect 5521 33382 5548 33438
rect 5604 33382 5631 33438
rect 5687 33382 5714 33438
rect 5770 33382 5797 33438
rect 5853 33382 5880 33438
rect 5936 33382 5963 33438
rect 6019 33382 6046 33438
rect 6102 33426 6129 33438
rect 6185 33426 6211 33438
rect 6267 33382 6293 33438
rect 6349 33382 6375 33438
rect 6431 33382 6457 33438
rect 6513 33382 6539 33438
rect 6595 33382 6621 33438
rect 6677 33382 6703 33438
rect 6759 33382 6785 33438
rect 6841 33382 6867 33438
rect 6923 33426 6949 33438
rect 7005 33426 7031 33438
rect 6923 33382 6929 33426
rect 7087 33382 7113 33438
rect 7169 33382 7195 33438
rect 7251 33426 8041 33438
rect 7251 33382 7765 33426
rect 4539 33374 5257 33382
rect 5309 33374 5323 33382
rect 5375 33374 6093 33382
rect 6145 33374 6159 33382
rect 6211 33374 6929 33382
rect 6981 33374 6995 33382
rect 7047 33374 7765 33382
rect 7817 33374 7831 33426
rect 7883 33382 8041 33426
rect 8097 33382 8124 33438
rect 8180 33382 8207 33438
rect 8263 33382 8290 33438
rect 8346 33382 8373 33438
rect 8429 33382 8456 33438
rect 8512 33382 8539 33438
rect 8595 33426 8622 33438
rect 8678 33426 8705 33438
rect 8595 33382 8601 33426
rect 8761 33382 8788 33438
rect 8844 33382 8871 33438
rect 8927 33382 8954 33438
rect 9010 33382 9037 33438
rect 9093 33382 9120 33438
rect 9176 33382 9203 33438
rect 9259 33382 9286 33438
rect 9342 33382 9369 33438
rect 9425 33426 9452 33438
rect 9508 33426 9535 33438
rect 9425 33382 9437 33426
rect 9591 33382 9618 33438
rect 9674 33382 9702 33438
rect 9758 33426 10397 33438
rect 9758 33382 10273 33426
rect 7883 33374 8601 33382
rect 8653 33374 8667 33382
rect 8719 33374 9437 33382
rect 9489 33374 9503 33382
rect 9555 33374 10273 33382
rect 10325 33374 10339 33426
rect 10391 33382 10397 33426
rect 10453 33382 10477 33438
rect 10533 33382 10557 33438
rect 10613 33382 10637 33438
rect 10693 33382 10717 33438
rect 10773 33382 10797 33438
rect 10853 33382 10877 33438
rect 10933 33382 10957 33438
rect 11013 33382 11037 33438
rect 11093 33426 11117 33438
rect 11173 33426 11197 33438
rect 11093 33382 11109 33426
rect 11173 33382 11175 33426
rect 11253 33382 11277 33438
rect 11333 33382 11357 33438
rect 11413 33382 11437 33438
rect 11493 33382 11517 33438
rect 11573 33382 11597 33438
rect 11653 33382 11677 33438
rect 11733 33382 11758 33438
rect 11814 33382 11839 33438
rect 11895 33382 11920 33438
rect 11976 33426 12001 33438
rect 12057 33426 13317 33438
rect 11997 33382 12001 33426
rect 10391 33374 11109 33382
rect 11161 33374 11175 33382
rect 11227 33374 11945 33382
rect 11997 33374 12011 33382
rect 12063 33374 12781 33426
rect 12833 33374 12847 33426
rect 12899 33374 13317 33426
rect 4305 33370 13317 33374
rect 3504 33368 13317 33370
rect 100 33344 2792 33356
rect 100 33292 2249 33344
rect 2301 33292 2315 33344
rect 2367 33292 2792 33344
rect 100 33280 2792 33292
rect 100 33228 2249 33280
rect 2301 33228 2315 33280
rect 2367 33228 2792 33280
rect 100 33216 2792 33228
rect 100 33164 2249 33216
rect 2301 33164 2315 33216
rect 2367 33164 2792 33216
rect 100 33152 2792 33164
rect 100 33100 2249 33152
rect 2301 33100 2315 33152
rect 2367 33100 2792 33152
rect 100 33088 2792 33100
rect 100 33036 2249 33088
rect 2301 33036 2315 33088
rect 2367 33036 2792 33088
rect 100 33024 2792 33036
rect 100 32972 2249 33024
rect 2301 32972 2315 33024
rect 2367 32972 2792 33024
rect 100 32960 2792 32972
rect 100 32908 2249 32960
rect 2301 32908 2315 32960
rect 2367 32908 2792 32960
rect 100 32896 2792 32908
rect 100 32844 2249 32896
rect 2301 32844 2315 32896
rect 2367 32844 2792 32896
rect 100 32832 2792 32844
rect 100 32780 2249 32832
rect 2301 32780 2315 32832
rect 2367 32780 2792 32832
rect 100 32768 2792 32780
rect 100 32716 2249 32768
rect 2301 32716 2315 32768
rect 2367 32726 2792 32768
tri 2792 32726 3002 32936 sw
rect 2367 32720 13602 32726
rect 2367 32716 3167 32720
rect 100 32704 3167 32716
rect 100 32652 2249 32704
rect 2301 32652 2315 32704
rect 2367 32668 3167 32704
rect 3219 32668 3233 32720
rect 3285 32668 4003 32720
rect 4055 32668 4069 32720
rect 4121 32668 4839 32720
rect 4891 32668 4905 32720
rect 4957 32668 5675 32720
rect 5727 32668 5741 32720
rect 5793 32668 6511 32720
rect 6563 32668 6577 32720
rect 6629 32668 7347 32720
rect 7399 32668 7413 32720
rect 7465 32668 8183 32720
rect 8235 32668 8249 32720
rect 8301 32668 9019 32720
rect 9071 32668 9085 32720
rect 9137 32668 9855 32720
rect 9907 32668 9921 32720
rect 9973 32668 10691 32720
rect 10743 32668 10757 32720
rect 10809 32668 11527 32720
rect 11579 32668 11593 32720
rect 11645 32668 12363 32720
rect 12415 32668 12429 32720
rect 12481 32668 13200 32720
rect 13252 32668 13270 32720
rect 13322 32668 13340 32720
rect 13392 32668 13410 32720
rect 13462 32668 13480 32720
rect 13532 32668 13550 32720
rect 2367 32654 13602 32668
rect 2367 32652 3167 32654
rect 100 32640 3167 32652
rect 100 32588 2249 32640
rect 2301 32588 2315 32640
rect 2367 32602 3167 32640
rect 3219 32602 3233 32654
rect 3285 32602 4003 32654
rect 4055 32602 4069 32654
rect 4121 32602 4839 32654
rect 4891 32602 4905 32654
rect 4957 32602 5675 32654
rect 5727 32602 5741 32654
rect 5793 32602 6511 32654
rect 6563 32602 6577 32654
rect 6629 32602 7347 32654
rect 7399 32602 7413 32654
rect 7465 32602 8183 32654
rect 8235 32602 8249 32654
rect 8301 32602 9019 32654
rect 9071 32602 9085 32654
rect 9137 32602 9855 32654
rect 9907 32602 9921 32654
rect 9973 32602 10691 32654
rect 10743 32602 10757 32654
rect 10809 32602 11527 32654
rect 11579 32602 11593 32654
rect 11645 32602 12363 32654
rect 12415 32602 12429 32654
rect 12481 32602 13200 32654
rect 13252 32602 13270 32654
rect 13322 32602 13340 32654
rect 13392 32602 13410 32654
rect 13462 32602 13480 32654
rect 13532 32602 13550 32654
rect 2367 32588 13602 32602
rect 100 32576 3167 32588
rect 100 32524 2249 32576
rect 2301 32524 2315 32576
rect 2367 32536 3167 32576
rect 3219 32536 3233 32588
rect 3285 32536 4003 32588
rect 4055 32536 4069 32588
rect 4121 32536 4839 32588
rect 4891 32536 4905 32588
rect 4957 32536 5675 32588
rect 5727 32536 5741 32588
rect 5793 32536 6511 32588
rect 6563 32536 6577 32588
rect 6629 32536 7347 32588
rect 7399 32536 7413 32588
rect 7465 32536 8183 32588
rect 8235 32536 8249 32588
rect 8301 32536 9019 32588
rect 9071 32536 9085 32588
rect 9137 32536 9855 32588
rect 9907 32536 9921 32588
rect 9973 32536 10691 32588
rect 10743 32536 10757 32588
rect 10809 32536 11527 32588
rect 11579 32536 11593 32588
rect 11645 32536 12363 32588
rect 12415 32536 12429 32588
rect 12481 32536 13200 32588
rect 13252 32536 13270 32588
rect 13322 32536 13340 32588
rect 13392 32536 13410 32588
rect 13462 32536 13480 32588
rect 13532 32536 13550 32588
rect 2367 32524 13602 32536
rect 100 32522 13602 32524
rect 100 32512 3167 32522
rect 100 32460 2249 32512
rect 2301 32460 2315 32512
rect 2367 32470 3167 32512
rect 3219 32470 3233 32522
rect 3285 32470 4003 32522
rect 4055 32470 4069 32522
rect 4121 32470 4839 32522
rect 4891 32470 4905 32522
rect 4957 32470 5675 32522
rect 5727 32470 5741 32522
rect 5793 32470 6511 32522
rect 6563 32470 6577 32522
rect 6629 32470 7347 32522
rect 7399 32470 7413 32522
rect 7465 32470 8183 32522
rect 8235 32470 8249 32522
rect 8301 32470 9019 32522
rect 9071 32470 9085 32522
rect 9137 32470 9855 32522
rect 9907 32470 9921 32522
rect 9973 32470 10691 32522
rect 10743 32470 10757 32522
rect 10809 32470 11527 32522
rect 11579 32470 11593 32522
rect 11645 32470 12363 32522
rect 12415 32470 12429 32522
rect 12481 32470 13200 32522
rect 13252 32470 13270 32522
rect 13322 32470 13340 32522
rect 13392 32470 13410 32522
rect 13462 32470 13480 32522
rect 13532 32470 13550 32522
rect 2367 32460 13602 32470
rect 100 32456 13602 32460
rect 100 32448 3167 32456
rect 100 32396 2249 32448
rect 2301 32396 2315 32448
rect 2367 32404 3167 32448
rect 3219 32404 3233 32456
rect 3285 32404 4003 32456
rect 4055 32404 4069 32456
rect 4121 32404 4839 32456
rect 4891 32404 4905 32456
rect 4957 32404 5675 32456
rect 5727 32404 5741 32456
rect 5793 32404 6511 32456
rect 6563 32404 6577 32456
rect 6629 32404 7347 32456
rect 7399 32404 7413 32456
rect 7465 32404 8183 32456
rect 8235 32404 8249 32456
rect 8301 32404 9019 32456
rect 9071 32404 9085 32456
rect 9137 32404 9855 32456
rect 9907 32404 9921 32456
rect 9973 32404 10691 32456
rect 10743 32404 10757 32456
rect 10809 32404 11527 32456
rect 11579 32404 11593 32456
rect 11645 32404 12363 32456
rect 12415 32404 12429 32456
rect 12481 32404 13200 32456
rect 13252 32404 13270 32456
rect 13322 32404 13340 32456
rect 13392 32404 13410 32456
rect 13462 32404 13480 32456
rect 13532 32404 13550 32456
rect 2367 32396 13602 32404
rect 100 32390 13602 32396
rect 100 32384 3167 32390
rect 100 32332 2249 32384
rect 2301 32332 2315 32384
rect 2367 32338 3167 32384
rect 3219 32338 3233 32390
rect 3285 32338 4003 32390
rect 4055 32338 4069 32390
rect 4121 32338 4839 32390
rect 4891 32338 4905 32390
rect 4957 32338 5675 32390
rect 5727 32338 5741 32390
rect 5793 32338 6511 32390
rect 6563 32338 6577 32390
rect 6629 32338 7347 32390
rect 7399 32338 7413 32390
rect 7465 32338 8183 32390
rect 8235 32338 8249 32390
rect 8301 32338 9019 32390
rect 9071 32338 9085 32390
rect 9137 32338 9855 32390
rect 9907 32338 9921 32390
rect 9973 32338 10691 32390
rect 10743 32338 10757 32390
rect 10809 32338 11527 32390
rect 11579 32338 11593 32390
rect 11645 32338 12363 32390
rect 12415 32338 12429 32390
rect 12481 32338 13200 32390
rect 13252 32338 13270 32390
rect 13322 32338 13340 32390
rect 13392 32338 13410 32390
rect 13462 32338 13480 32390
rect 13532 32338 13550 32390
rect 2367 32332 13602 32338
rect 100 32323 13602 32332
rect 100 32319 3167 32323
rect 100 32267 2249 32319
rect 2301 32267 2315 32319
rect 2367 32271 3167 32319
rect 3219 32271 3233 32323
rect 3285 32271 4003 32323
rect 4055 32271 4069 32323
rect 4121 32271 4839 32323
rect 4891 32271 4905 32323
rect 4957 32271 5675 32323
rect 5727 32271 5741 32323
rect 5793 32271 6511 32323
rect 6563 32271 6577 32323
rect 6629 32271 7347 32323
rect 7399 32271 7413 32323
rect 7465 32271 8183 32323
rect 8235 32271 8249 32323
rect 8301 32271 9019 32323
rect 9071 32271 9085 32323
rect 9137 32271 9855 32323
rect 9907 32271 9921 32323
rect 9973 32271 10691 32323
rect 10743 32271 10757 32323
rect 10809 32271 11527 32323
rect 11579 32271 11593 32323
rect 11645 32271 12363 32323
rect 12415 32271 12429 32323
rect 12481 32271 13200 32323
rect 13252 32271 13270 32323
rect 13322 32271 13340 32323
rect 13392 32271 13410 32323
rect 13462 32271 13480 32323
rect 13532 32271 13550 32323
rect 2367 32267 13602 32271
rect 100 32256 13602 32267
rect 100 32254 3167 32256
rect 100 32202 2249 32254
rect 2301 32202 2315 32254
rect 2367 32204 3167 32254
rect 3219 32204 3233 32256
rect 3285 32204 4003 32256
rect 4055 32204 4069 32256
rect 4121 32204 4839 32256
rect 4891 32204 4905 32256
rect 4957 32204 5675 32256
rect 5727 32204 5741 32256
rect 5793 32204 6511 32256
rect 6563 32204 6577 32256
rect 6629 32204 7347 32256
rect 7399 32204 7413 32256
rect 7465 32204 8183 32256
rect 8235 32204 8249 32256
rect 8301 32204 9019 32256
rect 9071 32204 9085 32256
rect 9137 32204 9855 32256
rect 9907 32204 9921 32256
rect 9973 32204 10691 32256
rect 10743 32204 10757 32256
rect 10809 32204 11527 32256
rect 11579 32204 11593 32256
rect 11645 32204 12363 32256
rect 12415 32204 12429 32256
rect 12481 32204 13200 32256
rect 13252 32204 13270 32256
rect 13322 32204 13340 32256
rect 13392 32204 13410 32256
rect 13462 32204 13480 32256
rect 13532 32204 13550 32256
rect 2367 32202 13602 32204
rect 100 32198 13602 32202
rect 100 32189 2792 32198
rect 100 32137 2249 32189
rect 2301 32137 2315 32189
rect 2367 32137 2792 32189
rect 100 32124 2792 32137
rect 100 32072 2249 32124
rect 2301 32072 2315 32124
rect 2367 32072 2792 32124
rect 100 32059 2792 32072
rect 100 32007 2249 32059
rect 2301 32007 2315 32059
rect 2367 32007 2792 32059
rect 100 31994 2792 32007
rect 100 31942 2249 31994
rect 2301 31942 2315 31994
rect 2367 31942 2792 31994
tri 2792 31988 3002 32198 nw
rect 100 31929 2792 31942
rect 100 31877 2249 31929
rect 2301 31877 2315 31929
rect 2367 31877 2792 31929
rect 100 31864 2792 31877
rect 100 31812 2249 31864
rect 2301 31812 2315 31864
rect 2367 31812 2792 31864
rect 100 31799 2792 31812
rect 100 31747 2249 31799
rect 2301 31747 2315 31799
rect 2367 31747 2792 31799
rect 100 31734 2792 31747
rect 100 31682 2249 31734
rect 2301 31682 2315 31734
rect 2367 31682 2792 31734
rect 100 31669 2792 31682
rect 100 31617 2249 31669
rect 2301 31617 2315 31669
rect 2367 31617 2792 31669
rect 100 31604 2792 31617
rect 100 31552 2249 31604
rect 2301 31552 2315 31604
rect 2367 31552 2792 31604
rect 100 31539 2792 31552
rect 100 31487 2249 31539
rect 2301 31487 2315 31539
rect 2367 31487 2792 31539
rect 100 31474 2792 31487
rect 100 31422 2249 31474
rect 2301 31422 2315 31474
rect 2367 31422 2792 31474
rect 100 31409 2792 31422
rect 100 31357 2249 31409
rect 2301 31357 2315 31409
rect 2367 31357 2792 31409
rect 3504 31896 13317 31898
rect 3504 31840 3513 31896
rect 3569 31892 3596 31896
rect 3652 31892 3679 31896
rect 3569 31840 3585 31892
rect 3735 31840 3762 31896
rect 3818 31840 3845 31896
rect 3901 31840 3928 31896
rect 3984 31840 4011 31896
rect 4067 31840 4094 31896
rect 4150 31840 4177 31896
rect 4233 31840 4260 31896
rect 4316 31892 13317 31896
rect 4316 31840 4421 31892
rect 4473 31840 4487 31892
rect 4539 31883 5257 31892
rect 5309 31883 5323 31892
rect 5375 31883 6093 31892
rect 6145 31883 6159 31892
rect 6211 31883 6929 31892
rect 4539 31840 5215 31883
rect 5375 31840 5377 31883
rect 3504 31827 5215 31840
rect 5271 31827 5296 31840
rect 5352 31827 5377 31840
rect 5433 31827 5458 31883
rect 5514 31827 5539 31883
rect 5595 31827 5620 31883
rect 5676 31827 5701 31883
rect 5757 31827 5782 31883
rect 5838 31827 5863 31883
rect 5919 31827 5944 31883
rect 6000 31827 6025 31883
rect 6081 31840 6093 31883
rect 6081 31827 6106 31840
rect 6162 31827 6186 31840
rect 6242 31827 6266 31883
rect 6322 31827 6346 31883
rect 6402 31840 6929 31883
rect 6981 31840 6995 31892
rect 7047 31840 7765 31892
rect 7817 31840 7831 31892
rect 7883 31883 8601 31892
rect 8653 31883 8667 31892
rect 8719 31883 9437 31892
rect 9489 31883 9503 31892
rect 9555 31883 10273 31892
rect 7883 31840 8572 31883
rect 8719 31840 8732 31883
rect 6402 31827 8572 31840
rect 8628 31827 8652 31840
rect 8708 31827 8732 31840
rect 8788 31827 8812 31883
rect 8868 31827 8893 31883
rect 8949 31827 8974 31883
rect 9030 31827 9055 31883
rect 9111 31827 9136 31883
rect 9192 31827 9217 31883
rect 9273 31827 9298 31883
rect 9354 31827 9379 31883
rect 9435 31840 9437 31883
rect 9435 31827 9460 31840
rect 9516 31827 9541 31840
rect 9597 31827 9622 31883
rect 9678 31827 9703 31883
rect 9759 31840 10273 31883
rect 10325 31840 10339 31892
rect 10391 31883 11109 31892
rect 11161 31883 11175 31892
rect 11227 31883 11945 31892
rect 11997 31883 12011 31892
rect 10391 31840 10871 31883
rect 9759 31827 10871 31840
rect 10927 31827 10951 31883
rect 11007 31827 11031 31883
rect 11087 31840 11109 31883
rect 11167 31840 11175 31883
rect 11087 31827 11111 31840
rect 11167 31827 11192 31840
rect 11248 31827 11273 31883
rect 11329 31827 11354 31883
rect 11410 31827 11435 31883
rect 11491 31827 11516 31883
rect 11572 31827 11597 31883
rect 11653 31827 11678 31883
rect 11734 31827 11759 31883
rect 11815 31827 11840 31883
rect 11896 31827 11921 31883
rect 11997 31840 12002 31883
rect 12063 31840 12781 31892
rect 12833 31840 12847 31892
rect 12899 31840 13317 31892
rect 11977 31827 12002 31840
rect 12058 31827 13317 31840
rect 3504 31826 13317 31827
rect 3504 31802 3585 31826
rect 3637 31802 3651 31826
rect 3703 31802 4421 31826
rect 3504 31746 3513 31802
rect 3569 31774 3585 31802
rect 3569 31760 3596 31774
rect 3652 31760 3679 31774
rect 3569 31746 3585 31760
rect 3735 31746 3762 31802
rect 3818 31746 3845 31802
rect 3901 31746 3928 31802
rect 3984 31746 4011 31802
rect 4067 31746 4094 31802
rect 4150 31746 4177 31802
rect 4233 31746 4260 31802
rect 4316 31774 4421 31802
rect 4473 31774 4487 31826
rect 4539 31795 5257 31826
rect 5309 31795 5323 31826
rect 5375 31795 6093 31826
rect 6145 31795 6159 31826
rect 6211 31795 6929 31826
rect 4539 31774 5215 31795
rect 5375 31774 5377 31795
rect 4316 31760 5215 31774
rect 5271 31760 5296 31774
rect 5352 31760 5377 31774
rect 4316 31746 4421 31760
rect 3504 31708 3585 31746
rect 3637 31708 3651 31746
rect 3703 31708 4421 31746
rect 4473 31708 4487 31760
rect 4539 31739 5215 31760
rect 5375 31739 5377 31760
rect 5433 31739 5458 31795
rect 5514 31739 5539 31795
rect 5595 31739 5620 31795
rect 5676 31739 5701 31795
rect 5757 31739 5782 31795
rect 5838 31739 5863 31795
rect 5919 31739 5944 31795
rect 6000 31739 6025 31795
rect 6081 31774 6093 31795
rect 6081 31760 6106 31774
rect 6162 31760 6186 31774
rect 6081 31739 6093 31760
rect 6242 31739 6266 31795
rect 6322 31739 6346 31795
rect 6402 31774 6929 31795
rect 6981 31774 6995 31826
rect 7047 31774 7765 31826
rect 7817 31774 7831 31826
rect 7883 31795 8601 31826
rect 8653 31795 8667 31826
rect 8719 31795 9437 31826
rect 9489 31795 9503 31826
rect 9555 31795 10273 31826
rect 7883 31774 8572 31795
rect 8719 31774 8732 31795
rect 6402 31760 8572 31774
rect 8628 31760 8652 31774
rect 8708 31760 8732 31774
rect 6402 31739 6929 31760
rect 4539 31708 5257 31739
rect 5309 31708 5323 31739
rect 5375 31708 6093 31739
rect 6145 31708 6159 31739
rect 6211 31708 6929 31739
rect 6981 31708 6995 31760
rect 7047 31708 7765 31760
rect 7817 31708 7831 31760
rect 7883 31739 8572 31760
rect 8719 31739 8732 31760
rect 8788 31739 8812 31795
rect 8868 31739 8893 31795
rect 8949 31739 8974 31795
rect 9030 31739 9055 31795
rect 9111 31739 9136 31795
rect 9192 31739 9217 31795
rect 9273 31739 9298 31795
rect 9354 31739 9379 31795
rect 9435 31774 9437 31795
rect 9435 31760 9460 31774
rect 9516 31760 9541 31774
rect 9435 31739 9437 31760
rect 9597 31739 9622 31795
rect 9678 31739 9703 31795
rect 9759 31774 10273 31795
rect 10325 31774 10339 31826
rect 10391 31795 11109 31826
rect 11161 31795 11175 31826
rect 11227 31795 11945 31826
rect 11997 31795 12011 31826
rect 10391 31774 10871 31795
rect 9759 31760 10871 31774
rect 9759 31739 10273 31760
rect 7883 31708 8601 31739
rect 8653 31708 8667 31739
rect 8719 31708 9437 31739
rect 9489 31708 9503 31739
rect 9555 31708 10273 31739
rect 10325 31708 10339 31760
rect 10391 31739 10871 31760
rect 10927 31739 10951 31795
rect 11007 31739 11031 31795
rect 11087 31774 11109 31795
rect 11167 31774 11175 31795
rect 11087 31760 11111 31774
rect 11167 31760 11192 31774
rect 11087 31739 11109 31760
rect 11167 31739 11175 31760
rect 11248 31739 11273 31795
rect 11329 31739 11354 31795
rect 11410 31739 11435 31795
rect 11491 31739 11516 31795
rect 11572 31739 11597 31795
rect 11653 31739 11678 31795
rect 11734 31739 11759 31795
rect 11815 31739 11840 31795
rect 11896 31739 11921 31795
rect 11997 31774 12002 31795
rect 12063 31774 12781 31826
rect 12833 31774 12847 31826
rect 12899 31774 13317 31826
rect 11977 31760 12002 31774
rect 12058 31760 13317 31774
rect 11997 31739 12002 31760
rect 10391 31708 11109 31739
rect 11161 31708 11175 31739
rect 11227 31708 11945 31739
rect 11997 31708 12011 31739
rect 12063 31708 12781 31760
rect 12833 31708 12847 31760
rect 12899 31708 13317 31760
rect 3504 31652 3513 31708
rect 3569 31694 3596 31708
rect 3652 31694 3679 31708
rect 3569 31652 3585 31694
rect 3735 31652 3762 31708
rect 3818 31652 3845 31708
rect 3901 31652 3928 31708
rect 3984 31652 4011 31708
rect 4067 31652 4094 31708
rect 4150 31652 4177 31708
rect 4233 31652 4260 31708
rect 4316 31707 13317 31708
rect 4316 31694 5215 31707
rect 5271 31694 5296 31707
rect 5352 31694 5377 31707
rect 4316 31652 4421 31694
rect 3504 31642 3585 31652
rect 3637 31642 3651 31652
rect 3703 31642 4421 31652
rect 4473 31642 4487 31694
rect 4539 31651 5215 31694
rect 5375 31651 5377 31694
rect 5433 31651 5458 31707
rect 5514 31651 5539 31707
rect 5595 31651 5620 31707
rect 5676 31651 5701 31707
rect 5757 31651 5782 31707
rect 5838 31651 5863 31707
rect 5919 31651 5944 31707
rect 6000 31651 6025 31707
rect 6081 31694 6106 31707
rect 6162 31694 6186 31707
rect 6081 31651 6093 31694
rect 6242 31651 6266 31707
rect 6322 31651 6346 31707
rect 6402 31694 8572 31707
rect 8628 31694 8652 31707
rect 8708 31694 8732 31707
rect 6402 31651 6929 31694
rect 4539 31642 5257 31651
rect 5309 31642 5323 31651
rect 5375 31642 6093 31651
rect 6145 31642 6159 31651
rect 6211 31642 6929 31651
rect 6981 31642 6995 31694
rect 7047 31642 7765 31694
rect 7817 31642 7831 31694
rect 7883 31651 8572 31694
rect 8719 31651 8732 31694
rect 8788 31651 8812 31707
rect 8868 31651 8893 31707
rect 8949 31651 8974 31707
rect 9030 31651 9055 31707
rect 9111 31651 9136 31707
rect 9192 31651 9217 31707
rect 9273 31651 9298 31707
rect 9354 31651 9379 31707
rect 9435 31694 9460 31707
rect 9516 31694 9541 31707
rect 9435 31651 9437 31694
rect 9597 31651 9622 31707
rect 9678 31651 9703 31707
rect 9759 31694 10871 31707
rect 9759 31651 10273 31694
rect 7883 31642 8601 31651
rect 8653 31642 8667 31651
rect 8719 31642 9437 31651
rect 9489 31642 9503 31651
rect 9555 31642 10273 31651
rect 10325 31642 10339 31694
rect 10391 31651 10871 31694
rect 10927 31651 10951 31707
rect 11007 31651 11031 31707
rect 11087 31694 11111 31707
rect 11167 31694 11192 31707
rect 11087 31651 11109 31694
rect 11167 31651 11175 31694
rect 11248 31651 11273 31707
rect 11329 31651 11354 31707
rect 11410 31651 11435 31707
rect 11491 31651 11516 31707
rect 11572 31651 11597 31707
rect 11653 31651 11678 31707
rect 11734 31651 11759 31707
rect 11815 31651 11840 31707
rect 11896 31651 11921 31707
rect 11977 31694 12002 31707
rect 12058 31694 13317 31707
rect 11997 31651 12002 31694
rect 10391 31642 11109 31651
rect 11161 31642 11175 31651
rect 11227 31642 11945 31651
rect 11997 31642 12011 31651
rect 12063 31642 12781 31694
rect 12833 31642 12847 31694
rect 12899 31642 13317 31694
rect 3504 31627 13317 31642
rect 3504 31614 3585 31627
rect 3637 31614 3651 31627
rect 3703 31614 4421 31627
rect 3504 31558 3513 31614
rect 3569 31575 3585 31614
rect 3569 31560 3596 31575
rect 3652 31560 3679 31575
rect 3569 31558 3585 31560
rect 3735 31558 3762 31614
rect 3818 31558 3845 31614
rect 3901 31558 3928 31614
rect 3984 31558 4011 31614
rect 4067 31558 4094 31614
rect 4150 31558 4177 31614
rect 4233 31558 4260 31614
rect 4316 31575 4421 31614
rect 4473 31575 4487 31627
rect 4539 31619 5257 31627
rect 5309 31619 5323 31627
rect 5375 31619 6093 31627
rect 6145 31619 6159 31627
rect 6211 31619 6929 31627
rect 4539 31575 5215 31619
rect 5375 31575 5377 31619
rect 4316 31563 5215 31575
rect 5271 31563 5296 31575
rect 5352 31563 5377 31575
rect 5433 31563 5458 31619
rect 5514 31563 5539 31619
rect 5595 31563 5620 31619
rect 5676 31563 5701 31619
rect 5757 31563 5782 31619
rect 5838 31563 5863 31619
rect 5919 31563 5944 31619
rect 6000 31563 6025 31619
rect 6081 31575 6093 31619
rect 6081 31563 6106 31575
rect 6162 31563 6186 31575
rect 6242 31563 6266 31619
rect 6322 31563 6346 31619
rect 6402 31575 6929 31619
rect 6981 31575 6995 31627
rect 7047 31575 7765 31627
rect 7817 31575 7831 31627
rect 7883 31619 8601 31627
rect 8653 31619 8667 31627
rect 8719 31619 9437 31627
rect 9489 31619 9503 31627
rect 9555 31619 10273 31627
rect 7883 31575 8572 31619
rect 8719 31575 8732 31619
rect 6402 31563 8572 31575
rect 8628 31563 8652 31575
rect 8708 31563 8732 31575
rect 8788 31563 8812 31619
rect 8868 31563 8893 31619
rect 8949 31563 8974 31619
rect 9030 31563 9055 31619
rect 9111 31563 9136 31619
rect 9192 31563 9217 31619
rect 9273 31563 9298 31619
rect 9354 31563 9379 31619
rect 9435 31575 9437 31619
rect 9435 31563 9460 31575
rect 9516 31563 9541 31575
rect 9597 31563 9622 31619
rect 9678 31563 9703 31619
rect 9759 31575 10273 31619
rect 10325 31575 10339 31627
rect 10391 31619 11109 31627
rect 11161 31619 11175 31627
rect 11227 31619 11945 31627
rect 11997 31619 12011 31627
rect 10391 31575 10871 31619
rect 9759 31563 10871 31575
rect 10927 31563 10951 31619
rect 11007 31563 11031 31619
rect 11087 31575 11109 31619
rect 11167 31575 11175 31619
rect 11087 31563 11111 31575
rect 11167 31563 11192 31575
rect 11248 31563 11273 31619
rect 11329 31563 11354 31619
rect 11410 31563 11435 31619
rect 11491 31563 11516 31619
rect 11572 31563 11597 31619
rect 11653 31563 11678 31619
rect 11734 31563 11759 31619
rect 11815 31563 11840 31619
rect 11896 31563 11921 31619
rect 11997 31575 12002 31619
rect 12063 31575 12781 31627
rect 12833 31575 12847 31627
rect 12899 31575 13317 31627
rect 11977 31563 12002 31575
rect 12058 31563 13317 31575
rect 4316 31560 13317 31563
rect 4316 31558 4421 31560
rect 3504 31520 3585 31558
rect 3637 31520 3651 31558
rect 3703 31520 4421 31558
rect 3504 31464 3513 31520
rect 3569 31508 3585 31520
rect 3569 31493 3596 31508
rect 3652 31493 3679 31508
rect 3569 31464 3585 31493
rect 3735 31464 3762 31520
rect 3818 31464 3845 31520
rect 3901 31464 3928 31520
rect 3984 31464 4011 31520
rect 4067 31464 4094 31520
rect 4150 31464 4177 31520
rect 4233 31464 4260 31520
rect 4316 31508 4421 31520
rect 4473 31508 4487 31560
rect 4539 31531 5257 31560
rect 5309 31531 5323 31560
rect 5375 31531 6093 31560
rect 6145 31531 6159 31560
rect 6211 31531 6929 31560
rect 4539 31508 5215 31531
rect 5375 31508 5377 31531
rect 4316 31493 5215 31508
rect 5271 31493 5296 31508
rect 5352 31493 5377 31508
rect 4316 31464 4421 31493
rect 3504 31441 3585 31464
rect 3637 31441 3651 31464
rect 3703 31441 4421 31464
rect 4473 31441 4487 31493
rect 4539 31475 5215 31493
rect 5375 31475 5377 31493
rect 5433 31475 5458 31531
rect 5514 31475 5539 31531
rect 5595 31475 5620 31531
rect 5676 31475 5701 31531
rect 5757 31475 5782 31531
rect 5838 31475 5863 31531
rect 5919 31475 5944 31531
rect 6000 31475 6025 31531
rect 6081 31508 6093 31531
rect 6081 31493 6106 31508
rect 6162 31493 6186 31508
rect 6081 31475 6093 31493
rect 6242 31475 6266 31531
rect 6322 31475 6346 31531
rect 6402 31508 6929 31531
rect 6981 31508 6995 31560
rect 7047 31508 7765 31560
rect 7817 31508 7831 31560
rect 7883 31531 8601 31560
rect 8653 31531 8667 31560
rect 8719 31531 9437 31560
rect 9489 31531 9503 31560
rect 9555 31531 10273 31560
rect 7883 31508 8572 31531
rect 8719 31508 8732 31531
rect 6402 31493 8572 31508
rect 8628 31493 8652 31508
rect 8708 31493 8732 31508
rect 6402 31475 6929 31493
rect 4539 31443 5257 31475
rect 5309 31443 5323 31475
rect 5375 31443 6093 31475
rect 6145 31443 6159 31475
rect 6211 31443 6929 31475
rect 4539 31441 5215 31443
rect 5375 31441 5377 31443
rect 3504 31426 5215 31441
rect 5271 31426 5296 31441
rect 5352 31426 5377 31441
rect 3504 31370 3513 31426
rect 3569 31374 3585 31426
rect 3569 31370 3596 31374
rect 3652 31370 3679 31374
rect 3735 31370 3762 31426
rect 3818 31370 3845 31426
rect 3901 31370 3928 31426
rect 3984 31370 4011 31426
rect 4067 31370 4094 31426
rect 4150 31370 4177 31426
rect 4233 31370 4260 31426
rect 4316 31374 4421 31426
rect 4473 31374 4487 31426
rect 4539 31387 5215 31426
rect 5375 31387 5377 31426
rect 5433 31387 5458 31443
rect 5514 31387 5539 31443
rect 5595 31387 5620 31443
rect 5676 31387 5701 31443
rect 5757 31387 5782 31443
rect 5838 31387 5863 31443
rect 5919 31387 5944 31443
rect 6000 31387 6025 31443
rect 6081 31441 6093 31443
rect 6081 31426 6106 31441
rect 6162 31426 6186 31441
rect 6081 31387 6093 31426
rect 6242 31387 6266 31443
rect 6322 31387 6346 31443
rect 6402 31441 6929 31443
rect 6981 31441 6995 31493
rect 7047 31441 7765 31493
rect 7817 31441 7831 31493
rect 7883 31475 8572 31493
rect 8719 31475 8732 31493
rect 8788 31475 8812 31531
rect 8868 31475 8893 31531
rect 8949 31475 8974 31531
rect 9030 31475 9055 31531
rect 9111 31475 9136 31531
rect 9192 31475 9217 31531
rect 9273 31475 9298 31531
rect 9354 31475 9379 31531
rect 9435 31508 9437 31531
rect 9435 31493 9460 31508
rect 9516 31493 9541 31508
rect 9435 31475 9437 31493
rect 9597 31475 9622 31531
rect 9678 31475 9703 31531
rect 9759 31508 10273 31531
rect 10325 31508 10339 31560
rect 10391 31531 11109 31560
rect 11161 31531 11175 31560
rect 11227 31531 11945 31560
rect 11997 31531 12011 31560
rect 10391 31508 10871 31531
rect 9759 31493 10871 31508
rect 9759 31475 10273 31493
rect 7883 31443 8601 31475
rect 8653 31443 8667 31475
rect 8719 31443 9437 31475
rect 9489 31443 9503 31475
rect 9555 31443 10273 31475
rect 7883 31441 8572 31443
rect 8719 31441 8732 31443
rect 6402 31426 8572 31441
rect 8628 31426 8652 31441
rect 8708 31426 8732 31441
rect 6402 31387 6929 31426
rect 4539 31374 5257 31387
rect 5309 31374 5323 31387
rect 5375 31374 6093 31387
rect 6145 31374 6159 31387
rect 6211 31374 6929 31387
rect 6981 31374 6995 31426
rect 7047 31374 7765 31426
rect 7817 31374 7831 31426
rect 7883 31387 8572 31426
rect 8719 31387 8732 31426
rect 8788 31387 8812 31443
rect 8868 31387 8893 31443
rect 8949 31387 8974 31443
rect 9030 31387 9055 31443
rect 9111 31387 9136 31443
rect 9192 31387 9217 31443
rect 9273 31387 9298 31443
rect 9354 31387 9379 31443
rect 9435 31441 9437 31443
rect 9435 31426 9460 31441
rect 9516 31426 9541 31441
rect 9435 31387 9437 31426
rect 9597 31387 9622 31443
rect 9678 31387 9703 31443
rect 9759 31441 10273 31443
rect 10325 31441 10339 31493
rect 10391 31475 10871 31493
rect 10927 31475 10951 31531
rect 11007 31475 11031 31531
rect 11087 31508 11109 31531
rect 11167 31508 11175 31531
rect 11087 31493 11111 31508
rect 11167 31493 11192 31508
rect 11087 31475 11109 31493
rect 11167 31475 11175 31493
rect 11248 31475 11273 31531
rect 11329 31475 11354 31531
rect 11410 31475 11435 31531
rect 11491 31475 11516 31531
rect 11572 31475 11597 31531
rect 11653 31475 11678 31531
rect 11734 31475 11759 31531
rect 11815 31475 11840 31531
rect 11896 31475 11921 31531
rect 11997 31508 12002 31531
rect 12063 31508 12781 31560
rect 12833 31508 12847 31560
rect 12899 31508 13317 31560
rect 11977 31493 12002 31508
rect 12058 31493 13317 31508
rect 11997 31475 12002 31493
rect 10391 31443 11109 31475
rect 11161 31443 11175 31475
rect 11227 31443 11945 31475
rect 11997 31443 12011 31475
rect 10391 31441 10871 31443
rect 9759 31426 10871 31441
rect 9759 31387 10273 31426
rect 7883 31374 8601 31387
rect 8653 31374 8667 31387
rect 8719 31374 9437 31387
rect 9489 31374 9503 31387
rect 9555 31374 10273 31387
rect 10325 31374 10339 31426
rect 10391 31387 10871 31426
rect 10927 31387 10951 31443
rect 11007 31387 11031 31443
rect 11087 31441 11109 31443
rect 11167 31441 11175 31443
rect 11087 31426 11111 31441
rect 11167 31426 11192 31441
rect 11087 31387 11109 31426
rect 11167 31387 11175 31426
rect 11248 31387 11273 31443
rect 11329 31387 11354 31443
rect 11410 31387 11435 31443
rect 11491 31387 11516 31443
rect 11572 31387 11597 31443
rect 11653 31387 11678 31443
rect 11734 31387 11759 31443
rect 11815 31387 11840 31443
rect 11896 31387 11921 31443
rect 11997 31441 12002 31443
rect 12063 31441 12781 31493
rect 12833 31441 12847 31493
rect 12899 31441 13317 31493
rect 11977 31426 12002 31441
rect 12058 31426 13317 31441
rect 11997 31387 12002 31426
rect 10391 31374 11109 31387
rect 11161 31374 11175 31387
rect 11227 31374 11945 31387
rect 11997 31374 12011 31387
rect 12063 31374 12781 31426
rect 12833 31374 12847 31426
rect 12899 31374 13317 31426
rect 4316 31370 13317 31374
rect 3504 31368 13317 31370
rect 100 31344 2792 31357
rect 100 31292 2249 31344
rect 2301 31292 2315 31344
rect 2367 31292 2792 31344
rect 100 31279 2792 31292
rect 100 31227 2249 31279
rect 2301 31227 2315 31279
rect 2367 31227 2792 31279
rect 100 31214 2792 31227
rect 100 31162 2249 31214
rect 2301 31162 2315 31214
rect 2367 31162 2792 31214
rect 100 31149 2792 31162
rect 100 31097 2249 31149
rect 2301 31097 2315 31149
rect 2367 31097 2792 31149
rect 100 31084 2792 31097
rect 100 31032 2249 31084
rect 2301 31032 2315 31084
rect 2367 31032 2792 31084
rect 100 31019 2792 31032
rect 100 30967 2249 31019
rect 2301 30967 2315 31019
rect 2367 30967 2792 31019
rect 100 30954 2792 30967
rect 100 30902 2249 30954
rect 2301 30902 2315 30954
rect 2367 30902 2792 30954
rect 100 30889 2792 30902
rect 100 30837 2249 30889
rect 2301 30837 2315 30889
rect 2367 30837 2792 30889
rect 100 30824 2792 30837
rect 100 30772 2249 30824
rect 2301 30772 2315 30824
rect 2367 30772 2792 30824
rect 100 30759 2792 30772
rect 100 30707 2249 30759
rect 2301 30707 2315 30759
rect 2367 30726 2792 30759
tri 2792 30726 3002 30936 sw
rect 2367 30720 13602 30726
rect 2367 30707 3167 30720
rect 100 30694 3167 30707
rect 100 30642 2249 30694
rect 2301 30642 2315 30694
rect 2367 30668 3167 30694
rect 3219 30668 3233 30720
rect 3285 30668 4003 30720
rect 4055 30668 4069 30720
rect 4121 30668 4839 30720
rect 4891 30668 4905 30720
rect 4957 30668 5675 30720
rect 5727 30668 5741 30720
rect 5793 30668 6511 30720
rect 6563 30668 6577 30720
rect 6629 30668 7347 30720
rect 7399 30668 7413 30720
rect 7465 30668 8183 30720
rect 8235 30668 8249 30720
rect 8301 30668 9019 30720
rect 9071 30668 9085 30720
rect 9137 30668 9855 30720
rect 9907 30668 9921 30720
rect 9973 30668 10691 30720
rect 10743 30668 10757 30720
rect 10809 30668 11527 30720
rect 11579 30668 11593 30720
rect 11645 30668 12363 30720
rect 12415 30668 12429 30720
rect 12481 30668 13200 30720
rect 13252 30668 13270 30720
rect 13322 30668 13340 30720
rect 13392 30668 13410 30720
rect 13462 30668 13480 30720
rect 13532 30668 13550 30720
rect 2367 30654 13602 30668
rect 2367 30642 3167 30654
rect 100 30629 3167 30642
rect 100 30577 2249 30629
rect 2301 30577 2315 30629
rect 2367 30602 3167 30629
rect 3219 30602 3233 30654
rect 3285 30602 4003 30654
rect 4055 30602 4069 30654
rect 4121 30602 4839 30654
rect 4891 30602 4905 30654
rect 4957 30602 5675 30654
rect 5727 30602 5741 30654
rect 5793 30602 6511 30654
rect 6563 30602 6577 30654
rect 6629 30602 7347 30654
rect 7399 30602 7413 30654
rect 7465 30602 8183 30654
rect 8235 30602 8249 30654
rect 8301 30602 9019 30654
rect 9071 30602 9085 30654
rect 9137 30602 9855 30654
rect 9907 30602 9921 30654
rect 9973 30602 10691 30654
rect 10743 30602 10757 30654
rect 10809 30602 11527 30654
rect 11579 30602 11593 30654
rect 11645 30602 12363 30654
rect 12415 30602 12429 30654
rect 12481 30602 13200 30654
rect 13252 30602 13270 30654
rect 13322 30602 13340 30654
rect 13392 30602 13410 30654
rect 13462 30602 13480 30654
rect 13532 30602 13550 30654
rect 2367 30588 13602 30602
rect 2367 30577 3167 30588
rect 100 30564 3167 30577
rect 100 30512 2249 30564
rect 2301 30512 2315 30564
rect 2367 30536 3167 30564
rect 3219 30536 3233 30588
rect 3285 30536 4003 30588
rect 4055 30536 4069 30588
rect 4121 30536 4839 30588
rect 4891 30536 4905 30588
rect 4957 30536 5675 30588
rect 5727 30536 5741 30588
rect 5793 30536 6511 30588
rect 6563 30536 6577 30588
rect 6629 30536 7347 30588
rect 7399 30536 7413 30588
rect 7465 30536 8183 30588
rect 8235 30536 8249 30588
rect 8301 30536 9019 30588
rect 9071 30536 9085 30588
rect 9137 30536 9855 30588
rect 9907 30536 9921 30588
rect 9973 30536 10691 30588
rect 10743 30536 10757 30588
rect 10809 30536 11527 30588
rect 11579 30536 11593 30588
rect 11645 30536 12363 30588
rect 12415 30536 12429 30588
rect 12481 30536 13200 30588
rect 13252 30536 13270 30588
rect 13322 30536 13340 30588
rect 13392 30536 13410 30588
rect 13462 30536 13480 30588
rect 13532 30536 13550 30588
rect 2367 30522 13602 30536
rect 2367 30512 3167 30522
rect 100 30499 3167 30512
rect 100 30447 2249 30499
rect 2301 30447 2315 30499
rect 2367 30470 3167 30499
rect 3219 30470 3233 30522
rect 3285 30470 4003 30522
rect 4055 30470 4069 30522
rect 4121 30470 4839 30522
rect 4891 30470 4905 30522
rect 4957 30470 5675 30522
rect 5727 30470 5741 30522
rect 5793 30470 6511 30522
rect 6563 30470 6577 30522
rect 6629 30470 7347 30522
rect 7399 30470 7413 30522
rect 7465 30470 8183 30522
rect 8235 30470 8249 30522
rect 8301 30470 9019 30522
rect 9071 30470 9085 30522
rect 9137 30470 9855 30522
rect 9907 30470 9921 30522
rect 9973 30470 10691 30522
rect 10743 30470 10757 30522
rect 10809 30470 11527 30522
rect 11579 30470 11593 30522
rect 11645 30470 12363 30522
rect 12415 30470 12429 30522
rect 12481 30470 13200 30522
rect 13252 30470 13270 30522
rect 13322 30470 13340 30522
rect 13392 30470 13410 30522
rect 13462 30470 13480 30522
rect 13532 30470 13550 30522
rect 2367 30456 13602 30470
rect 2367 30447 3167 30456
rect 100 30434 3167 30447
rect 100 30382 2249 30434
rect 2301 30382 2315 30434
rect 2367 30404 3167 30434
rect 3219 30404 3233 30456
rect 3285 30404 4003 30456
rect 4055 30404 4069 30456
rect 4121 30404 4839 30456
rect 4891 30404 4905 30456
rect 4957 30404 5675 30456
rect 5727 30404 5741 30456
rect 5793 30404 6511 30456
rect 6563 30404 6577 30456
rect 6629 30404 7347 30456
rect 7399 30404 7413 30456
rect 7465 30404 8183 30456
rect 8235 30404 8249 30456
rect 8301 30404 9019 30456
rect 9071 30404 9085 30456
rect 9137 30404 9855 30456
rect 9907 30404 9921 30456
rect 9973 30404 10691 30456
rect 10743 30404 10757 30456
rect 10809 30404 11527 30456
rect 11579 30404 11593 30456
rect 11645 30404 12363 30456
rect 12415 30404 12429 30456
rect 12481 30404 13200 30456
rect 13252 30404 13270 30456
rect 13322 30404 13340 30456
rect 13392 30404 13410 30456
rect 13462 30404 13480 30456
rect 13532 30404 13550 30456
rect 2367 30390 13602 30404
rect 2367 30382 3167 30390
rect 100 30369 3167 30382
rect 100 30317 2249 30369
rect 2301 30317 2315 30369
rect 2367 30338 3167 30369
rect 3219 30338 3233 30390
rect 3285 30338 4003 30390
rect 4055 30338 4069 30390
rect 4121 30338 4839 30390
rect 4891 30338 4905 30390
rect 4957 30338 5675 30390
rect 5727 30338 5741 30390
rect 5793 30338 6511 30390
rect 6563 30338 6577 30390
rect 6629 30338 7347 30390
rect 7399 30338 7413 30390
rect 7465 30338 8183 30390
rect 8235 30338 8249 30390
rect 8301 30338 9019 30390
rect 9071 30338 9085 30390
rect 9137 30338 9855 30390
rect 9907 30338 9921 30390
rect 9973 30338 10691 30390
rect 10743 30338 10757 30390
rect 10809 30338 11527 30390
rect 11579 30338 11593 30390
rect 11645 30338 12363 30390
rect 12415 30338 12429 30390
rect 12481 30338 13200 30390
rect 13252 30338 13270 30390
rect 13322 30338 13340 30390
rect 13392 30338 13410 30390
rect 13462 30338 13480 30390
rect 13532 30338 13550 30390
rect 2367 30323 13602 30338
rect 2367 30317 3167 30323
rect 100 30304 3167 30317
rect 100 30252 2249 30304
rect 2301 30252 2315 30304
rect 2367 30271 3167 30304
rect 3219 30271 3233 30323
rect 3285 30271 4003 30323
rect 4055 30271 4069 30323
rect 4121 30271 4839 30323
rect 4891 30271 4905 30323
rect 4957 30271 5675 30323
rect 5727 30271 5741 30323
rect 5793 30271 6511 30323
rect 6563 30271 6577 30323
rect 6629 30271 7347 30323
rect 7399 30271 7413 30323
rect 7465 30271 8183 30323
rect 8235 30271 8249 30323
rect 8301 30271 9019 30323
rect 9071 30271 9085 30323
rect 9137 30271 9855 30323
rect 9907 30271 9921 30323
rect 9973 30271 10691 30323
rect 10743 30271 10757 30323
rect 10809 30271 11527 30323
rect 11579 30271 11593 30323
rect 11645 30271 12363 30323
rect 12415 30271 12429 30323
rect 12481 30271 13200 30323
rect 13252 30271 13270 30323
rect 13322 30271 13340 30323
rect 13392 30271 13410 30323
rect 13462 30271 13480 30323
rect 13532 30271 13550 30323
rect 2367 30256 13602 30271
rect 2367 30252 3167 30256
rect 100 30239 3167 30252
rect 100 30187 2249 30239
rect 2301 30187 2315 30239
rect 2367 30204 3167 30239
rect 3219 30204 3233 30256
rect 3285 30204 4003 30256
rect 4055 30204 4069 30256
rect 4121 30204 4839 30256
rect 4891 30204 4905 30256
rect 4957 30204 5675 30256
rect 5727 30204 5741 30256
rect 5793 30204 6511 30256
rect 6563 30204 6577 30256
rect 6629 30204 7347 30256
rect 7399 30204 7413 30256
rect 7465 30204 8183 30256
rect 8235 30204 8249 30256
rect 8301 30204 9019 30256
rect 9071 30204 9085 30256
rect 9137 30204 9855 30256
rect 9907 30204 9921 30256
rect 9973 30204 10691 30256
rect 10743 30204 10757 30256
rect 10809 30204 11527 30256
rect 11579 30204 11593 30256
rect 11645 30204 12363 30256
rect 12415 30204 12429 30256
rect 12481 30204 13200 30256
rect 13252 30204 13270 30256
rect 13322 30204 13340 30256
rect 13392 30204 13410 30256
rect 13462 30204 13480 30256
rect 13532 30204 13550 30256
rect 2367 30198 13602 30204
rect 2367 30187 2792 30198
rect 100 30174 2792 30187
rect 100 30122 2249 30174
rect 2301 30122 2315 30174
rect 2367 30122 2792 30174
rect 100 30109 2792 30122
rect 100 30057 2249 30109
rect 2301 30057 2315 30109
rect 2367 30057 2792 30109
rect 100 30044 2792 30057
rect 100 29992 2249 30044
rect 2301 29992 2315 30044
rect 2367 29992 2792 30044
rect 100 29979 2792 29992
tri 2792 29988 3002 30198 nw
rect 100 29927 2249 29979
rect 2301 29927 2315 29979
rect 2367 29927 2792 29979
rect 100 29914 2792 29927
rect 100 29862 2249 29914
rect 2301 29862 2315 29914
rect 2367 29862 2792 29914
rect 100 29849 2792 29862
rect 100 29797 2249 29849
rect 2301 29797 2315 29849
rect 2367 29797 2792 29849
rect 100 29784 2792 29797
rect 100 29732 2249 29784
rect 2301 29732 2315 29784
rect 2367 29732 2792 29784
rect 100 29719 2792 29732
rect 100 29667 2249 29719
rect 2301 29667 2315 29719
rect 2367 29667 2792 29719
rect 100 29654 2792 29667
rect 100 29602 2249 29654
rect 2301 29602 2315 29654
rect 2367 29602 2792 29654
rect 100 29589 2792 29602
rect 100 29537 2249 29589
rect 2301 29537 2315 29589
rect 2367 29537 2792 29589
rect 100 29524 2792 29537
rect 100 29472 2249 29524
rect 2301 29472 2315 29524
rect 2367 29472 2792 29524
rect 100 29459 2792 29472
rect 100 29407 2249 29459
rect 2301 29407 2315 29459
rect 2367 29407 2792 29459
rect 100 29394 2792 29407
rect 100 29342 2249 29394
rect 2301 29342 2315 29394
rect 2367 29342 2792 29394
rect 3504 29896 13317 29898
rect 3504 29840 3513 29896
rect 3569 29892 3596 29896
rect 3652 29892 3679 29896
rect 3569 29840 3585 29892
rect 3735 29840 3762 29896
rect 3818 29840 3845 29896
rect 3901 29840 3928 29896
rect 3984 29840 4011 29896
rect 4067 29840 4094 29896
rect 4150 29840 4177 29896
rect 4233 29840 4260 29896
rect 4316 29892 13317 29896
rect 4316 29840 4421 29892
rect 4473 29840 4487 29892
rect 4539 29883 5257 29892
rect 5309 29883 5323 29892
rect 5375 29883 6093 29892
rect 6145 29883 6159 29892
rect 6211 29883 6929 29892
rect 4539 29840 5215 29883
rect 5375 29840 5377 29883
rect 3504 29827 5215 29840
rect 5271 29827 5296 29840
rect 5352 29827 5377 29840
rect 5433 29827 5458 29883
rect 5514 29827 5539 29883
rect 5595 29827 5620 29883
rect 5676 29827 5701 29883
rect 5757 29827 5782 29883
rect 5838 29827 5863 29883
rect 5919 29827 5944 29883
rect 6000 29827 6025 29883
rect 6081 29840 6093 29883
rect 6081 29827 6106 29840
rect 6162 29827 6186 29840
rect 6242 29827 6266 29883
rect 6322 29827 6346 29883
rect 6402 29840 6929 29883
rect 6981 29840 6995 29892
rect 7047 29840 7765 29892
rect 7817 29840 7831 29892
rect 7883 29883 8601 29892
rect 8653 29883 8667 29892
rect 8719 29883 9437 29892
rect 9489 29883 9503 29892
rect 9555 29883 10273 29892
rect 7883 29840 8572 29883
rect 8719 29840 8732 29883
rect 6402 29827 8572 29840
rect 8628 29827 8652 29840
rect 8708 29827 8732 29840
rect 8788 29827 8812 29883
rect 8868 29827 8893 29883
rect 8949 29827 8974 29883
rect 9030 29827 9055 29883
rect 9111 29827 9136 29883
rect 9192 29827 9217 29883
rect 9273 29827 9298 29883
rect 9354 29827 9379 29883
rect 9435 29840 9437 29883
rect 9435 29827 9460 29840
rect 9516 29827 9541 29840
rect 9597 29827 9622 29883
rect 9678 29827 9703 29883
rect 9759 29840 10273 29883
rect 10325 29840 10339 29892
rect 10391 29883 11109 29892
rect 11161 29883 11175 29892
rect 11227 29883 11945 29892
rect 11997 29883 12011 29892
rect 10391 29840 10871 29883
rect 9759 29827 10871 29840
rect 10927 29827 10951 29883
rect 11007 29827 11031 29883
rect 11087 29840 11109 29883
rect 11167 29840 11175 29883
rect 11087 29827 11111 29840
rect 11167 29827 11192 29840
rect 11248 29827 11273 29883
rect 11329 29827 11354 29883
rect 11410 29827 11435 29883
rect 11491 29827 11516 29883
rect 11572 29827 11597 29883
rect 11653 29827 11678 29883
rect 11734 29827 11759 29883
rect 11815 29827 11840 29883
rect 11896 29827 11921 29883
rect 11997 29840 12002 29883
rect 12063 29840 12781 29892
rect 12833 29840 12847 29892
rect 12899 29840 13317 29892
rect 11977 29827 12002 29840
rect 12058 29827 13317 29840
rect 3504 29826 13317 29827
rect 3504 29802 3585 29826
rect 3637 29802 3651 29826
rect 3703 29802 4421 29826
rect 3504 29746 3513 29802
rect 3569 29774 3585 29802
rect 3569 29760 3596 29774
rect 3652 29760 3679 29774
rect 3569 29746 3585 29760
rect 3735 29746 3762 29802
rect 3818 29746 3845 29802
rect 3901 29746 3928 29802
rect 3984 29746 4011 29802
rect 4067 29746 4094 29802
rect 4150 29746 4177 29802
rect 4233 29746 4260 29802
rect 4316 29774 4421 29802
rect 4473 29774 4487 29826
rect 4539 29795 5257 29826
rect 5309 29795 5323 29826
rect 5375 29795 6093 29826
rect 6145 29795 6159 29826
rect 6211 29795 6929 29826
rect 4539 29774 5215 29795
rect 5375 29774 5377 29795
rect 4316 29760 5215 29774
rect 5271 29760 5296 29774
rect 5352 29760 5377 29774
rect 4316 29746 4421 29760
rect 3504 29708 3585 29746
rect 3637 29708 3651 29746
rect 3703 29708 4421 29746
rect 4473 29708 4487 29760
rect 4539 29739 5215 29760
rect 5375 29739 5377 29760
rect 5433 29739 5458 29795
rect 5514 29739 5539 29795
rect 5595 29739 5620 29795
rect 5676 29739 5701 29795
rect 5757 29739 5782 29795
rect 5838 29739 5863 29795
rect 5919 29739 5944 29795
rect 6000 29739 6025 29795
rect 6081 29774 6093 29795
rect 6081 29760 6106 29774
rect 6162 29760 6186 29774
rect 6081 29739 6093 29760
rect 6242 29739 6266 29795
rect 6322 29739 6346 29795
rect 6402 29774 6929 29795
rect 6981 29774 6995 29826
rect 7047 29774 7765 29826
rect 7817 29774 7831 29826
rect 7883 29795 8601 29826
rect 8653 29795 8667 29826
rect 8719 29795 9437 29826
rect 9489 29795 9503 29826
rect 9555 29795 10273 29826
rect 7883 29774 8572 29795
rect 8719 29774 8732 29795
rect 6402 29760 8572 29774
rect 8628 29760 8652 29774
rect 8708 29760 8732 29774
rect 6402 29739 6929 29760
rect 4539 29708 5257 29739
rect 5309 29708 5323 29739
rect 5375 29708 6093 29739
rect 6145 29708 6159 29739
rect 6211 29708 6929 29739
rect 6981 29708 6995 29760
rect 7047 29708 7765 29760
rect 7817 29708 7831 29760
rect 7883 29739 8572 29760
rect 8719 29739 8732 29760
rect 8788 29739 8812 29795
rect 8868 29739 8893 29795
rect 8949 29739 8974 29795
rect 9030 29739 9055 29795
rect 9111 29739 9136 29795
rect 9192 29739 9217 29795
rect 9273 29739 9298 29795
rect 9354 29739 9379 29795
rect 9435 29774 9437 29795
rect 9435 29760 9460 29774
rect 9516 29760 9541 29774
rect 9435 29739 9437 29760
rect 9597 29739 9622 29795
rect 9678 29739 9703 29795
rect 9759 29774 10273 29795
rect 10325 29774 10339 29826
rect 10391 29795 11109 29826
rect 11161 29795 11175 29826
rect 11227 29795 11945 29826
rect 11997 29795 12011 29826
rect 10391 29774 10871 29795
rect 9759 29760 10871 29774
rect 9759 29739 10273 29760
rect 7883 29708 8601 29739
rect 8653 29708 8667 29739
rect 8719 29708 9437 29739
rect 9489 29708 9503 29739
rect 9555 29708 10273 29739
rect 10325 29708 10339 29760
rect 10391 29739 10871 29760
rect 10927 29739 10951 29795
rect 11007 29739 11031 29795
rect 11087 29774 11109 29795
rect 11167 29774 11175 29795
rect 11087 29760 11111 29774
rect 11167 29760 11192 29774
rect 11087 29739 11109 29760
rect 11167 29739 11175 29760
rect 11248 29739 11273 29795
rect 11329 29739 11354 29795
rect 11410 29739 11435 29795
rect 11491 29739 11516 29795
rect 11572 29739 11597 29795
rect 11653 29739 11678 29795
rect 11734 29739 11759 29795
rect 11815 29739 11840 29795
rect 11896 29739 11921 29795
rect 11997 29774 12002 29795
rect 12063 29774 12781 29826
rect 12833 29774 12847 29826
rect 12899 29774 13317 29826
rect 11977 29760 12002 29774
rect 12058 29760 13317 29774
rect 11997 29739 12002 29760
rect 10391 29708 11109 29739
rect 11161 29708 11175 29739
rect 11227 29708 11945 29739
rect 11997 29708 12011 29739
rect 12063 29708 12781 29760
rect 12833 29708 12847 29760
rect 12899 29708 13317 29760
rect 3504 29652 3513 29708
rect 3569 29694 3596 29708
rect 3652 29694 3679 29708
rect 3569 29652 3585 29694
rect 3735 29652 3762 29708
rect 3818 29652 3845 29708
rect 3901 29652 3928 29708
rect 3984 29652 4011 29708
rect 4067 29652 4094 29708
rect 4150 29652 4177 29708
rect 4233 29652 4260 29708
rect 4316 29707 13317 29708
rect 4316 29694 5215 29707
rect 5271 29694 5296 29707
rect 5352 29694 5377 29707
rect 4316 29652 4421 29694
rect 3504 29642 3585 29652
rect 3637 29642 3651 29652
rect 3703 29642 4421 29652
rect 4473 29642 4487 29694
rect 4539 29651 5215 29694
rect 5375 29651 5377 29694
rect 5433 29651 5458 29707
rect 5514 29651 5539 29707
rect 5595 29651 5620 29707
rect 5676 29651 5701 29707
rect 5757 29651 5782 29707
rect 5838 29651 5863 29707
rect 5919 29651 5944 29707
rect 6000 29651 6025 29707
rect 6081 29694 6106 29707
rect 6162 29694 6186 29707
rect 6081 29651 6093 29694
rect 6242 29651 6266 29707
rect 6322 29651 6346 29707
rect 6402 29694 8572 29707
rect 8628 29694 8652 29707
rect 8708 29694 8732 29707
rect 6402 29651 6929 29694
rect 4539 29642 5257 29651
rect 5309 29642 5323 29651
rect 5375 29642 6093 29651
rect 6145 29642 6159 29651
rect 6211 29642 6929 29651
rect 6981 29642 6995 29694
rect 7047 29642 7765 29694
rect 7817 29642 7831 29694
rect 7883 29651 8572 29694
rect 8719 29651 8732 29694
rect 8788 29651 8812 29707
rect 8868 29651 8893 29707
rect 8949 29651 8974 29707
rect 9030 29651 9055 29707
rect 9111 29651 9136 29707
rect 9192 29651 9217 29707
rect 9273 29651 9298 29707
rect 9354 29651 9379 29707
rect 9435 29694 9460 29707
rect 9516 29694 9541 29707
rect 9435 29651 9437 29694
rect 9597 29651 9622 29707
rect 9678 29651 9703 29707
rect 9759 29694 10871 29707
rect 9759 29651 10273 29694
rect 7883 29642 8601 29651
rect 8653 29642 8667 29651
rect 8719 29642 9437 29651
rect 9489 29642 9503 29651
rect 9555 29642 10273 29651
rect 10325 29642 10339 29694
rect 10391 29651 10871 29694
rect 10927 29651 10951 29707
rect 11007 29651 11031 29707
rect 11087 29694 11111 29707
rect 11167 29694 11192 29707
rect 11087 29651 11109 29694
rect 11167 29651 11175 29694
rect 11248 29651 11273 29707
rect 11329 29651 11354 29707
rect 11410 29651 11435 29707
rect 11491 29651 11516 29707
rect 11572 29651 11597 29707
rect 11653 29651 11678 29707
rect 11734 29651 11759 29707
rect 11815 29651 11840 29707
rect 11896 29651 11921 29707
rect 11977 29694 12002 29707
rect 12058 29694 13317 29707
rect 11997 29651 12002 29694
rect 10391 29642 11109 29651
rect 11161 29642 11175 29651
rect 11227 29642 11945 29651
rect 11997 29642 12011 29651
rect 12063 29642 12781 29694
rect 12833 29642 12847 29694
rect 12899 29642 13317 29694
rect 3504 29627 13317 29642
rect 3504 29614 3585 29627
rect 3637 29614 3651 29627
rect 3703 29614 4421 29627
rect 3504 29558 3513 29614
rect 3569 29575 3585 29614
rect 3569 29560 3596 29575
rect 3652 29560 3679 29575
rect 3569 29558 3585 29560
rect 3735 29558 3762 29614
rect 3818 29558 3845 29614
rect 3901 29558 3928 29614
rect 3984 29558 4011 29614
rect 4067 29558 4094 29614
rect 4150 29558 4177 29614
rect 4233 29558 4260 29614
rect 4316 29575 4421 29614
rect 4473 29575 4487 29627
rect 4539 29619 5257 29627
rect 5309 29619 5323 29627
rect 5375 29619 6093 29627
rect 6145 29619 6159 29627
rect 6211 29619 6929 29627
rect 4539 29575 5215 29619
rect 5375 29575 5377 29619
rect 4316 29563 5215 29575
rect 5271 29563 5296 29575
rect 5352 29563 5377 29575
rect 5433 29563 5458 29619
rect 5514 29563 5539 29619
rect 5595 29563 5620 29619
rect 5676 29563 5701 29619
rect 5757 29563 5782 29619
rect 5838 29563 5863 29619
rect 5919 29563 5944 29619
rect 6000 29563 6025 29619
rect 6081 29575 6093 29619
rect 6081 29563 6106 29575
rect 6162 29563 6186 29575
rect 6242 29563 6266 29619
rect 6322 29563 6346 29619
rect 6402 29575 6929 29619
rect 6981 29575 6995 29627
rect 7047 29575 7765 29627
rect 7817 29575 7831 29627
rect 7883 29619 8601 29627
rect 8653 29619 8667 29627
rect 8719 29619 9437 29627
rect 9489 29619 9503 29627
rect 9555 29619 10273 29627
rect 7883 29575 8572 29619
rect 8719 29575 8732 29619
rect 6402 29563 8572 29575
rect 8628 29563 8652 29575
rect 8708 29563 8732 29575
rect 8788 29563 8812 29619
rect 8868 29563 8893 29619
rect 8949 29563 8974 29619
rect 9030 29563 9055 29619
rect 9111 29563 9136 29619
rect 9192 29563 9217 29619
rect 9273 29563 9298 29619
rect 9354 29563 9379 29619
rect 9435 29575 9437 29619
rect 9435 29563 9460 29575
rect 9516 29563 9541 29575
rect 9597 29563 9622 29619
rect 9678 29563 9703 29619
rect 9759 29575 10273 29619
rect 10325 29575 10339 29627
rect 10391 29619 11109 29627
rect 11161 29619 11175 29627
rect 11227 29619 11945 29627
rect 11997 29619 12011 29627
rect 10391 29575 10871 29619
rect 9759 29563 10871 29575
rect 10927 29563 10951 29619
rect 11007 29563 11031 29619
rect 11087 29575 11109 29619
rect 11167 29575 11175 29619
rect 11087 29563 11111 29575
rect 11167 29563 11192 29575
rect 11248 29563 11273 29619
rect 11329 29563 11354 29619
rect 11410 29563 11435 29619
rect 11491 29563 11516 29619
rect 11572 29563 11597 29619
rect 11653 29563 11678 29619
rect 11734 29563 11759 29619
rect 11815 29563 11840 29619
rect 11896 29563 11921 29619
rect 11997 29575 12002 29619
rect 12063 29575 12781 29627
rect 12833 29575 12847 29627
rect 12899 29575 13317 29627
rect 11977 29563 12002 29575
rect 12058 29563 13317 29575
rect 4316 29560 13317 29563
rect 4316 29558 4421 29560
rect 3504 29520 3585 29558
rect 3637 29520 3651 29558
rect 3703 29520 4421 29558
rect 3504 29464 3513 29520
rect 3569 29508 3585 29520
rect 3569 29493 3596 29508
rect 3652 29493 3679 29508
rect 3569 29464 3585 29493
rect 3735 29464 3762 29520
rect 3818 29464 3845 29520
rect 3901 29464 3928 29520
rect 3984 29464 4011 29520
rect 4067 29464 4094 29520
rect 4150 29464 4177 29520
rect 4233 29464 4260 29520
rect 4316 29508 4421 29520
rect 4473 29508 4487 29560
rect 4539 29531 5257 29560
rect 5309 29531 5323 29560
rect 5375 29531 6093 29560
rect 6145 29531 6159 29560
rect 6211 29531 6929 29560
rect 4539 29508 5215 29531
rect 5375 29508 5377 29531
rect 4316 29493 5215 29508
rect 5271 29493 5296 29508
rect 5352 29493 5377 29508
rect 4316 29464 4421 29493
rect 3504 29441 3585 29464
rect 3637 29441 3651 29464
rect 3703 29441 4421 29464
rect 4473 29441 4487 29493
rect 4539 29475 5215 29493
rect 5375 29475 5377 29493
rect 5433 29475 5458 29531
rect 5514 29475 5539 29531
rect 5595 29475 5620 29531
rect 5676 29475 5701 29531
rect 5757 29475 5782 29531
rect 5838 29475 5863 29531
rect 5919 29475 5944 29531
rect 6000 29475 6025 29531
rect 6081 29508 6093 29531
rect 6081 29493 6106 29508
rect 6162 29493 6186 29508
rect 6081 29475 6093 29493
rect 6242 29475 6266 29531
rect 6322 29475 6346 29531
rect 6402 29508 6929 29531
rect 6981 29508 6995 29560
rect 7047 29508 7765 29560
rect 7817 29508 7831 29560
rect 7883 29531 8601 29560
rect 8653 29531 8667 29560
rect 8719 29531 9437 29560
rect 9489 29531 9503 29560
rect 9555 29531 10273 29560
rect 7883 29508 8572 29531
rect 8719 29508 8732 29531
rect 6402 29493 8572 29508
rect 8628 29493 8652 29508
rect 8708 29493 8732 29508
rect 6402 29475 6929 29493
rect 4539 29443 5257 29475
rect 5309 29443 5323 29475
rect 5375 29443 6093 29475
rect 6145 29443 6159 29475
rect 6211 29443 6929 29475
rect 4539 29441 5215 29443
rect 5375 29441 5377 29443
rect 3504 29426 5215 29441
rect 5271 29426 5296 29441
rect 5352 29426 5377 29441
rect 3504 29370 3513 29426
rect 3569 29374 3585 29426
rect 3569 29370 3596 29374
rect 3652 29370 3679 29374
rect 3735 29370 3762 29426
rect 3818 29370 3845 29426
rect 3901 29370 3928 29426
rect 3984 29370 4011 29426
rect 4067 29370 4094 29426
rect 4150 29370 4177 29426
rect 4233 29370 4260 29426
rect 4316 29374 4421 29426
rect 4473 29374 4487 29426
rect 4539 29387 5215 29426
rect 5375 29387 5377 29426
rect 5433 29387 5458 29443
rect 5514 29387 5539 29443
rect 5595 29387 5620 29443
rect 5676 29387 5701 29443
rect 5757 29387 5782 29443
rect 5838 29387 5863 29443
rect 5919 29387 5944 29443
rect 6000 29387 6025 29443
rect 6081 29441 6093 29443
rect 6081 29426 6106 29441
rect 6162 29426 6186 29441
rect 6081 29387 6093 29426
rect 6242 29387 6266 29443
rect 6322 29387 6346 29443
rect 6402 29441 6929 29443
rect 6981 29441 6995 29493
rect 7047 29441 7765 29493
rect 7817 29441 7831 29493
rect 7883 29475 8572 29493
rect 8719 29475 8732 29493
rect 8788 29475 8812 29531
rect 8868 29475 8893 29531
rect 8949 29475 8974 29531
rect 9030 29475 9055 29531
rect 9111 29475 9136 29531
rect 9192 29475 9217 29531
rect 9273 29475 9298 29531
rect 9354 29475 9379 29531
rect 9435 29508 9437 29531
rect 9435 29493 9460 29508
rect 9516 29493 9541 29508
rect 9435 29475 9437 29493
rect 9597 29475 9622 29531
rect 9678 29475 9703 29531
rect 9759 29508 10273 29531
rect 10325 29508 10339 29560
rect 10391 29531 11109 29560
rect 11161 29531 11175 29560
rect 11227 29531 11945 29560
rect 11997 29531 12011 29560
rect 10391 29508 10871 29531
rect 9759 29493 10871 29508
rect 9759 29475 10273 29493
rect 7883 29443 8601 29475
rect 8653 29443 8667 29475
rect 8719 29443 9437 29475
rect 9489 29443 9503 29475
rect 9555 29443 10273 29475
rect 7883 29441 8572 29443
rect 8719 29441 8732 29443
rect 6402 29426 8572 29441
rect 8628 29426 8652 29441
rect 8708 29426 8732 29441
rect 6402 29387 6929 29426
rect 4539 29374 5257 29387
rect 5309 29374 5323 29387
rect 5375 29374 6093 29387
rect 6145 29374 6159 29387
rect 6211 29374 6929 29387
rect 6981 29374 6995 29426
rect 7047 29374 7765 29426
rect 7817 29374 7831 29426
rect 7883 29387 8572 29426
rect 8719 29387 8732 29426
rect 8788 29387 8812 29443
rect 8868 29387 8893 29443
rect 8949 29387 8974 29443
rect 9030 29387 9055 29443
rect 9111 29387 9136 29443
rect 9192 29387 9217 29443
rect 9273 29387 9298 29443
rect 9354 29387 9379 29443
rect 9435 29441 9437 29443
rect 9435 29426 9460 29441
rect 9516 29426 9541 29441
rect 9435 29387 9437 29426
rect 9597 29387 9622 29443
rect 9678 29387 9703 29443
rect 9759 29441 10273 29443
rect 10325 29441 10339 29493
rect 10391 29475 10871 29493
rect 10927 29475 10951 29531
rect 11007 29475 11031 29531
rect 11087 29508 11109 29531
rect 11167 29508 11175 29531
rect 11087 29493 11111 29508
rect 11167 29493 11192 29508
rect 11087 29475 11109 29493
rect 11167 29475 11175 29493
rect 11248 29475 11273 29531
rect 11329 29475 11354 29531
rect 11410 29475 11435 29531
rect 11491 29475 11516 29531
rect 11572 29475 11597 29531
rect 11653 29475 11678 29531
rect 11734 29475 11759 29531
rect 11815 29475 11840 29531
rect 11896 29475 11921 29531
rect 11997 29508 12002 29531
rect 12063 29508 12781 29560
rect 12833 29508 12847 29560
rect 12899 29508 13317 29560
rect 11977 29493 12002 29508
rect 12058 29493 13317 29508
rect 11997 29475 12002 29493
rect 10391 29443 11109 29475
rect 11161 29443 11175 29475
rect 11227 29443 11945 29475
rect 11997 29443 12011 29475
rect 10391 29441 10871 29443
rect 9759 29426 10871 29441
rect 9759 29387 10273 29426
rect 7883 29374 8601 29387
rect 8653 29374 8667 29387
rect 8719 29374 9437 29387
rect 9489 29374 9503 29387
rect 9555 29374 10273 29387
rect 10325 29374 10339 29426
rect 10391 29387 10871 29426
rect 10927 29387 10951 29443
rect 11007 29387 11031 29443
rect 11087 29441 11109 29443
rect 11167 29441 11175 29443
rect 11087 29426 11111 29441
rect 11167 29426 11192 29441
rect 11087 29387 11109 29426
rect 11167 29387 11175 29426
rect 11248 29387 11273 29443
rect 11329 29387 11354 29443
rect 11410 29387 11435 29443
rect 11491 29387 11516 29443
rect 11572 29387 11597 29443
rect 11653 29387 11678 29443
rect 11734 29387 11759 29443
rect 11815 29387 11840 29443
rect 11896 29387 11921 29443
rect 11997 29441 12002 29443
rect 12063 29441 12781 29493
rect 12833 29441 12847 29493
rect 12899 29441 13317 29493
rect 11977 29426 12002 29441
rect 12058 29426 13317 29441
rect 11997 29387 12002 29426
rect 10391 29374 11109 29387
rect 11161 29374 11175 29387
rect 11227 29374 11945 29387
rect 11997 29374 12011 29387
rect 12063 29374 12781 29426
rect 12833 29374 12847 29426
rect 12899 29374 13317 29426
rect 4316 29370 13317 29374
rect 3504 29368 13317 29370
rect 100 29329 2792 29342
rect 100 29277 2249 29329
rect 2301 29277 2315 29329
rect 2367 29277 2792 29329
rect 100 29264 2792 29277
rect 100 29212 2249 29264
rect 2301 29212 2315 29264
rect 2367 29212 2792 29264
rect 100 29199 2792 29212
rect 100 29147 2249 29199
rect 2301 29147 2315 29199
rect 2367 29147 2792 29199
rect 100 29134 2792 29147
rect 100 29082 2249 29134
rect 2301 29082 2315 29134
rect 2367 29082 2792 29134
rect 100 29069 2792 29082
rect 100 29017 2249 29069
rect 2301 29017 2315 29069
rect 2367 29017 2792 29069
rect 100 29004 2792 29017
rect 100 28952 2249 29004
rect 2301 28952 2315 29004
rect 2367 28952 2792 29004
rect 100 28939 2792 28952
rect 100 28887 2249 28939
rect 2301 28887 2315 28939
rect 2367 28887 2792 28939
rect 100 28726 2792 28887
tri 2792 28726 3002 28936 sw
rect 100 28720 13602 28726
rect 100 28668 4839 28720
rect 4891 28668 4905 28720
rect 4957 28668 5675 28720
rect 5727 28668 5741 28720
rect 5793 28668 6511 28720
rect 6563 28668 6577 28720
rect 6629 28668 7347 28720
rect 7399 28668 7413 28720
rect 7465 28668 8183 28720
rect 8235 28668 8249 28720
rect 8301 28668 9019 28720
rect 9071 28668 9085 28720
rect 9137 28668 9855 28720
rect 9907 28668 9921 28720
rect 9973 28668 10691 28720
rect 10743 28668 10757 28720
rect 10809 28668 11527 28720
rect 11579 28668 11593 28720
rect 11645 28668 12363 28720
rect 12415 28668 12429 28720
rect 12481 28668 13200 28720
rect 13252 28668 13270 28720
rect 13322 28668 13340 28720
rect 13392 28668 13410 28720
rect 13462 28668 13480 28720
rect 13532 28668 13550 28720
rect 100 28654 13602 28668
rect 100 28602 4839 28654
rect 4891 28602 4905 28654
rect 4957 28602 5675 28654
rect 5727 28602 5741 28654
rect 5793 28602 6511 28654
rect 6563 28602 6577 28654
rect 6629 28602 7347 28654
rect 7399 28602 7413 28654
rect 7465 28602 8183 28654
rect 8235 28602 8249 28654
rect 8301 28602 9019 28654
rect 9071 28602 9085 28654
rect 9137 28602 9855 28654
rect 9907 28602 9921 28654
rect 9973 28602 10691 28654
rect 10743 28602 10757 28654
rect 10809 28602 11527 28654
rect 11579 28602 11593 28654
rect 11645 28602 12363 28654
rect 12415 28602 12429 28654
rect 12481 28602 13200 28654
rect 13252 28602 13270 28654
rect 13322 28602 13340 28654
rect 13392 28602 13410 28654
rect 13462 28602 13480 28654
rect 13532 28602 13550 28654
rect 100 28588 13602 28602
rect 100 28536 4839 28588
rect 4891 28536 4905 28588
rect 4957 28536 5675 28588
rect 5727 28536 5741 28588
rect 5793 28536 6511 28588
rect 6563 28536 6577 28588
rect 6629 28536 7347 28588
rect 7399 28536 7413 28588
rect 7465 28536 8183 28588
rect 8235 28536 8249 28588
rect 8301 28536 9019 28588
rect 9071 28536 9085 28588
rect 9137 28536 9855 28588
rect 9907 28536 9921 28588
rect 9973 28536 10691 28588
rect 10743 28536 10757 28588
rect 10809 28536 11527 28588
rect 11579 28536 11593 28588
rect 11645 28536 12363 28588
rect 12415 28536 12429 28588
rect 12481 28536 13200 28588
rect 13252 28536 13270 28588
rect 13322 28536 13340 28588
rect 13392 28536 13410 28588
rect 13462 28536 13480 28588
rect 13532 28536 13550 28588
rect 100 28522 13602 28536
rect 100 28470 4839 28522
rect 4891 28470 4905 28522
rect 4957 28470 5675 28522
rect 5727 28470 5741 28522
rect 5793 28470 6511 28522
rect 6563 28470 6577 28522
rect 6629 28470 7347 28522
rect 7399 28470 7413 28522
rect 7465 28470 8183 28522
rect 8235 28470 8249 28522
rect 8301 28470 9019 28522
rect 9071 28470 9085 28522
rect 9137 28470 9855 28522
rect 9907 28470 9921 28522
rect 9973 28470 10691 28522
rect 10743 28470 10757 28522
rect 10809 28470 11527 28522
rect 11579 28470 11593 28522
rect 11645 28470 12363 28522
rect 12415 28470 12429 28522
rect 12481 28470 13200 28522
rect 13252 28470 13270 28522
rect 13322 28470 13340 28522
rect 13392 28470 13410 28522
rect 13462 28470 13480 28522
rect 13532 28470 13550 28522
rect 100 28456 13602 28470
rect 100 28404 4839 28456
rect 4891 28404 4905 28456
rect 4957 28404 5675 28456
rect 5727 28404 5741 28456
rect 5793 28404 6511 28456
rect 6563 28404 6577 28456
rect 6629 28404 7347 28456
rect 7399 28404 7413 28456
rect 7465 28404 8183 28456
rect 8235 28404 8249 28456
rect 8301 28404 9019 28456
rect 9071 28404 9085 28456
rect 9137 28404 9855 28456
rect 9907 28404 9921 28456
rect 9973 28404 10691 28456
rect 10743 28404 10757 28456
rect 10809 28404 11527 28456
rect 11579 28404 11593 28456
rect 11645 28404 12363 28456
rect 12415 28404 12429 28456
rect 12481 28404 13200 28456
rect 13252 28404 13270 28456
rect 13322 28404 13340 28456
rect 13392 28404 13410 28456
rect 13462 28404 13480 28456
rect 13532 28404 13550 28456
rect 100 28390 13602 28404
rect 100 28338 4839 28390
rect 4891 28338 4905 28390
rect 4957 28338 5675 28390
rect 5727 28338 5741 28390
rect 5793 28338 6511 28390
rect 6563 28338 6577 28390
rect 6629 28338 7347 28390
rect 7399 28338 7413 28390
rect 7465 28338 8183 28390
rect 8235 28338 8249 28390
rect 8301 28338 9019 28390
rect 9071 28338 9085 28390
rect 9137 28338 9855 28390
rect 9907 28338 9921 28390
rect 9973 28338 10691 28390
rect 10743 28338 10757 28390
rect 10809 28338 11527 28390
rect 11579 28338 11593 28390
rect 11645 28338 12363 28390
rect 12415 28338 12429 28390
rect 12481 28338 13200 28390
rect 13252 28338 13270 28390
rect 13322 28338 13340 28390
rect 13392 28338 13410 28390
rect 13462 28338 13480 28390
rect 13532 28338 13550 28390
rect 100 28323 13602 28338
rect 100 28271 4839 28323
rect 4891 28271 4905 28323
rect 4957 28271 5675 28323
rect 5727 28271 5741 28323
rect 5793 28271 6511 28323
rect 6563 28271 6577 28323
rect 6629 28271 7347 28323
rect 7399 28271 7413 28323
rect 7465 28271 8183 28323
rect 8235 28271 8249 28323
rect 8301 28271 9019 28323
rect 9071 28271 9085 28323
rect 9137 28271 9855 28323
rect 9907 28271 9921 28323
rect 9973 28271 10691 28323
rect 10743 28271 10757 28323
rect 10809 28271 11527 28323
rect 11579 28271 11593 28323
rect 11645 28271 12363 28323
rect 12415 28271 12429 28323
rect 12481 28271 13200 28323
rect 13252 28271 13270 28323
rect 13322 28271 13340 28323
rect 13392 28271 13410 28323
rect 13462 28271 13480 28323
rect 13532 28271 13550 28323
rect 100 28256 13602 28271
rect 100 28204 4839 28256
rect 4891 28204 4905 28256
rect 4957 28204 5675 28256
rect 5727 28204 5741 28256
rect 5793 28204 6511 28256
rect 6563 28204 6577 28256
rect 6629 28204 7347 28256
rect 7399 28204 7413 28256
rect 7465 28204 8183 28256
rect 8235 28204 8249 28256
rect 8301 28204 9019 28256
rect 9071 28204 9085 28256
rect 9137 28204 9855 28256
rect 9907 28204 9921 28256
rect 9973 28204 10691 28256
rect 10743 28204 10757 28256
rect 10809 28204 11527 28256
rect 11579 28204 11593 28256
rect 11645 28204 12363 28256
rect 12415 28204 12429 28256
rect 12481 28204 13200 28256
rect 13252 28204 13270 28256
rect 13322 28204 13340 28256
rect 13392 28204 13410 28256
rect 13462 28204 13480 28256
rect 13532 28204 13550 28256
rect 100 28198 13602 28204
rect 100 26726 2792 28198
tri 2792 27988 3002 28198 nw
rect 3438 27896 13317 27898
rect 3438 27840 3452 27896
rect 3508 27840 3532 27896
rect 3588 27840 3612 27896
rect 3668 27840 3693 27896
rect 3749 27840 3774 27896
rect 3830 27840 3855 27896
rect 3911 27840 3936 27896
rect 3992 27840 4017 27896
rect 4073 27840 4098 27896
rect 4154 27840 4179 27896
rect 4235 27840 4260 27896
rect 4316 27892 13317 27896
rect 4316 27883 5257 27892
rect 5309 27883 5323 27892
rect 5375 27883 6093 27892
rect 6145 27883 6159 27892
rect 6211 27883 6929 27892
rect 4316 27840 5215 27883
rect 5375 27840 5377 27883
rect 3438 27827 5215 27840
rect 5271 27827 5296 27840
rect 5352 27827 5377 27840
rect 5433 27827 5458 27883
rect 5514 27827 5539 27883
rect 5595 27827 5620 27883
rect 5676 27827 5701 27883
rect 5757 27827 5782 27883
rect 5838 27827 5863 27883
rect 5919 27827 5944 27883
rect 6000 27827 6025 27883
rect 6081 27840 6093 27883
rect 6081 27827 6106 27840
rect 6162 27827 6186 27840
rect 6242 27827 6266 27883
rect 6322 27827 6346 27883
rect 6402 27840 6929 27883
rect 6981 27840 6995 27892
rect 7047 27840 7765 27892
rect 7817 27840 7831 27892
rect 7883 27883 8601 27892
rect 8653 27883 8667 27892
rect 8719 27883 9437 27892
rect 9489 27883 9503 27892
rect 9555 27883 10273 27892
rect 7883 27840 8572 27883
rect 8719 27840 8732 27883
rect 6402 27827 8572 27840
rect 8628 27827 8652 27840
rect 8708 27827 8732 27840
rect 8788 27827 8812 27883
rect 8868 27827 8893 27883
rect 8949 27827 8974 27883
rect 9030 27827 9055 27883
rect 9111 27827 9136 27883
rect 9192 27827 9217 27883
rect 9273 27827 9298 27883
rect 9354 27827 9379 27883
rect 9435 27840 9437 27883
rect 9435 27827 9460 27840
rect 9516 27827 9541 27840
rect 9597 27827 9622 27883
rect 9678 27827 9703 27883
rect 9759 27840 10273 27883
rect 10325 27840 10339 27892
rect 10391 27883 11109 27892
rect 11161 27883 11175 27892
rect 11227 27883 11945 27892
rect 11997 27883 12011 27892
rect 10391 27840 10871 27883
rect 9759 27827 10871 27840
rect 10927 27827 10951 27883
rect 11007 27827 11031 27883
rect 11087 27840 11109 27883
rect 11167 27840 11175 27883
rect 11087 27827 11111 27840
rect 11167 27827 11192 27840
rect 11248 27827 11273 27883
rect 11329 27827 11354 27883
rect 11410 27827 11435 27883
rect 11491 27827 11516 27883
rect 11572 27827 11597 27883
rect 11653 27827 11678 27883
rect 11734 27827 11759 27883
rect 11815 27827 11840 27883
rect 11896 27827 11921 27883
rect 11997 27840 12002 27883
rect 12063 27840 12781 27892
rect 12833 27840 12847 27892
rect 12899 27840 13317 27892
rect 11977 27827 12002 27840
rect 12058 27827 13317 27840
rect 3438 27826 13317 27827
rect 3438 27802 5257 27826
rect 3438 27746 3452 27802
rect 3508 27746 3532 27802
rect 3588 27746 3612 27802
rect 3668 27746 3693 27802
rect 3749 27746 3774 27802
rect 3830 27746 3855 27802
rect 3911 27746 3936 27802
rect 3992 27746 4017 27802
rect 4073 27746 4098 27802
rect 4154 27746 4179 27802
rect 4235 27746 4260 27802
rect 4316 27795 5257 27802
rect 5309 27795 5323 27826
rect 5375 27795 6093 27826
rect 6145 27795 6159 27826
rect 6211 27795 6929 27826
rect 4316 27746 5215 27795
rect 5375 27774 5377 27795
rect 5271 27760 5296 27774
rect 5352 27760 5377 27774
rect 3438 27739 5215 27746
rect 5375 27739 5377 27760
rect 5433 27739 5458 27795
rect 5514 27739 5539 27795
rect 5595 27739 5620 27795
rect 5676 27739 5701 27795
rect 5757 27739 5782 27795
rect 5838 27739 5863 27795
rect 5919 27739 5944 27795
rect 6000 27739 6025 27795
rect 6081 27774 6093 27795
rect 6081 27760 6106 27774
rect 6162 27760 6186 27774
rect 6081 27739 6093 27760
rect 6242 27739 6266 27795
rect 6322 27739 6346 27795
rect 6402 27774 6929 27795
rect 6981 27774 6995 27826
rect 7047 27774 7765 27826
rect 7817 27774 7831 27826
rect 7883 27795 8601 27826
rect 8653 27795 8667 27826
rect 8719 27795 9437 27826
rect 9489 27795 9503 27826
rect 9555 27795 10273 27826
rect 7883 27774 8572 27795
rect 8719 27774 8732 27795
rect 6402 27760 8572 27774
rect 8628 27760 8652 27774
rect 8708 27760 8732 27774
rect 6402 27739 6929 27760
rect 3438 27708 5257 27739
rect 5309 27708 5323 27739
rect 5375 27708 6093 27739
rect 6145 27708 6159 27739
rect 6211 27708 6929 27739
rect 6981 27708 6995 27760
rect 7047 27708 7765 27760
rect 7817 27708 7831 27760
rect 7883 27739 8572 27760
rect 8719 27739 8732 27760
rect 8788 27739 8812 27795
rect 8868 27739 8893 27795
rect 8949 27739 8974 27795
rect 9030 27739 9055 27795
rect 9111 27739 9136 27795
rect 9192 27739 9217 27795
rect 9273 27739 9298 27795
rect 9354 27739 9379 27795
rect 9435 27774 9437 27795
rect 9435 27760 9460 27774
rect 9516 27760 9541 27774
rect 9435 27739 9437 27760
rect 9597 27739 9622 27795
rect 9678 27739 9703 27795
rect 9759 27774 10273 27795
rect 10325 27774 10339 27826
rect 10391 27795 11109 27826
rect 11161 27795 11175 27826
rect 11227 27795 11945 27826
rect 11997 27795 12011 27826
rect 10391 27774 10871 27795
rect 9759 27760 10871 27774
rect 9759 27739 10273 27760
rect 7883 27708 8601 27739
rect 8653 27708 8667 27739
rect 8719 27708 9437 27739
rect 9489 27708 9503 27739
rect 9555 27708 10273 27739
rect 10325 27708 10339 27760
rect 10391 27739 10871 27760
rect 10927 27739 10951 27795
rect 11007 27739 11031 27795
rect 11087 27774 11109 27795
rect 11167 27774 11175 27795
rect 11087 27760 11111 27774
rect 11167 27760 11192 27774
rect 11087 27739 11109 27760
rect 11167 27739 11175 27760
rect 11248 27739 11273 27795
rect 11329 27739 11354 27795
rect 11410 27739 11435 27795
rect 11491 27739 11516 27795
rect 11572 27739 11597 27795
rect 11653 27739 11678 27795
rect 11734 27739 11759 27795
rect 11815 27739 11840 27795
rect 11896 27739 11921 27795
rect 11997 27774 12002 27795
rect 12063 27774 12781 27826
rect 12833 27774 12847 27826
rect 12899 27774 13317 27826
rect 11977 27760 12002 27774
rect 12058 27760 13317 27774
rect 11997 27739 12002 27760
rect 10391 27708 11109 27739
rect 11161 27708 11175 27739
rect 11227 27708 11945 27739
rect 11997 27708 12011 27739
rect 12063 27708 12781 27760
rect 12833 27708 12847 27760
rect 12899 27708 13317 27760
rect 3438 27652 3452 27708
rect 3508 27652 3532 27708
rect 3588 27652 3612 27708
rect 3668 27652 3693 27708
rect 3749 27652 3774 27708
rect 3830 27652 3855 27708
rect 3911 27652 3936 27708
rect 3992 27652 4017 27708
rect 4073 27652 4098 27708
rect 4154 27652 4179 27708
rect 4235 27652 4260 27708
rect 4316 27707 13317 27708
rect 4316 27652 5215 27707
rect 5271 27694 5296 27707
rect 5352 27694 5377 27707
rect 3438 27651 5215 27652
rect 5375 27651 5377 27694
rect 5433 27651 5458 27707
rect 5514 27651 5539 27707
rect 5595 27651 5620 27707
rect 5676 27651 5701 27707
rect 5757 27651 5782 27707
rect 5838 27651 5863 27707
rect 5919 27651 5944 27707
rect 6000 27651 6025 27707
rect 6081 27694 6106 27707
rect 6162 27694 6186 27707
rect 6081 27651 6093 27694
rect 6242 27651 6266 27707
rect 6322 27651 6346 27707
rect 6402 27694 8572 27707
rect 8628 27694 8652 27707
rect 8708 27694 8732 27707
rect 6402 27651 6929 27694
rect 3438 27642 5257 27651
rect 5309 27642 5323 27651
rect 5375 27642 6093 27651
rect 6145 27642 6159 27651
rect 6211 27642 6929 27651
rect 6981 27642 6995 27694
rect 7047 27642 7765 27694
rect 7817 27642 7831 27694
rect 7883 27651 8572 27694
rect 8719 27651 8732 27694
rect 8788 27651 8812 27707
rect 8868 27651 8893 27707
rect 8949 27651 8974 27707
rect 9030 27651 9055 27707
rect 9111 27651 9136 27707
rect 9192 27651 9217 27707
rect 9273 27651 9298 27707
rect 9354 27651 9379 27707
rect 9435 27694 9460 27707
rect 9516 27694 9541 27707
rect 9435 27651 9437 27694
rect 9597 27651 9622 27707
rect 9678 27651 9703 27707
rect 9759 27694 10871 27707
rect 9759 27651 10273 27694
rect 7883 27642 8601 27651
rect 8653 27642 8667 27651
rect 8719 27642 9437 27651
rect 9489 27642 9503 27651
rect 9555 27642 10273 27651
rect 10325 27642 10339 27694
rect 10391 27651 10871 27694
rect 10927 27651 10951 27707
rect 11007 27651 11031 27707
rect 11087 27694 11111 27707
rect 11167 27694 11192 27707
rect 11087 27651 11109 27694
rect 11167 27651 11175 27694
rect 11248 27651 11273 27707
rect 11329 27651 11354 27707
rect 11410 27651 11435 27707
rect 11491 27651 11516 27707
rect 11572 27651 11597 27707
rect 11653 27651 11678 27707
rect 11734 27651 11759 27707
rect 11815 27651 11840 27707
rect 11896 27651 11921 27707
rect 11977 27694 12002 27707
rect 12058 27694 13317 27707
rect 11997 27651 12002 27694
rect 10391 27642 11109 27651
rect 11161 27642 11175 27651
rect 11227 27642 11945 27651
rect 11997 27642 12011 27651
rect 12063 27642 12781 27694
rect 12833 27642 12847 27694
rect 12899 27642 13317 27694
rect 3438 27627 13317 27642
rect 3438 27619 5257 27627
rect 5309 27619 5323 27627
rect 5375 27619 6093 27627
rect 6145 27619 6159 27627
rect 6211 27619 6929 27627
rect 3438 27614 5215 27619
rect 3438 27558 3452 27614
rect 3508 27558 3532 27614
rect 3588 27558 3612 27614
rect 3668 27558 3693 27614
rect 3749 27558 3774 27614
rect 3830 27558 3855 27614
rect 3911 27558 3936 27614
rect 3992 27558 4017 27614
rect 4073 27558 4098 27614
rect 4154 27558 4179 27614
rect 4235 27558 4260 27614
rect 4316 27563 5215 27614
rect 5375 27575 5377 27619
rect 5271 27563 5296 27575
rect 5352 27563 5377 27575
rect 5433 27563 5458 27619
rect 5514 27563 5539 27619
rect 5595 27563 5620 27619
rect 5676 27563 5701 27619
rect 5757 27563 5782 27619
rect 5838 27563 5863 27619
rect 5919 27563 5944 27619
rect 6000 27563 6025 27619
rect 6081 27575 6093 27619
rect 6081 27563 6106 27575
rect 6162 27563 6186 27575
rect 6242 27563 6266 27619
rect 6322 27563 6346 27619
rect 6402 27575 6929 27619
rect 6981 27575 6995 27627
rect 7047 27575 7765 27627
rect 7817 27575 7831 27627
rect 7883 27619 8601 27627
rect 8653 27619 8667 27627
rect 8719 27619 9437 27627
rect 9489 27619 9503 27627
rect 9555 27619 10273 27627
rect 7883 27575 8572 27619
rect 8719 27575 8732 27619
rect 6402 27563 8572 27575
rect 8628 27563 8652 27575
rect 8708 27563 8732 27575
rect 8788 27563 8812 27619
rect 8868 27563 8893 27619
rect 8949 27563 8974 27619
rect 9030 27563 9055 27619
rect 9111 27563 9136 27619
rect 9192 27563 9217 27619
rect 9273 27563 9298 27619
rect 9354 27563 9379 27619
rect 9435 27575 9437 27619
rect 9435 27563 9460 27575
rect 9516 27563 9541 27575
rect 9597 27563 9622 27619
rect 9678 27563 9703 27619
rect 9759 27575 10273 27619
rect 10325 27575 10339 27627
rect 10391 27619 11109 27627
rect 11161 27619 11175 27627
rect 11227 27619 11945 27627
rect 11997 27619 12011 27627
rect 10391 27575 10871 27619
rect 9759 27563 10871 27575
rect 10927 27563 10951 27619
rect 11007 27563 11031 27619
rect 11087 27575 11109 27619
rect 11167 27575 11175 27619
rect 11087 27563 11111 27575
rect 11167 27563 11192 27575
rect 11248 27563 11273 27619
rect 11329 27563 11354 27619
rect 11410 27563 11435 27619
rect 11491 27563 11516 27619
rect 11572 27563 11597 27619
rect 11653 27563 11678 27619
rect 11734 27563 11759 27619
rect 11815 27563 11840 27619
rect 11896 27563 11921 27619
rect 11997 27575 12002 27619
rect 12063 27575 12781 27627
rect 12833 27575 12847 27627
rect 12899 27575 13317 27627
rect 11977 27563 12002 27575
rect 12058 27563 13317 27575
rect 4316 27560 13317 27563
rect 4316 27558 5257 27560
rect 3438 27531 5257 27558
rect 5309 27531 5323 27560
rect 5375 27531 6093 27560
rect 6145 27531 6159 27560
rect 6211 27531 6929 27560
rect 3438 27520 5215 27531
rect 3438 27464 3452 27520
rect 3508 27464 3532 27520
rect 3588 27464 3612 27520
rect 3668 27464 3693 27520
rect 3749 27464 3774 27520
rect 3830 27464 3855 27520
rect 3911 27464 3936 27520
rect 3992 27464 4017 27520
rect 4073 27464 4098 27520
rect 4154 27464 4179 27520
rect 4235 27464 4260 27520
rect 4316 27475 5215 27520
rect 5375 27508 5377 27531
rect 5271 27493 5296 27508
rect 5352 27493 5377 27508
rect 5375 27475 5377 27493
rect 5433 27475 5458 27531
rect 5514 27475 5539 27531
rect 5595 27475 5620 27531
rect 5676 27475 5701 27531
rect 5757 27475 5782 27531
rect 5838 27475 5863 27531
rect 5919 27475 5944 27531
rect 6000 27475 6025 27531
rect 6081 27508 6093 27531
rect 6081 27493 6106 27508
rect 6162 27493 6186 27508
rect 6081 27475 6093 27493
rect 6242 27475 6266 27531
rect 6322 27475 6346 27531
rect 6402 27508 6929 27531
rect 6981 27508 6995 27560
rect 7047 27508 7765 27560
rect 7817 27508 7831 27560
rect 7883 27531 8601 27560
rect 8653 27531 8667 27560
rect 8719 27531 9437 27560
rect 9489 27531 9503 27560
rect 9555 27531 10273 27560
rect 7883 27508 8572 27531
rect 8719 27508 8732 27531
rect 6402 27493 8572 27508
rect 8628 27493 8652 27508
rect 8708 27493 8732 27508
rect 6402 27475 6929 27493
rect 4316 27464 5257 27475
rect 3438 27443 5257 27464
rect 5309 27443 5323 27475
rect 5375 27443 6093 27475
rect 6145 27443 6159 27475
rect 6211 27443 6929 27475
rect 3438 27426 5215 27443
rect 5375 27441 5377 27443
rect 5271 27426 5296 27441
rect 5352 27426 5377 27441
rect 3438 27370 3452 27426
rect 3508 27370 3532 27426
rect 3588 27370 3612 27426
rect 3668 27370 3693 27426
rect 3749 27370 3774 27426
rect 3830 27370 3855 27426
rect 3911 27370 3936 27426
rect 3992 27370 4017 27426
rect 4073 27370 4098 27426
rect 4154 27370 4179 27426
rect 4235 27370 4260 27426
rect 4316 27387 5215 27426
rect 5375 27387 5377 27426
rect 5433 27387 5458 27443
rect 5514 27387 5539 27443
rect 5595 27387 5620 27443
rect 5676 27387 5701 27443
rect 5757 27387 5782 27443
rect 5838 27387 5863 27443
rect 5919 27387 5944 27443
rect 6000 27387 6025 27443
rect 6081 27441 6093 27443
rect 6081 27426 6106 27441
rect 6162 27426 6186 27441
rect 6081 27387 6093 27426
rect 6242 27387 6266 27443
rect 6322 27387 6346 27443
rect 6402 27441 6929 27443
rect 6981 27441 6995 27493
rect 7047 27441 7765 27493
rect 7817 27441 7831 27493
rect 7883 27475 8572 27493
rect 8719 27475 8732 27493
rect 8788 27475 8812 27531
rect 8868 27475 8893 27531
rect 8949 27475 8974 27531
rect 9030 27475 9055 27531
rect 9111 27475 9136 27531
rect 9192 27475 9217 27531
rect 9273 27475 9298 27531
rect 9354 27475 9379 27531
rect 9435 27508 9437 27531
rect 9435 27493 9460 27508
rect 9516 27493 9541 27508
rect 9435 27475 9437 27493
rect 9597 27475 9622 27531
rect 9678 27475 9703 27531
rect 9759 27508 10273 27531
rect 10325 27508 10339 27560
rect 10391 27531 11109 27560
rect 11161 27531 11175 27560
rect 11227 27531 11945 27560
rect 11997 27531 12011 27560
rect 10391 27508 10871 27531
rect 9759 27493 10871 27508
rect 9759 27475 10273 27493
rect 7883 27443 8601 27475
rect 8653 27443 8667 27475
rect 8719 27443 9437 27475
rect 9489 27443 9503 27475
rect 9555 27443 10273 27475
rect 7883 27441 8572 27443
rect 8719 27441 8732 27443
rect 6402 27426 8572 27441
rect 8628 27426 8652 27441
rect 8708 27426 8732 27441
rect 6402 27387 6929 27426
rect 4316 27374 5257 27387
rect 5309 27374 5323 27387
rect 5375 27374 6093 27387
rect 6145 27374 6159 27387
rect 6211 27374 6929 27387
rect 6981 27374 6995 27426
rect 7047 27374 7765 27426
rect 7817 27374 7831 27426
rect 7883 27387 8572 27426
rect 8719 27387 8732 27426
rect 8788 27387 8812 27443
rect 8868 27387 8893 27443
rect 8949 27387 8974 27443
rect 9030 27387 9055 27443
rect 9111 27387 9136 27443
rect 9192 27387 9217 27443
rect 9273 27387 9298 27443
rect 9354 27387 9379 27443
rect 9435 27441 9437 27443
rect 9435 27426 9460 27441
rect 9516 27426 9541 27441
rect 9435 27387 9437 27426
rect 9597 27387 9622 27443
rect 9678 27387 9703 27443
rect 9759 27441 10273 27443
rect 10325 27441 10339 27493
rect 10391 27475 10871 27493
rect 10927 27475 10951 27531
rect 11007 27475 11031 27531
rect 11087 27508 11109 27531
rect 11167 27508 11175 27531
rect 11087 27493 11111 27508
rect 11167 27493 11192 27508
rect 11087 27475 11109 27493
rect 11167 27475 11175 27493
rect 11248 27475 11273 27531
rect 11329 27475 11354 27531
rect 11410 27475 11435 27531
rect 11491 27475 11516 27531
rect 11572 27475 11597 27531
rect 11653 27475 11678 27531
rect 11734 27475 11759 27531
rect 11815 27475 11840 27531
rect 11896 27475 11921 27531
rect 11997 27508 12002 27531
rect 12063 27508 12781 27560
rect 12833 27508 12847 27560
rect 12899 27508 13317 27560
rect 11977 27493 12002 27508
rect 12058 27493 13317 27508
rect 11997 27475 12002 27493
rect 10391 27443 11109 27475
rect 11161 27443 11175 27475
rect 11227 27443 11945 27475
rect 11997 27443 12011 27475
rect 10391 27441 10871 27443
rect 9759 27426 10871 27441
rect 9759 27387 10273 27426
rect 7883 27374 8601 27387
rect 8653 27374 8667 27387
rect 8719 27374 9437 27387
rect 9489 27374 9503 27387
rect 9555 27374 10273 27387
rect 10325 27374 10339 27426
rect 10391 27387 10871 27426
rect 10927 27387 10951 27443
rect 11007 27387 11031 27443
rect 11087 27441 11109 27443
rect 11167 27441 11175 27443
rect 11087 27426 11111 27441
rect 11167 27426 11192 27441
rect 11087 27387 11109 27426
rect 11167 27387 11175 27426
rect 11248 27387 11273 27443
rect 11329 27387 11354 27443
rect 11410 27387 11435 27443
rect 11491 27387 11516 27443
rect 11572 27387 11597 27443
rect 11653 27387 11678 27443
rect 11734 27387 11759 27443
rect 11815 27387 11840 27443
rect 11896 27387 11921 27443
rect 11997 27441 12002 27443
rect 12063 27441 12781 27493
rect 12833 27441 12847 27493
rect 12899 27441 13317 27493
rect 11977 27426 12002 27441
rect 12058 27426 13317 27441
rect 11997 27387 12002 27426
rect 10391 27374 11109 27387
rect 11161 27374 11175 27387
rect 11227 27374 11945 27387
rect 11997 27374 12011 27387
rect 12063 27374 12781 27426
rect 12833 27374 12847 27426
rect 12899 27374 13317 27426
rect 4316 27370 13317 27374
rect 3438 27368 13317 27370
tri 2792 26726 3002 26936 sw
rect 100 26720 13602 26726
rect 100 26668 4839 26720
rect 4891 26668 4905 26720
rect 4957 26668 5675 26720
rect 5727 26668 5741 26720
rect 5793 26668 6511 26720
rect 6563 26668 6577 26720
rect 6629 26668 7347 26720
rect 7399 26668 7413 26720
rect 7465 26668 8183 26720
rect 8235 26668 8249 26720
rect 8301 26668 9019 26720
rect 9071 26668 9085 26720
rect 9137 26668 9855 26720
rect 9907 26668 9921 26720
rect 9973 26668 10691 26720
rect 10743 26668 10757 26720
rect 10809 26668 11527 26720
rect 11579 26668 11593 26720
rect 11645 26668 12363 26720
rect 12415 26668 12429 26720
rect 12481 26668 13200 26720
rect 13252 26668 13270 26720
rect 13322 26668 13340 26720
rect 13392 26668 13410 26720
rect 13462 26668 13480 26720
rect 13532 26668 13550 26720
rect 100 26654 13602 26668
rect 100 26602 4839 26654
rect 4891 26602 4905 26654
rect 4957 26602 5675 26654
rect 5727 26602 5741 26654
rect 5793 26602 6511 26654
rect 6563 26602 6577 26654
rect 6629 26602 7347 26654
rect 7399 26602 7413 26654
rect 7465 26602 8183 26654
rect 8235 26602 8249 26654
rect 8301 26602 9019 26654
rect 9071 26602 9085 26654
rect 9137 26602 9855 26654
rect 9907 26602 9921 26654
rect 9973 26602 10691 26654
rect 10743 26602 10757 26654
rect 10809 26602 11527 26654
rect 11579 26602 11593 26654
rect 11645 26602 12363 26654
rect 12415 26602 12429 26654
rect 12481 26602 13200 26654
rect 13252 26602 13270 26654
rect 13322 26602 13340 26654
rect 13392 26602 13410 26654
rect 13462 26602 13480 26654
rect 13532 26602 13550 26654
rect 100 26588 13602 26602
rect 100 26536 4839 26588
rect 4891 26536 4905 26588
rect 4957 26536 5675 26588
rect 5727 26536 5741 26588
rect 5793 26536 6511 26588
rect 6563 26536 6577 26588
rect 6629 26536 7347 26588
rect 7399 26536 7413 26588
rect 7465 26536 8183 26588
rect 8235 26536 8249 26588
rect 8301 26536 9019 26588
rect 9071 26536 9085 26588
rect 9137 26536 9855 26588
rect 9907 26536 9921 26588
rect 9973 26536 10691 26588
rect 10743 26536 10757 26588
rect 10809 26536 11527 26588
rect 11579 26536 11593 26588
rect 11645 26536 12363 26588
rect 12415 26536 12429 26588
rect 12481 26536 13200 26588
rect 13252 26536 13270 26588
rect 13322 26536 13340 26588
rect 13392 26536 13410 26588
rect 13462 26536 13480 26588
rect 13532 26536 13550 26588
rect 100 26522 13602 26536
rect 100 26470 4839 26522
rect 4891 26470 4905 26522
rect 4957 26470 5675 26522
rect 5727 26470 5741 26522
rect 5793 26470 6511 26522
rect 6563 26470 6577 26522
rect 6629 26470 7347 26522
rect 7399 26470 7413 26522
rect 7465 26470 8183 26522
rect 8235 26470 8249 26522
rect 8301 26470 9019 26522
rect 9071 26470 9085 26522
rect 9137 26470 9855 26522
rect 9907 26470 9921 26522
rect 9973 26470 10691 26522
rect 10743 26470 10757 26522
rect 10809 26470 11527 26522
rect 11579 26470 11593 26522
rect 11645 26470 12363 26522
rect 12415 26470 12429 26522
rect 12481 26470 13200 26522
rect 13252 26470 13270 26522
rect 13322 26470 13340 26522
rect 13392 26470 13410 26522
rect 13462 26470 13480 26522
rect 13532 26470 13550 26522
rect 100 26456 13602 26470
rect 100 26404 4839 26456
rect 4891 26404 4905 26456
rect 4957 26404 5675 26456
rect 5727 26404 5741 26456
rect 5793 26404 6511 26456
rect 6563 26404 6577 26456
rect 6629 26404 7347 26456
rect 7399 26404 7413 26456
rect 7465 26404 8183 26456
rect 8235 26404 8249 26456
rect 8301 26404 9019 26456
rect 9071 26404 9085 26456
rect 9137 26404 9855 26456
rect 9907 26404 9921 26456
rect 9973 26404 10691 26456
rect 10743 26404 10757 26456
rect 10809 26404 11527 26456
rect 11579 26404 11593 26456
rect 11645 26404 12363 26456
rect 12415 26404 12429 26456
rect 12481 26404 13200 26456
rect 13252 26404 13270 26456
rect 13322 26404 13340 26456
rect 13392 26404 13410 26456
rect 13462 26404 13480 26456
rect 13532 26404 13550 26456
rect 100 26389 13602 26404
rect 100 26337 4839 26389
rect 4891 26337 4905 26389
rect 4957 26337 5675 26389
rect 5727 26337 5741 26389
rect 5793 26337 6511 26389
rect 6563 26337 6577 26389
rect 6629 26337 7347 26389
rect 7399 26337 7413 26389
rect 7465 26337 8183 26389
rect 8235 26337 8249 26389
rect 8301 26337 9019 26389
rect 9071 26337 9085 26389
rect 9137 26337 9855 26389
rect 9907 26337 9921 26389
rect 9973 26337 10691 26389
rect 10743 26337 10757 26389
rect 10809 26337 11527 26389
rect 11579 26337 11593 26389
rect 11645 26337 12363 26389
rect 12415 26337 12429 26389
rect 12481 26337 13200 26389
rect 13252 26337 13270 26389
rect 13322 26337 13340 26389
rect 13392 26337 13410 26389
rect 13462 26337 13480 26389
rect 13532 26337 13550 26389
rect 100 26322 13602 26337
rect 100 26270 4839 26322
rect 4891 26270 4905 26322
rect 4957 26270 5675 26322
rect 5727 26270 5741 26322
rect 5793 26270 6511 26322
rect 6563 26270 6577 26322
rect 6629 26270 7347 26322
rect 7399 26270 7413 26322
rect 7465 26270 8183 26322
rect 8235 26270 8249 26322
rect 8301 26270 9019 26322
rect 9071 26270 9085 26322
rect 9137 26270 9855 26322
rect 9907 26270 9921 26322
rect 9973 26270 10691 26322
rect 10743 26270 10757 26322
rect 10809 26270 11527 26322
rect 11579 26270 11593 26322
rect 11645 26270 12363 26322
rect 12415 26270 12429 26322
rect 12481 26270 13200 26322
rect 13252 26270 13270 26322
rect 13322 26270 13340 26322
rect 13392 26270 13410 26322
rect 13462 26270 13480 26322
rect 13532 26270 13550 26322
rect 100 26255 13602 26270
rect 100 26203 4839 26255
rect 4891 26203 4905 26255
rect 4957 26203 5675 26255
rect 5727 26203 5741 26255
rect 5793 26203 6511 26255
rect 6563 26203 6577 26255
rect 6629 26203 7347 26255
rect 7399 26203 7413 26255
rect 7465 26203 8183 26255
rect 8235 26203 8249 26255
rect 8301 26203 9019 26255
rect 9071 26203 9085 26255
rect 9137 26203 9855 26255
rect 9907 26203 9921 26255
rect 9973 26203 10691 26255
rect 10743 26203 10757 26255
rect 10809 26203 11527 26255
rect 11579 26203 11593 26255
rect 11645 26203 12363 26255
rect 12415 26203 12429 26255
rect 12481 26203 13200 26255
rect 13252 26203 13270 26255
rect 13322 26203 13340 26255
rect 13392 26203 13410 26255
rect 13462 26203 13480 26255
rect 13532 26203 13550 26255
rect 100 26197 13602 26203
rect 100 14901 2792 26197
tri 2792 25987 3002 26197 nw
rect 3434 25891 13317 25897
rect 3434 25882 5257 25891
rect 5309 25882 5323 25891
rect 5375 25882 6093 25891
rect 6145 25882 6159 25891
rect 6211 25882 6929 25891
rect 3434 25826 3443 25882
rect 3499 25826 3525 25882
rect 3581 25826 3607 25882
rect 3663 25826 3689 25882
rect 3745 25826 3771 25882
rect 3827 25826 3853 25882
rect 3909 25826 3935 25882
rect 3991 25826 4017 25882
rect 4073 25826 4098 25882
rect 4154 25826 4179 25882
rect 4235 25826 4260 25882
rect 4316 25826 5215 25882
rect 5375 25839 5377 25882
rect 5271 25826 5296 25839
rect 5352 25826 5377 25839
rect 5433 25826 5458 25882
rect 5514 25826 5539 25882
rect 5595 25826 5620 25882
rect 5676 25826 5701 25882
rect 5757 25826 5782 25882
rect 5838 25826 5863 25882
rect 5919 25826 5944 25882
rect 6000 25826 6025 25882
rect 6081 25839 6093 25882
rect 6081 25826 6106 25839
rect 6162 25826 6186 25839
rect 6242 25826 6266 25882
rect 6322 25826 6346 25882
rect 6402 25839 6929 25882
rect 6981 25839 6995 25891
rect 7047 25839 7765 25891
rect 7817 25839 7831 25891
rect 7883 25882 8601 25891
rect 8653 25882 8667 25891
rect 8719 25882 9437 25891
rect 9489 25882 9503 25891
rect 9555 25882 10273 25891
rect 7883 25839 8572 25882
rect 8719 25839 8732 25882
rect 6402 25826 8572 25839
rect 8628 25826 8652 25839
rect 8708 25826 8732 25839
rect 8788 25826 8812 25882
rect 8868 25826 8893 25882
rect 8949 25826 8974 25882
rect 9030 25826 9055 25882
rect 9111 25826 9136 25882
rect 9192 25826 9217 25882
rect 9273 25826 9298 25882
rect 9354 25826 9379 25882
rect 9435 25839 9437 25882
rect 9435 25826 9460 25839
rect 9516 25826 9541 25839
rect 9597 25826 9622 25882
rect 9678 25826 9703 25882
rect 9759 25839 10273 25882
rect 10325 25839 10339 25891
rect 10391 25882 11109 25891
rect 11161 25882 11175 25891
rect 11227 25882 11945 25891
rect 11997 25882 12011 25891
rect 10391 25839 10871 25882
rect 9759 25826 10871 25839
rect 10927 25826 10951 25882
rect 11007 25826 11031 25882
rect 11087 25839 11109 25882
rect 11167 25839 11175 25882
rect 11087 25826 11111 25839
rect 11167 25826 11192 25839
rect 11248 25826 11273 25882
rect 11329 25826 11354 25882
rect 11410 25826 11435 25882
rect 11491 25826 11516 25882
rect 11572 25826 11597 25882
rect 11653 25826 11678 25882
rect 11734 25826 11759 25882
rect 11815 25826 11840 25882
rect 11896 25826 11921 25882
rect 11997 25839 12002 25882
rect 12063 25839 12781 25891
rect 12833 25839 12847 25891
rect 12899 25839 13317 25891
rect 11977 25826 12002 25839
rect 12058 25826 13317 25839
rect 3434 25825 13317 25826
rect 3434 25794 5257 25825
rect 5309 25794 5323 25825
rect 5375 25794 6093 25825
rect 6145 25794 6159 25825
rect 6211 25794 6929 25825
rect 3434 25738 3443 25794
rect 3499 25738 3525 25794
rect 3581 25738 3607 25794
rect 3663 25738 3689 25794
rect 3745 25738 3771 25794
rect 3827 25738 3853 25794
rect 3909 25738 3935 25794
rect 3991 25738 4017 25794
rect 4073 25738 4098 25794
rect 4154 25738 4179 25794
rect 4235 25738 4260 25794
rect 4316 25738 5215 25794
rect 5375 25773 5377 25794
rect 5271 25759 5296 25773
rect 5352 25759 5377 25773
rect 5375 25738 5377 25759
rect 5433 25738 5458 25794
rect 5514 25738 5539 25794
rect 5595 25738 5620 25794
rect 5676 25738 5701 25794
rect 5757 25738 5782 25794
rect 5838 25738 5863 25794
rect 5919 25738 5944 25794
rect 6000 25738 6025 25794
rect 6081 25773 6093 25794
rect 6081 25759 6106 25773
rect 6162 25759 6186 25773
rect 6081 25738 6093 25759
rect 6242 25738 6266 25794
rect 6322 25738 6346 25794
rect 6402 25773 6929 25794
rect 6981 25773 6995 25825
rect 7047 25773 7765 25825
rect 7817 25773 7831 25825
rect 7883 25794 8601 25825
rect 8653 25794 8667 25825
rect 8719 25794 9437 25825
rect 9489 25794 9503 25825
rect 9555 25794 10273 25825
rect 7883 25773 8572 25794
rect 8719 25773 8732 25794
rect 6402 25759 8572 25773
rect 8628 25759 8652 25773
rect 8708 25759 8732 25773
rect 6402 25738 6929 25759
rect 3434 25707 5257 25738
rect 5309 25707 5323 25738
rect 5375 25707 6093 25738
rect 6145 25707 6159 25738
rect 6211 25707 6929 25738
rect 6981 25707 6995 25759
rect 7047 25707 7765 25759
rect 7817 25707 7831 25759
rect 7883 25738 8572 25759
rect 8719 25738 8732 25759
rect 8788 25738 8812 25794
rect 8868 25738 8893 25794
rect 8949 25738 8974 25794
rect 9030 25738 9055 25794
rect 9111 25738 9136 25794
rect 9192 25738 9217 25794
rect 9273 25738 9298 25794
rect 9354 25738 9379 25794
rect 9435 25773 9437 25794
rect 9435 25759 9460 25773
rect 9516 25759 9541 25773
rect 9435 25738 9437 25759
rect 9597 25738 9622 25794
rect 9678 25738 9703 25794
rect 9759 25773 10273 25794
rect 10325 25773 10339 25825
rect 10391 25794 11109 25825
rect 11161 25794 11175 25825
rect 11227 25794 11945 25825
rect 11997 25794 12011 25825
rect 10391 25773 10871 25794
rect 9759 25759 10871 25773
rect 9759 25738 10273 25759
rect 7883 25707 8601 25738
rect 8653 25707 8667 25738
rect 8719 25707 9437 25738
rect 9489 25707 9503 25738
rect 9555 25707 10273 25738
rect 10325 25707 10339 25759
rect 10391 25738 10871 25759
rect 10927 25738 10951 25794
rect 11007 25738 11031 25794
rect 11087 25773 11109 25794
rect 11167 25773 11175 25794
rect 11087 25759 11111 25773
rect 11167 25759 11192 25773
rect 11087 25738 11109 25759
rect 11167 25738 11175 25759
rect 11248 25738 11273 25794
rect 11329 25738 11354 25794
rect 11410 25738 11435 25794
rect 11491 25738 11516 25794
rect 11572 25738 11597 25794
rect 11653 25738 11678 25794
rect 11734 25738 11759 25794
rect 11815 25738 11840 25794
rect 11896 25738 11921 25794
rect 11997 25773 12002 25794
rect 12063 25773 12781 25825
rect 12833 25773 12847 25825
rect 12899 25773 13317 25825
rect 11977 25759 12002 25773
rect 12058 25759 13317 25773
rect 11997 25738 12002 25759
rect 10391 25707 11109 25738
rect 11161 25707 11175 25738
rect 11227 25707 11945 25738
rect 11997 25707 12011 25738
rect 12063 25707 12781 25759
rect 12833 25707 12847 25759
rect 12899 25707 13317 25759
rect 3434 25706 13317 25707
rect 3434 25650 3443 25706
rect 3499 25650 3525 25706
rect 3581 25650 3607 25706
rect 3663 25650 3689 25706
rect 3745 25650 3771 25706
rect 3827 25650 3853 25706
rect 3909 25650 3935 25706
rect 3991 25650 4017 25706
rect 4073 25650 4098 25706
rect 4154 25650 4179 25706
rect 4235 25650 4260 25706
rect 4316 25650 5215 25706
rect 5271 25693 5296 25706
rect 5352 25693 5377 25706
rect 5375 25650 5377 25693
rect 5433 25650 5458 25706
rect 5514 25650 5539 25706
rect 5595 25650 5620 25706
rect 5676 25650 5701 25706
rect 5757 25650 5782 25706
rect 5838 25650 5863 25706
rect 5919 25650 5944 25706
rect 6000 25650 6025 25706
rect 6081 25693 6106 25706
rect 6162 25693 6186 25706
rect 6081 25650 6093 25693
rect 6242 25650 6266 25706
rect 6322 25650 6346 25706
rect 6402 25693 8572 25706
rect 8628 25693 8652 25706
rect 8708 25693 8732 25706
rect 6402 25650 6929 25693
rect 3434 25641 5257 25650
rect 5309 25641 5323 25650
rect 5375 25641 6093 25650
rect 6145 25641 6159 25650
rect 6211 25641 6929 25650
rect 6981 25641 6995 25693
rect 7047 25641 7765 25693
rect 7817 25641 7831 25693
rect 7883 25650 8572 25693
rect 8719 25650 8732 25693
rect 8788 25650 8812 25706
rect 8868 25650 8893 25706
rect 8949 25650 8974 25706
rect 9030 25650 9055 25706
rect 9111 25650 9136 25706
rect 9192 25650 9217 25706
rect 9273 25650 9298 25706
rect 9354 25650 9379 25706
rect 9435 25693 9460 25706
rect 9516 25693 9541 25706
rect 9435 25650 9437 25693
rect 9597 25650 9622 25706
rect 9678 25650 9703 25706
rect 9759 25693 10871 25706
rect 9759 25650 10273 25693
rect 7883 25641 8601 25650
rect 8653 25641 8667 25650
rect 8719 25641 9437 25650
rect 9489 25641 9503 25650
rect 9555 25641 10273 25650
rect 10325 25641 10339 25693
rect 10391 25650 10871 25693
rect 10927 25650 10951 25706
rect 11007 25650 11031 25706
rect 11087 25693 11111 25706
rect 11167 25693 11192 25706
rect 11087 25650 11109 25693
rect 11167 25650 11175 25693
rect 11248 25650 11273 25706
rect 11329 25650 11354 25706
rect 11410 25650 11435 25706
rect 11491 25650 11516 25706
rect 11572 25650 11597 25706
rect 11653 25650 11678 25706
rect 11734 25650 11759 25706
rect 11815 25650 11840 25706
rect 11896 25650 11921 25706
rect 11977 25693 12002 25706
rect 12058 25693 13317 25706
rect 11997 25650 12002 25693
rect 10391 25641 11109 25650
rect 11161 25641 11175 25650
rect 11227 25641 11945 25650
rect 11997 25641 12011 25650
rect 12063 25641 12781 25693
rect 12833 25641 12847 25693
rect 12899 25641 13317 25693
rect 3434 25626 13317 25641
rect 3434 25618 5257 25626
rect 5309 25618 5323 25626
rect 5375 25618 6093 25626
rect 6145 25618 6159 25626
rect 6211 25618 6929 25626
rect 3434 25562 3443 25618
rect 3499 25562 3525 25618
rect 3581 25562 3607 25618
rect 3663 25562 3689 25618
rect 3745 25562 3771 25618
rect 3827 25562 3853 25618
rect 3909 25562 3935 25618
rect 3991 25562 4017 25618
rect 4073 25562 4098 25618
rect 4154 25562 4179 25618
rect 4235 25562 4260 25618
rect 4316 25562 5215 25618
rect 5375 25574 5377 25618
rect 5271 25562 5296 25574
rect 5352 25562 5377 25574
rect 5433 25562 5458 25618
rect 5514 25562 5539 25618
rect 5595 25562 5620 25618
rect 5676 25562 5701 25618
rect 5757 25562 5782 25618
rect 5838 25562 5863 25618
rect 5919 25562 5944 25618
rect 6000 25562 6025 25618
rect 6081 25574 6093 25618
rect 6081 25562 6106 25574
rect 6162 25562 6186 25574
rect 6242 25562 6266 25618
rect 6322 25562 6346 25618
rect 6402 25574 6929 25618
rect 6981 25574 6995 25626
rect 7047 25574 7765 25626
rect 7817 25574 7831 25626
rect 7883 25618 8601 25626
rect 8653 25618 8667 25626
rect 8719 25618 9437 25626
rect 9489 25618 9503 25626
rect 9555 25618 10273 25626
rect 7883 25574 8572 25618
rect 8719 25574 8732 25618
rect 6402 25562 8572 25574
rect 8628 25562 8652 25574
rect 8708 25562 8732 25574
rect 8788 25562 8812 25618
rect 8868 25562 8893 25618
rect 8949 25562 8974 25618
rect 9030 25562 9055 25618
rect 9111 25562 9136 25618
rect 9192 25562 9217 25618
rect 9273 25562 9298 25618
rect 9354 25562 9379 25618
rect 9435 25574 9437 25618
rect 9435 25562 9460 25574
rect 9516 25562 9541 25574
rect 9597 25562 9622 25618
rect 9678 25562 9703 25618
rect 9759 25574 10273 25618
rect 10325 25574 10339 25626
rect 10391 25618 11109 25626
rect 11161 25618 11175 25626
rect 11227 25618 11945 25626
rect 11997 25618 12011 25626
rect 10391 25574 10871 25618
rect 9759 25562 10871 25574
rect 10927 25562 10951 25618
rect 11007 25562 11031 25618
rect 11087 25574 11109 25618
rect 11167 25574 11175 25618
rect 11087 25562 11111 25574
rect 11167 25562 11192 25574
rect 11248 25562 11273 25618
rect 11329 25562 11354 25618
rect 11410 25562 11435 25618
rect 11491 25562 11516 25618
rect 11572 25562 11597 25618
rect 11653 25562 11678 25618
rect 11734 25562 11759 25618
rect 11815 25562 11840 25618
rect 11896 25562 11921 25618
rect 11997 25574 12002 25618
rect 12063 25574 12781 25626
rect 12833 25574 12847 25626
rect 12899 25574 13317 25626
rect 11977 25562 12002 25574
rect 12058 25562 13317 25574
rect 3434 25559 13317 25562
rect 3434 25530 5257 25559
rect 5309 25530 5323 25559
rect 5375 25530 6093 25559
rect 6145 25530 6159 25559
rect 6211 25530 6929 25559
rect 3434 25474 3443 25530
rect 3499 25474 3525 25530
rect 3581 25474 3607 25530
rect 3663 25474 3689 25530
rect 3745 25474 3771 25530
rect 3827 25474 3853 25530
rect 3909 25474 3935 25530
rect 3991 25474 4017 25530
rect 4073 25474 4098 25530
rect 4154 25474 4179 25530
rect 4235 25474 4260 25530
rect 4316 25474 5215 25530
rect 5375 25507 5377 25530
rect 5271 25492 5296 25507
rect 5352 25492 5377 25507
rect 5375 25474 5377 25492
rect 5433 25474 5458 25530
rect 5514 25474 5539 25530
rect 5595 25474 5620 25530
rect 5676 25474 5701 25530
rect 5757 25474 5782 25530
rect 5838 25474 5863 25530
rect 5919 25474 5944 25530
rect 6000 25474 6025 25530
rect 6081 25507 6093 25530
rect 6081 25492 6106 25507
rect 6162 25492 6186 25507
rect 6081 25474 6093 25492
rect 6242 25474 6266 25530
rect 6322 25474 6346 25530
rect 6402 25507 6929 25530
rect 6981 25507 6995 25559
rect 7047 25507 7765 25559
rect 7817 25507 7831 25559
rect 7883 25530 8601 25559
rect 8653 25530 8667 25559
rect 8719 25530 9437 25559
rect 9489 25530 9503 25559
rect 9555 25530 10273 25559
rect 7883 25507 8572 25530
rect 8719 25507 8732 25530
rect 6402 25492 8572 25507
rect 8628 25492 8652 25507
rect 8708 25492 8732 25507
rect 6402 25474 6929 25492
rect 3434 25442 5257 25474
rect 5309 25442 5323 25474
rect 5375 25442 6093 25474
rect 6145 25442 6159 25474
rect 6211 25442 6929 25474
rect 3434 25386 3443 25442
rect 3499 25386 3525 25442
rect 3581 25386 3607 25442
rect 3663 25386 3689 25442
rect 3745 25386 3771 25442
rect 3827 25386 3853 25442
rect 3909 25386 3935 25442
rect 3991 25386 4017 25442
rect 4073 25386 4098 25442
rect 4154 25386 4179 25442
rect 4235 25386 4260 25442
rect 4316 25386 5215 25442
rect 5375 25440 5377 25442
rect 5271 25425 5296 25440
rect 5352 25425 5377 25440
rect 5375 25386 5377 25425
rect 5433 25386 5458 25442
rect 5514 25386 5539 25442
rect 5595 25386 5620 25442
rect 5676 25386 5701 25442
rect 5757 25386 5782 25442
rect 5838 25386 5863 25442
rect 5919 25386 5944 25442
rect 6000 25386 6025 25442
rect 6081 25440 6093 25442
rect 6081 25425 6106 25440
rect 6162 25425 6186 25440
rect 6081 25386 6093 25425
rect 6242 25386 6266 25442
rect 6322 25386 6346 25442
rect 6402 25440 6929 25442
rect 6981 25440 6995 25492
rect 7047 25440 7765 25492
rect 7817 25440 7831 25492
rect 7883 25474 8572 25492
rect 8719 25474 8732 25492
rect 8788 25474 8812 25530
rect 8868 25474 8893 25530
rect 8949 25474 8974 25530
rect 9030 25474 9055 25530
rect 9111 25474 9136 25530
rect 9192 25474 9217 25530
rect 9273 25474 9298 25530
rect 9354 25474 9379 25530
rect 9435 25507 9437 25530
rect 9435 25492 9460 25507
rect 9516 25492 9541 25507
rect 9435 25474 9437 25492
rect 9597 25474 9622 25530
rect 9678 25474 9703 25530
rect 9759 25507 10273 25530
rect 10325 25507 10339 25559
rect 10391 25530 11109 25559
rect 11161 25530 11175 25559
rect 11227 25530 11945 25559
rect 11997 25530 12011 25559
rect 10391 25507 10871 25530
rect 9759 25492 10871 25507
rect 9759 25474 10273 25492
rect 7883 25442 8601 25474
rect 8653 25442 8667 25474
rect 8719 25442 9437 25474
rect 9489 25442 9503 25474
rect 9555 25442 10273 25474
rect 7883 25440 8572 25442
rect 8719 25440 8732 25442
rect 6402 25425 8572 25440
rect 8628 25425 8652 25440
rect 8708 25425 8732 25440
rect 6402 25386 6929 25425
rect 3434 25373 5257 25386
rect 5309 25373 5323 25386
rect 5375 25373 6093 25386
rect 6145 25373 6159 25386
rect 6211 25373 6929 25386
rect 6981 25373 6995 25425
rect 7047 25373 7765 25425
rect 7817 25373 7831 25425
rect 7883 25386 8572 25425
rect 8719 25386 8732 25425
rect 8788 25386 8812 25442
rect 8868 25386 8893 25442
rect 8949 25386 8974 25442
rect 9030 25386 9055 25442
rect 9111 25386 9136 25442
rect 9192 25386 9217 25442
rect 9273 25386 9298 25442
rect 9354 25386 9379 25442
rect 9435 25440 9437 25442
rect 9435 25425 9460 25440
rect 9516 25425 9541 25440
rect 9435 25386 9437 25425
rect 9597 25386 9622 25442
rect 9678 25386 9703 25442
rect 9759 25440 10273 25442
rect 10325 25440 10339 25492
rect 10391 25474 10871 25492
rect 10927 25474 10951 25530
rect 11007 25474 11031 25530
rect 11087 25507 11109 25530
rect 11167 25507 11175 25530
rect 11087 25492 11111 25507
rect 11167 25492 11192 25507
rect 11087 25474 11109 25492
rect 11167 25474 11175 25492
rect 11248 25474 11273 25530
rect 11329 25474 11354 25530
rect 11410 25474 11435 25530
rect 11491 25474 11516 25530
rect 11572 25474 11597 25530
rect 11653 25474 11678 25530
rect 11734 25474 11759 25530
rect 11815 25474 11840 25530
rect 11896 25474 11921 25530
rect 11997 25507 12002 25530
rect 12063 25507 12781 25559
rect 12833 25507 12847 25559
rect 12899 25507 13317 25559
rect 11977 25492 12002 25507
rect 12058 25492 13317 25507
rect 11997 25474 12002 25492
rect 10391 25442 11109 25474
rect 11161 25442 11175 25474
rect 11227 25442 11945 25474
rect 11997 25442 12011 25474
rect 10391 25440 10871 25442
rect 9759 25425 10871 25440
rect 9759 25386 10273 25425
rect 7883 25373 8601 25386
rect 8653 25373 8667 25386
rect 8719 25373 9437 25386
rect 9489 25373 9503 25386
rect 9555 25373 10273 25386
rect 10325 25373 10339 25425
rect 10391 25386 10871 25425
rect 10927 25386 10951 25442
rect 11007 25386 11031 25442
rect 11087 25440 11109 25442
rect 11167 25440 11175 25442
rect 11087 25425 11111 25440
rect 11167 25425 11192 25440
rect 11087 25386 11109 25425
rect 11167 25386 11175 25425
rect 11248 25386 11273 25442
rect 11329 25386 11354 25442
rect 11410 25386 11435 25442
rect 11491 25386 11516 25442
rect 11572 25386 11597 25442
rect 11653 25386 11678 25442
rect 11734 25386 11759 25442
rect 11815 25386 11840 25442
rect 11896 25386 11921 25442
rect 11997 25440 12002 25442
rect 12063 25440 12781 25492
rect 12833 25440 12847 25492
rect 12899 25440 13317 25492
rect 11977 25425 12002 25440
rect 12058 25425 13317 25440
rect 11997 25386 12002 25425
rect 10391 25373 11109 25386
rect 11161 25373 11175 25386
rect 11227 25373 11945 25386
rect 11997 25373 12011 25386
rect 12063 25373 12781 25425
rect 12833 25373 12847 25425
rect 12899 25373 13317 25425
rect 3434 25367 13317 25373
rect 3756 23697 5075 23703
rect 3756 23645 3757 23697
rect 3809 23645 3831 23697
rect 3883 23651 5075 23697
rect 5127 23651 5151 23703
rect 5203 23651 5226 23703
rect 5278 23651 5301 23703
rect 5353 23651 5376 23703
rect 5428 23651 5451 23703
rect 5503 23651 5509 23703
rect 3883 23645 5509 23651
rect 3756 23627 5509 23645
rect 3756 23625 5075 23627
rect 3756 23573 3757 23625
rect 3809 23573 3831 23625
rect 3883 23575 5075 23625
rect 5127 23575 5151 23627
rect 5203 23575 5226 23627
rect 5278 23575 5301 23627
rect 5353 23575 5376 23627
rect 5428 23575 5451 23627
rect 5503 23575 5509 23627
rect 3883 23573 5509 23575
rect 3756 23553 5509 23573
rect 3756 23501 3757 23553
rect 3809 23501 3831 23553
rect 3883 23551 5509 23553
rect 3883 23501 5075 23551
rect 3756 23499 5075 23501
rect 5127 23499 5151 23551
rect 5203 23499 5226 23551
rect 5278 23499 5301 23551
rect 5353 23499 5376 23551
rect 5428 23499 5451 23551
rect 5503 23499 5509 23551
rect 3756 23480 5509 23499
rect 3756 23428 3757 23480
rect 3809 23428 3831 23480
rect 3883 23475 5509 23480
rect 3883 23428 5075 23475
rect 3756 23423 5075 23428
rect 5127 23423 5151 23475
rect 5203 23423 5226 23475
rect 5278 23423 5301 23475
rect 5353 23423 5376 23475
rect 5428 23423 5451 23475
rect 5503 23423 5509 23475
rect 3756 23422 5509 23423
rect 3756 21723 3762 21775
rect 3814 21723 3826 21775
rect 3878 21723 5073 21775
rect 5125 21723 5140 21775
rect 5192 21723 5206 21775
rect 5258 21723 5272 21775
rect 5324 21723 5330 21775
rect 4911 19702 4917 19754
rect 4969 19702 4981 19754
rect 5033 19702 5039 19754
rect 4911 18055 5039 19702
rect 4911 18003 4917 18055
rect 4969 18003 4981 18055
rect 5033 18003 5039 18055
rect 4731 16809 4849 16815
rect 4783 16757 4797 16809
rect 4731 16706 4849 16757
rect 4480 16657 4662 16663
rect 4480 16605 4481 16657
rect 4533 16605 4545 16657
rect 4597 16605 4609 16657
rect 4661 16605 4662 16657
rect 4480 16545 4662 16605
rect 4480 16493 4481 16545
rect 4533 16493 4545 16545
rect 4597 16493 4609 16545
rect 4661 16493 4662 16545
rect 4480 16433 4662 16493
rect 4480 16381 4481 16433
rect 4533 16381 4545 16433
rect 4597 16381 4609 16433
rect 4661 16381 4662 16433
rect 4480 16066 4662 16381
rect 4480 16014 4481 16066
rect 4533 16014 4545 16066
rect 4597 16014 4609 16066
rect 4661 16014 4662 16066
rect 4480 15922 4662 16014
rect 4480 15870 4481 15922
rect 4533 15870 4545 15922
rect 4597 15870 4609 15922
rect 4661 15870 4662 15922
rect 4480 15778 4662 15870
rect 4480 15726 4481 15778
rect 4533 15726 4545 15778
rect 4597 15726 4609 15778
rect 4661 15726 4662 15778
rect 4480 15634 4662 15726
rect 4480 15582 4481 15634
rect 4533 15582 4545 15634
rect 4597 15582 4609 15634
rect 4661 15582 4662 15634
rect 4480 15490 4662 15582
rect 4480 15438 4481 15490
rect 4533 15438 4545 15490
rect 4597 15438 4609 15490
rect 4661 15438 4662 15490
rect 4480 15346 4662 15438
rect 4480 15294 4481 15346
rect 4533 15294 4545 15346
rect 4597 15294 4609 15346
rect 4661 15294 4662 15346
rect 4480 15202 4662 15294
rect 4480 15150 4481 15202
rect 4533 15150 4545 15202
rect 4597 15150 4609 15202
rect 4661 15150 4662 15202
rect 4480 15144 4662 15150
rect 4783 16654 4797 16706
rect 4731 16603 4849 16654
rect 4783 16551 4797 16603
rect 100 14869 2760 14901
tri 2760 14869 2792 14901 nw
rect 4731 15042 4849 16551
rect 4911 16271 5039 18003
rect 4911 16219 4917 16271
rect 4969 16219 4981 16271
rect 5033 16219 5039 16271
rect 4911 16209 5039 16219
rect 13200 19706 13602 19712
rect 13252 19654 13270 19706
rect 13322 19654 13340 19706
rect 13392 19654 13410 19706
rect 13462 19654 13480 19706
rect 13532 19654 13550 19706
rect 13200 19642 13602 19654
rect 13252 19590 13270 19642
rect 13322 19590 13340 19642
rect 13392 19590 13410 19642
rect 13462 19590 13480 19642
rect 13532 19590 13550 19642
rect 13200 19578 13602 19590
rect 13252 19526 13270 19578
rect 13322 19526 13340 19578
rect 13392 19526 13410 19578
rect 13462 19526 13480 19578
rect 13532 19526 13550 19578
rect 13200 19514 13602 19526
rect 13252 19462 13270 19514
rect 13322 19462 13340 19514
rect 13392 19462 13410 19514
rect 13462 19462 13480 19514
rect 13532 19462 13550 19514
rect 13200 19450 13602 19462
rect 13252 19398 13270 19450
rect 13322 19398 13340 19450
rect 13392 19398 13410 19450
rect 13462 19398 13480 19450
rect 13532 19398 13550 19450
rect 13200 19386 13602 19398
rect 13252 19334 13270 19386
rect 13322 19334 13340 19386
rect 13392 19334 13410 19386
rect 13462 19334 13480 19386
rect 13532 19334 13550 19386
rect 13200 19322 13602 19334
rect 13252 19270 13270 19322
rect 13322 19270 13340 19322
rect 13392 19270 13410 19322
rect 13462 19270 13480 19322
rect 13532 19270 13550 19322
rect 13200 19258 13602 19270
rect 13252 19206 13270 19258
rect 13322 19206 13340 19258
rect 13392 19206 13410 19258
rect 13462 19206 13480 19258
rect 13532 19206 13550 19258
rect 13200 19194 13602 19206
rect 13252 19142 13270 19194
rect 13322 19142 13340 19194
rect 13392 19142 13410 19194
rect 13462 19142 13480 19194
rect 13532 19142 13550 19194
rect 13200 19130 13602 19142
rect 13252 19078 13270 19130
rect 13322 19078 13340 19130
rect 13392 19078 13410 19130
rect 13462 19078 13480 19130
rect 13532 19078 13550 19130
rect 13200 19066 13602 19078
rect 13252 19014 13270 19066
rect 13322 19014 13340 19066
rect 13392 19014 13410 19066
rect 13462 19014 13480 19066
rect 13532 19014 13550 19066
rect 13200 19002 13602 19014
rect 13252 18950 13270 19002
rect 13322 18950 13340 19002
rect 13392 18950 13410 19002
rect 13462 18950 13480 19002
rect 13532 18950 13550 19002
rect 13200 18938 13602 18950
rect 13252 18886 13270 18938
rect 13322 18886 13340 18938
rect 13392 18886 13410 18938
rect 13462 18886 13480 18938
rect 13532 18886 13550 18938
rect 13200 18874 13602 18886
rect 13252 18822 13270 18874
rect 13322 18822 13340 18874
rect 13392 18822 13410 18874
rect 13462 18822 13480 18874
rect 13532 18822 13550 18874
rect 13200 18810 13602 18822
rect 13252 18758 13270 18810
rect 13322 18758 13340 18810
rect 13392 18758 13410 18810
rect 13462 18758 13480 18810
rect 13532 18758 13550 18810
rect 13200 18746 13602 18758
rect 13252 18694 13270 18746
rect 13322 18694 13340 18746
rect 13392 18694 13410 18746
rect 13462 18694 13480 18746
rect 13532 18694 13550 18746
rect 13200 18682 13602 18694
rect 13252 18630 13270 18682
rect 13322 18630 13340 18682
rect 13392 18630 13410 18682
rect 13462 18630 13480 18682
rect 13532 18630 13550 18682
rect 13200 18618 13602 18630
rect 13252 18566 13270 18618
rect 13322 18566 13340 18618
rect 13392 18566 13410 18618
rect 13462 18566 13480 18618
rect 13532 18566 13550 18618
rect 13200 18554 13602 18566
rect 13252 18502 13270 18554
rect 13322 18502 13340 18554
rect 13392 18502 13410 18554
rect 13462 18502 13480 18554
rect 13532 18502 13550 18554
rect 13200 18490 13602 18502
rect 13252 18438 13270 18490
rect 13322 18438 13340 18490
rect 13392 18438 13410 18490
rect 13462 18438 13480 18490
rect 13532 18438 13550 18490
rect 13200 18426 13602 18438
rect 13252 18374 13270 18426
rect 13322 18374 13340 18426
rect 13392 18374 13410 18426
rect 13462 18374 13480 18426
rect 13532 18374 13550 18426
rect 13200 18362 13602 18374
rect 13252 18310 13270 18362
rect 13322 18310 13340 18362
rect 13392 18310 13410 18362
rect 13462 18310 13480 18362
rect 13532 18310 13550 18362
rect 13200 18298 13602 18310
rect 13252 18246 13270 18298
rect 13322 18246 13340 18298
rect 13392 18246 13410 18298
rect 13462 18246 13480 18298
rect 13532 18246 13550 18298
rect 13200 18234 13602 18246
rect 13252 18182 13270 18234
rect 13322 18182 13340 18234
rect 13392 18182 13410 18234
rect 13462 18182 13480 18234
rect 13532 18182 13550 18234
rect 13200 18170 13602 18182
rect 13252 18118 13270 18170
rect 13322 18118 13340 18170
rect 13392 18118 13410 18170
rect 13462 18118 13480 18170
rect 13532 18118 13550 18170
rect 13200 18106 13602 18118
rect 13252 18054 13270 18106
rect 13322 18054 13340 18106
rect 13392 18054 13410 18106
rect 13462 18054 13480 18106
rect 13532 18054 13550 18106
rect 13200 18042 13602 18054
rect 13252 17990 13270 18042
rect 13322 17990 13340 18042
rect 13392 17990 13410 18042
rect 13462 17990 13480 18042
rect 13532 17990 13550 18042
rect 13200 17978 13602 17990
rect 13252 17926 13270 17978
rect 13322 17926 13340 17978
rect 13392 17926 13410 17978
rect 13462 17926 13480 17978
rect 13532 17926 13550 17978
rect 13200 17914 13602 17926
rect 13252 17862 13270 17914
rect 13322 17862 13340 17914
rect 13392 17862 13410 17914
rect 13462 17862 13480 17914
rect 13532 17862 13550 17914
rect 13200 17850 13602 17862
rect 13252 17798 13270 17850
rect 13322 17798 13340 17850
rect 13392 17798 13410 17850
rect 13462 17798 13480 17850
rect 13532 17798 13550 17850
rect 13200 17786 13602 17798
rect 13252 17734 13270 17786
rect 13322 17734 13340 17786
rect 13392 17734 13410 17786
rect 13462 17734 13480 17786
rect 13532 17734 13550 17786
rect 13200 17722 13602 17734
rect 13252 17670 13270 17722
rect 13322 17670 13340 17722
rect 13392 17670 13410 17722
rect 13462 17670 13480 17722
rect 13532 17670 13550 17722
rect 13200 17658 13602 17670
rect 13252 17606 13270 17658
rect 13322 17606 13340 17658
rect 13392 17606 13410 17658
rect 13462 17606 13480 17658
rect 13532 17606 13550 17658
rect 13200 17594 13602 17606
rect 13252 17542 13270 17594
rect 13322 17542 13340 17594
rect 13392 17542 13410 17594
rect 13462 17542 13480 17594
rect 13532 17542 13550 17594
rect 13200 17530 13602 17542
rect 13252 17478 13270 17530
rect 13322 17478 13340 17530
rect 13392 17478 13410 17530
rect 13462 17478 13480 17530
rect 13532 17478 13550 17530
rect 13200 17466 13602 17478
rect 13252 17414 13270 17466
rect 13322 17414 13340 17466
rect 13392 17414 13410 17466
rect 13462 17414 13480 17466
rect 13532 17414 13550 17466
rect 13200 17402 13602 17414
rect 13252 17350 13270 17402
rect 13322 17350 13340 17402
rect 13392 17350 13410 17402
rect 13462 17350 13480 17402
rect 13532 17350 13550 17402
rect 13200 17338 13602 17350
rect 13252 17286 13270 17338
rect 13322 17286 13340 17338
rect 13392 17286 13410 17338
rect 13462 17286 13480 17338
rect 13532 17286 13550 17338
rect 13200 17274 13602 17286
rect 13252 17222 13270 17274
rect 13322 17222 13340 17274
rect 13392 17222 13410 17274
rect 13462 17222 13480 17274
rect 13532 17222 13550 17274
rect 13200 17210 13602 17222
rect 13252 17158 13270 17210
rect 13322 17158 13340 17210
rect 13392 17158 13410 17210
rect 13462 17158 13480 17210
rect 13532 17158 13550 17210
rect 13200 17146 13602 17158
rect 13252 17094 13270 17146
rect 13322 17094 13340 17146
rect 13392 17094 13410 17146
rect 13462 17094 13480 17146
rect 13532 17094 13550 17146
rect 13200 17082 13602 17094
rect 13252 17030 13270 17082
rect 13322 17030 13340 17082
rect 13392 17030 13410 17082
rect 13462 17030 13480 17082
rect 13532 17030 13550 17082
rect 13200 17018 13602 17030
rect 13252 16966 13270 17018
rect 13322 16966 13340 17018
rect 13392 16966 13410 17018
rect 13462 16966 13480 17018
rect 13532 16966 13550 17018
rect 13200 16954 13602 16966
rect 13252 16902 13270 16954
rect 13322 16902 13340 16954
rect 13392 16902 13410 16954
rect 13462 16902 13480 16954
rect 13532 16902 13550 16954
rect 13200 16890 13602 16902
rect 13252 16838 13270 16890
rect 13322 16838 13340 16890
rect 13392 16838 13410 16890
rect 13462 16838 13480 16890
rect 13532 16838 13550 16890
rect 13200 16826 13602 16838
rect 13252 16774 13270 16826
rect 13322 16774 13340 16826
rect 13392 16774 13410 16826
rect 13462 16774 13480 16826
rect 13532 16774 13550 16826
rect 13200 16762 13602 16774
rect 13252 16710 13270 16762
rect 13322 16710 13340 16762
rect 13392 16710 13410 16762
rect 13462 16710 13480 16762
rect 13532 16710 13550 16762
rect 13200 16698 13602 16710
rect 13252 16646 13270 16698
rect 13322 16646 13340 16698
rect 13392 16646 13410 16698
rect 13462 16646 13480 16698
rect 13532 16646 13550 16698
rect 13200 16634 13602 16646
rect 13252 16582 13270 16634
rect 13322 16582 13340 16634
rect 13392 16582 13410 16634
rect 13462 16582 13480 16634
rect 13532 16582 13550 16634
rect 13200 16570 13602 16582
rect 13252 16518 13270 16570
rect 13322 16518 13340 16570
rect 13392 16518 13410 16570
rect 13462 16518 13480 16570
rect 13532 16518 13550 16570
rect 13200 16506 13602 16518
rect 13252 16454 13270 16506
rect 13322 16454 13340 16506
rect 13392 16454 13410 16506
rect 13462 16454 13480 16506
rect 13532 16454 13550 16506
rect 13200 16442 13602 16454
rect 13252 16390 13270 16442
rect 13322 16390 13340 16442
rect 13392 16390 13410 16442
rect 13462 16390 13480 16442
rect 13532 16390 13550 16442
rect 13200 16378 13602 16390
rect 13252 16326 13270 16378
rect 13322 16326 13340 16378
rect 13392 16326 13410 16378
rect 13462 16326 13480 16378
rect 13532 16326 13550 16378
rect 13200 16314 13602 16326
rect 13252 16262 13270 16314
rect 13322 16262 13340 16314
rect 13392 16262 13410 16314
rect 13462 16262 13480 16314
rect 13532 16262 13550 16314
rect 13200 16250 13602 16262
rect 4783 14990 4797 15042
rect 4731 14921 4849 14990
rect 4783 14869 4797 14921
rect 13252 16198 13270 16250
rect 13322 16198 13340 16250
rect 13392 16198 13410 16250
rect 13462 16198 13480 16250
rect 13532 16198 13550 16250
rect 13200 16186 13602 16198
rect 13252 16134 13270 16186
rect 13322 16134 13340 16186
rect 13392 16134 13410 16186
rect 13462 16134 13480 16186
rect 13532 16134 13550 16186
rect 13200 16122 13602 16134
rect 13252 16070 13270 16122
rect 13322 16070 13340 16122
rect 13392 16070 13410 16122
rect 13462 16070 13480 16122
rect 13532 16070 13550 16122
rect 13200 16058 13602 16070
rect 13252 16006 13270 16058
rect 13322 16006 13340 16058
rect 13392 16006 13410 16058
rect 13462 16006 13480 16058
rect 13532 16006 13550 16058
rect 13200 15994 13602 16006
rect 13252 15942 13270 15994
rect 13322 15942 13340 15994
rect 13392 15942 13410 15994
rect 13462 15942 13480 15994
rect 13532 15942 13550 15994
rect 13200 15930 13602 15942
rect 13252 15878 13270 15930
rect 13322 15878 13340 15930
rect 13392 15878 13410 15930
rect 13462 15878 13480 15930
rect 13532 15878 13550 15930
rect 13200 15866 13602 15878
rect 13252 15814 13270 15866
rect 13322 15814 13340 15866
rect 13392 15814 13410 15866
rect 13462 15814 13480 15866
rect 13532 15814 13550 15866
rect 13200 15802 13602 15814
rect 13252 15750 13270 15802
rect 13322 15750 13340 15802
rect 13392 15750 13410 15802
rect 13462 15750 13480 15802
rect 13532 15750 13550 15802
rect 13200 15738 13602 15750
rect 13252 15686 13270 15738
rect 13322 15686 13340 15738
rect 13392 15686 13410 15738
rect 13462 15686 13480 15738
rect 13532 15686 13550 15738
rect 13200 15674 13602 15686
rect 13252 15622 13270 15674
rect 13322 15622 13340 15674
rect 13392 15622 13410 15674
rect 13462 15622 13480 15674
rect 13532 15622 13550 15674
rect 13200 15610 13602 15622
rect 13252 15558 13270 15610
rect 13322 15558 13340 15610
rect 13392 15558 13410 15610
rect 13462 15558 13480 15610
rect 13532 15558 13550 15610
rect 13200 15546 13602 15558
rect 13252 15494 13270 15546
rect 13322 15494 13340 15546
rect 13392 15494 13410 15546
rect 13462 15494 13480 15546
rect 13532 15494 13550 15546
rect 13200 15482 13602 15494
rect 13252 15430 13270 15482
rect 13322 15430 13340 15482
rect 13392 15430 13410 15482
rect 13462 15430 13480 15482
rect 13532 15430 13550 15482
rect 13200 15418 13602 15430
rect 13252 15366 13270 15418
rect 13322 15366 13340 15418
rect 13392 15366 13410 15418
rect 13462 15366 13480 15418
rect 13532 15366 13550 15418
rect 13200 15354 13602 15366
rect 13252 15302 13270 15354
rect 13322 15302 13340 15354
rect 13392 15302 13410 15354
rect 13462 15302 13480 15354
rect 13532 15302 13550 15354
rect 13200 15290 13602 15302
rect 13252 15238 13270 15290
rect 13322 15238 13340 15290
rect 13392 15238 13410 15290
rect 13462 15238 13480 15290
rect 13532 15238 13550 15290
rect 13200 15226 13602 15238
rect 13252 15174 13270 15226
rect 13322 15174 13340 15226
rect 13392 15174 13410 15226
rect 13462 15174 13480 15226
rect 13532 15174 13550 15226
rect 13200 15162 13602 15174
rect 13252 15110 13270 15162
rect 13322 15110 13340 15162
rect 13392 15110 13410 15162
rect 13462 15110 13480 15162
rect 13532 15110 13550 15162
rect 13200 15098 13602 15110
rect 13252 15046 13270 15098
rect 13322 15046 13340 15098
rect 13392 15046 13410 15098
rect 13462 15046 13480 15098
rect 13532 15046 13550 15098
rect 13200 15034 13602 15046
rect 13252 14982 13270 15034
rect 13322 14982 13340 15034
rect 13392 14982 13410 15034
rect 13462 14982 13480 15034
rect 13532 14982 13550 15034
rect 13200 14970 13602 14982
rect 13252 14918 13270 14970
rect 13322 14918 13340 14970
rect 13392 14918 13410 14970
rect 13462 14918 13480 14970
rect 13532 14918 13550 14970
rect 13200 14906 13602 14918
rect 100 14863 2754 14869
tri 2754 14863 2760 14869 nw
rect 4731 14863 4849 14869
tri 13177 14863 13200 14886 se
rect 100 4997 2750 14863
tri 2750 14859 2754 14863 nw
tri 13173 14859 13177 14863 se
rect 13177 14859 13200 14863
tri 13168 14854 13173 14859 se
rect 13173 14854 13200 14859
rect 13252 14854 13270 14906
rect 13322 14854 13340 14906
rect 13392 14854 13410 14906
rect 13462 14854 13480 14906
rect 13532 14854 13550 14906
tri 13602 14863 13625 14886 sw
rect 13602 14854 13625 14863
tri 13156 14842 13168 14854 se
rect 13168 14842 13625 14854
tri 13104 14790 13156 14842 se
rect 13156 14790 13200 14842
rect 13252 14790 13270 14842
rect 13322 14790 13340 14842
rect 13392 14790 13410 14842
rect 13462 14790 13480 14842
rect 13532 14790 13550 14842
rect 13602 14790 13625 14842
tri 13092 14778 13104 14790 se
rect 13104 14778 13625 14790
tri 13040 14726 13092 14778 se
rect 13092 14726 13200 14778
rect 13252 14726 13270 14778
rect 13322 14726 13340 14778
rect 13392 14726 13410 14778
rect 13462 14726 13480 14778
rect 13532 14726 13550 14778
rect 13602 14726 13625 14778
tri 13625 14726 13762 14863 sw
rect 3227 14720 14940 14726
rect 3279 14668 3293 14720
rect 3345 14668 3781 14720
rect 3833 14668 3847 14720
rect 3899 14668 4335 14720
rect 4387 14668 4401 14720
rect 4453 14668 4889 14720
rect 4941 14668 4955 14720
rect 5007 14668 5443 14720
rect 5495 14668 5509 14720
rect 5561 14668 5997 14720
rect 6049 14668 6063 14720
rect 6115 14668 6551 14720
rect 6603 14668 6617 14720
rect 6669 14668 7105 14720
rect 7157 14668 7171 14720
rect 7223 14668 7659 14720
rect 7711 14668 7725 14720
rect 7777 14668 8213 14720
rect 8265 14668 8279 14720
rect 8331 14668 8767 14720
rect 8819 14668 8833 14720
rect 8885 14668 9321 14720
rect 9373 14668 9387 14720
rect 9439 14668 9875 14720
rect 9927 14668 9941 14720
rect 9993 14668 10429 14720
rect 10481 14668 10495 14720
rect 10547 14668 10983 14720
rect 11035 14668 11049 14720
rect 11101 14668 11537 14720
rect 11589 14668 11603 14720
rect 11655 14668 12091 14720
rect 12143 14668 12157 14720
rect 12209 14668 12645 14720
rect 12697 14668 12711 14720
rect 12763 14714 14940 14720
rect 12763 14668 13200 14714
rect 3227 14662 13200 14668
rect 13252 14662 13270 14714
rect 13322 14662 13340 14714
rect 13392 14662 13410 14714
rect 13462 14662 13480 14714
rect 13532 14662 13550 14714
rect 13602 14662 14940 14714
rect 3227 14654 14940 14662
rect 3279 14602 3293 14654
rect 3345 14602 3781 14654
rect 3833 14602 3847 14654
rect 3899 14602 4335 14654
rect 4387 14602 4401 14654
rect 4453 14602 4889 14654
rect 4941 14602 4955 14654
rect 5007 14602 5443 14654
rect 5495 14602 5509 14654
rect 5561 14602 5997 14654
rect 6049 14602 6063 14654
rect 6115 14602 6551 14654
rect 6603 14602 6617 14654
rect 6669 14602 7105 14654
rect 7157 14602 7171 14654
rect 7223 14602 7659 14654
rect 7711 14602 7725 14654
rect 7777 14602 8213 14654
rect 8265 14602 8279 14654
rect 8331 14602 8767 14654
rect 8819 14602 8833 14654
rect 8885 14602 9321 14654
rect 9373 14602 9387 14654
rect 9439 14602 9875 14654
rect 9927 14602 9941 14654
rect 9993 14602 10429 14654
rect 10481 14602 10495 14654
rect 10547 14602 10983 14654
rect 11035 14602 11049 14654
rect 11101 14602 11537 14654
rect 11589 14602 11603 14654
rect 11655 14602 12091 14654
rect 12143 14602 12157 14654
rect 12209 14602 12645 14654
rect 12697 14602 12711 14654
rect 12763 14650 14940 14654
rect 12763 14602 13200 14650
rect 3227 14598 13200 14602
rect 13252 14598 13270 14650
rect 13322 14598 13340 14650
rect 13392 14598 13410 14650
rect 13462 14598 13480 14650
rect 13532 14598 13550 14650
rect 13602 14598 14940 14650
rect 3227 14588 14940 14598
rect 3279 14536 3293 14588
rect 3345 14536 3781 14588
rect 3833 14536 3847 14588
rect 3899 14536 4335 14588
rect 4387 14536 4401 14588
rect 4453 14536 4889 14588
rect 4941 14536 4955 14588
rect 5007 14536 5443 14588
rect 5495 14536 5509 14588
rect 5561 14536 5997 14588
rect 6049 14536 6063 14588
rect 6115 14536 6551 14588
rect 6603 14536 6617 14588
rect 6669 14536 7105 14588
rect 7157 14536 7171 14588
rect 7223 14536 7659 14588
rect 7711 14536 7725 14588
rect 7777 14536 8213 14588
rect 8265 14536 8279 14588
rect 8331 14536 8767 14588
rect 8819 14536 8833 14588
rect 8885 14536 9321 14588
rect 9373 14536 9387 14588
rect 9439 14536 9875 14588
rect 9927 14536 9941 14588
rect 9993 14536 10429 14588
rect 10481 14536 10495 14588
rect 10547 14536 10983 14588
rect 11035 14536 11049 14588
rect 11101 14536 11537 14588
rect 11589 14536 11603 14588
rect 11655 14536 12091 14588
rect 12143 14536 12157 14588
rect 12209 14536 12645 14588
rect 12697 14536 12711 14588
rect 12763 14586 14940 14588
rect 12763 14536 13200 14586
rect 3227 14534 13200 14536
rect 13252 14534 13270 14586
rect 13322 14534 13340 14586
rect 13392 14534 13410 14586
rect 13462 14534 13480 14586
rect 13532 14534 13550 14586
rect 13602 14534 14940 14586
rect 3227 14522 14940 14534
rect 3279 14470 3293 14522
rect 3345 14470 3781 14522
rect 3833 14470 3847 14522
rect 3899 14470 4335 14522
rect 4387 14470 4401 14522
rect 4453 14470 4889 14522
rect 4941 14470 4955 14522
rect 5007 14470 5443 14522
rect 5495 14470 5509 14522
rect 5561 14470 5997 14522
rect 6049 14470 6063 14522
rect 6115 14470 6551 14522
rect 6603 14470 6617 14522
rect 6669 14470 7105 14522
rect 7157 14470 7171 14522
rect 7223 14470 7659 14522
rect 7711 14470 7725 14522
rect 7777 14470 8213 14522
rect 8265 14470 8279 14522
rect 8331 14470 8767 14522
rect 8819 14470 8833 14522
rect 8885 14470 9321 14522
rect 9373 14470 9387 14522
rect 9439 14470 9875 14522
rect 9927 14470 9941 14522
rect 9993 14470 10429 14522
rect 10481 14470 10495 14522
rect 10547 14470 10983 14522
rect 11035 14470 11049 14522
rect 11101 14470 11537 14522
rect 11589 14470 11603 14522
rect 11655 14470 12091 14522
rect 12143 14470 12157 14522
rect 12209 14470 12645 14522
rect 12697 14470 12711 14522
rect 12763 14470 13200 14522
rect 13252 14470 13270 14522
rect 13322 14470 13340 14522
rect 13392 14470 13410 14522
rect 13462 14470 13480 14522
rect 13532 14470 13550 14522
rect 13602 14470 14940 14522
rect 3227 14458 14940 14470
rect 3227 14456 13200 14458
rect 3279 14404 3293 14456
rect 3345 14404 3781 14456
rect 3833 14404 3847 14456
rect 3899 14404 4335 14456
rect 4387 14404 4401 14456
rect 4453 14404 4889 14456
rect 4941 14404 4955 14456
rect 5007 14404 5443 14456
rect 5495 14404 5509 14456
rect 5561 14404 5997 14456
rect 6049 14404 6063 14456
rect 6115 14404 6551 14456
rect 6603 14404 6617 14456
rect 6669 14404 7105 14456
rect 7157 14404 7171 14456
rect 7223 14404 7659 14456
rect 7711 14404 7725 14456
rect 7777 14404 8213 14456
rect 8265 14404 8279 14456
rect 8331 14404 8767 14456
rect 8819 14404 8833 14456
rect 8885 14404 9321 14456
rect 9373 14404 9387 14456
rect 9439 14404 9875 14456
rect 9927 14404 9941 14456
rect 9993 14404 10429 14456
rect 10481 14404 10495 14456
rect 10547 14404 10983 14456
rect 11035 14404 11049 14456
rect 11101 14404 11537 14456
rect 11589 14404 11603 14456
rect 11655 14404 12091 14456
rect 12143 14404 12157 14456
rect 12209 14404 12645 14456
rect 12697 14404 12711 14456
rect 12763 14406 13200 14456
rect 13252 14406 13270 14458
rect 13322 14406 13340 14458
rect 13392 14406 13410 14458
rect 13462 14406 13480 14458
rect 13532 14406 13550 14458
rect 13602 14406 14940 14458
rect 12763 14404 14940 14406
rect 3227 14394 14940 14404
rect 3227 14390 13200 14394
rect 3279 14338 3293 14390
rect 3345 14338 3781 14390
rect 3833 14338 3847 14390
rect 3899 14338 4335 14390
rect 4387 14338 4401 14390
rect 4453 14338 4889 14390
rect 4941 14338 4955 14390
rect 5007 14338 5443 14390
rect 5495 14338 5509 14390
rect 5561 14338 5997 14390
rect 6049 14338 6063 14390
rect 6115 14338 6551 14390
rect 6603 14338 6617 14390
rect 6669 14338 7105 14390
rect 7157 14338 7171 14390
rect 7223 14338 7659 14390
rect 7711 14338 7725 14390
rect 7777 14338 8213 14390
rect 8265 14338 8279 14390
rect 8331 14338 8767 14390
rect 8819 14338 8833 14390
rect 8885 14338 9321 14390
rect 9373 14338 9387 14390
rect 9439 14338 9875 14390
rect 9927 14338 9941 14390
rect 9993 14338 10429 14390
rect 10481 14338 10495 14390
rect 10547 14338 10983 14390
rect 11035 14338 11049 14390
rect 11101 14338 11537 14390
rect 11589 14338 11603 14390
rect 11655 14338 12091 14390
rect 12143 14338 12157 14390
rect 12209 14338 12645 14390
rect 12697 14338 12711 14390
rect 12763 14342 13200 14390
rect 13252 14342 13270 14394
rect 13322 14342 13340 14394
rect 13392 14342 13410 14394
rect 13462 14342 13480 14394
rect 13532 14342 13550 14394
rect 13602 14342 14940 14394
rect 12763 14338 14940 14342
rect 3227 14330 14940 14338
rect 3227 14323 13200 14330
rect 3279 14271 3293 14323
rect 3345 14271 3781 14323
rect 3833 14271 3847 14323
rect 3899 14271 4335 14323
rect 4387 14271 4401 14323
rect 4453 14271 4889 14323
rect 4941 14271 4955 14323
rect 5007 14271 5443 14323
rect 5495 14271 5509 14323
rect 5561 14271 5997 14323
rect 6049 14271 6063 14323
rect 6115 14271 6551 14323
rect 6603 14271 6617 14323
rect 6669 14271 7105 14323
rect 7157 14271 7171 14323
rect 7223 14271 7659 14323
rect 7711 14271 7725 14323
rect 7777 14271 8213 14323
rect 8265 14271 8279 14323
rect 8331 14271 8767 14323
rect 8819 14271 8833 14323
rect 8885 14271 9321 14323
rect 9373 14271 9387 14323
rect 9439 14271 9875 14323
rect 9927 14271 9941 14323
rect 9993 14271 10429 14323
rect 10481 14271 10495 14323
rect 10547 14271 10983 14323
rect 11035 14271 11049 14323
rect 11101 14271 11537 14323
rect 11589 14271 11603 14323
rect 11655 14271 12091 14323
rect 12143 14271 12157 14323
rect 12209 14271 12645 14323
rect 12697 14271 12711 14323
rect 12763 14278 13200 14323
rect 13252 14278 13270 14330
rect 13322 14278 13340 14330
rect 13392 14278 13410 14330
rect 13462 14278 13480 14330
rect 13532 14278 13550 14330
rect 13602 14278 14940 14330
rect 12763 14271 14940 14278
rect 3227 14266 14940 14271
rect 3227 14256 13200 14266
rect 3279 14204 3293 14256
rect 3345 14204 3781 14256
rect 3833 14204 3847 14256
rect 3899 14204 4335 14256
rect 4387 14204 4401 14256
rect 4453 14204 4889 14256
rect 4941 14204 4955 14256
rect 5007 14204 5443 14256
rect 5495 14204 5509 14256
rect 5561 14204 5997 14256
rect 6049 14204 6063 14256
rect 6115 14204 6551 14256
rect 6603 14204 6617 14256
rect 6669 14204 7105 14256
rect 7157 14204 7171 14256
rect 7223 14204 7659 14256
rect 7711 14204 7725 14256
rect 7777 14204 8213 14256
rect 8265 14204 8279 14256
rect 8331 14204 8767 14256
rect 8819 14204 8833 14256
rect 8885 14204 9321 14256
rect 9373 14204 9387 14256
rect 9439 14204 9875 14256
rect 9927 14204 9941 14256
rect 9993 14204 10429 14256
rect 10481 14204 10495 14256
rect 10547 14204 10983 14256
rect 11035 14204 11049 14256
rect 11101 14204 11537 14256
rect 11589 14204 11603 14256
rect 11655 14204 12091 14256
rect 12143 14204 12157 14256
rect 12209 14204 12645 14256
rect 12697 14204 12711 14256
rect 12763 14214 13200 14256
rect 13252 14214 13270 14266
rect 13322 14214 13340 14266
rect 13392 14214 13410 14266
rect 13462 14214 13480 14266
rect 13532 14214 13550 14266
rect 13602 14214 14940 14266
rect 12763 14204 14940 14214
rect 3227 14202 14940 14204
rect 3227 14198 13200 14202
tri 12989 14150 13037 14198 ne
rect 13037 14150 13200 14198
rect 13252 14150 13270 14202
rect 13322 14150 13340 14202
rect 13392 14150 13410 14202
rect 13462 14150 13480 14202
rect 13532 14150 13550 14202
rect 13602 14150 14940 14202
tri 13037 14138 13049 14150 ne
rect 13049 14138 14940 14150
tri 13049 14086 13101 14138 ne
rect 13101 14086 13200 14138
rect 13252 14086 13270 14138
rect 13322 14086 13340 14138
rect 13392 14086 13410 14138
rect 13462 14086 13480 14138
rect 13532 14086 13550 14138
rect 13602 14086 14940 14138
tri 13101 14074 13113 14086 ne
rect 13113 14074 14940 14086
tri 13113 14022 13165 14074 ne
rect 13165 14022 13200 14074
rect 13252 14022 13270 14074
rect 13322 14022 13340 14074
rect 13392 14022 13410 14074
rect 13462 14022 13480 14074
rect 13532 14022 13550 14074
rect 13602 14022 14940 14074
tri 13165 14010 13177 14022 ne
rect 13177 14010 14940 14022
tri 13177 13988 13199 14010 ne
rect 13199 13958 13200 14010
rect 13252 13958 13270 14010
rect 13322 13958 13340 14010
rect 13392 13958 13410 14010
rect 13462 13958 13480 14010
rect 13532 13958 13550 14010
rect 13602 13958 14940 14010
rect 13199 13946 14940 13958
rect 2950 13892 13040 13898
rect 3002 13840 3016 13892
rect 3068 13840 3504 13892
rect 3556 13840 3570 13892
rect 3622 13840 4058 13892
rect 4110 13840 4124 13892
rect 4176 13840 4612 13892
rect 4664 13840 4678 13892
rect 4730 13840 5166 13892
rect 5218 13840 5232 13892
rect 5284 13840 5720 13892
rect 5772 13840 5786 13892
rect 5838 13840 6274 13892
rect 6326 13840 6340 13892
rect 6392 13840 6828 13892
rect 6880 13840 6894 13892
rect 6946 13840 7382 13892
rect 7434 13840 7448 13892
rect 7500 13877 7936 13892
rect 7988 13877 8002 13892
rect 8054 13877 8490 13892
rect 8542 13877 8556 13892
rect 8608 13877 9044 13892
rect 9096 13877 9110 13892
rect 9162 13877 9598 13892
rect 9650 13877 9664 13892
rect 9716 13877 10152 13892
rect 7500 13840 7691 13877
rect 2950 13826 7691 13840
rect 3002 13774 3016 13826
rect 3068 13774 3504 13826
rect 3556 13774 3570 13826
rect 3622 13774 4058 13826
rect 4110 13774 4124 13826
rect 4176 13774 4612 13826
rect 4664 13774 4678 13826
rect 4730 13774 5166 13826
rect 5218 13774 5232 13826
rect 5284 13774 5720 13826
rect 5772 13774 5786 13826
rect 5838 13774 6274 13826
rect 6326 13774 6340 13826
rect 6392 13774 6828 13826
rect 6880 13774 6894 13826
rect 6946 13774 7382 13826
rect 7434 13774 7448 13826
rect 7500 13821 7691 13826
rect 7747 13821 7775 13877
rect 7831 13821 7858 13877
rect 7914 13840 7936 13877
rect 7997 13840 8002 13877
rect 7914 13826 7941 13840
rect 7997 13826 8024 13840
rect 7914 13821 7936 13826
rect 7997 13821 8002 13826
rect 8080 13821 8107 13877
rect 8163 13821 8190 13877
rect 8246 13821 8273 13877
rect 8329 13821 8356 13877
rect 8412 13821 8439 13877
rect 8495 13826 8522 13840
rect 8578 13826 8605 13840
rect 8661 13821 8688 13877
rect 8744 13821 8771 13877
rect 8827 13821 8854 13877
rect 8910 13821 8937 13877
rect 8993 13821 9020 13877
rect 9096 13840 9103 13877
rect 9162 13840 9186 13877
rect 9076 13826 9103 13840
rect 9159 13826 9186 13840
rect 9096 13821 9103 13826
rect 9162 13821 9186 13826
rect 9242 13821 9269 13877
rect 9325 13821 9352 13877
rect 9408 13821 9435 13877
rect 9491 13821 9518 13877
rect 9574 13840 9598 13877
rect 9657 13840 9664 13877
rect 9574 13826 9601 13840
rect 9657 13826 9684 13840
rect 9574 13821 9598 13826
rect 9657 13821 9664 13826
rect 9740 13821 9767 13877
rect 9823 13840 10152 13877
rect 10204 13840 10218 13892
rect 10270 13840 10706 13892
rect 10758 13840 10772 13892
rect 10824 13840 11260 13892
rect 11312 13840 11326 13892
rect 11378 13840 11814 13892
rect 11866 13840 11880 13892
rect 11932 13840 12368 13892
rect 12420 13840 12434 13892
rect 12486 13840 12922 13892
rect 12974 13840 12988 13892
rect 9823 13826 13040 13840
rect 9823 13821 10152 13826
rect 7500 13789 7936 13821
rect 7988 13789 8002 13821
rect 8054 13789 8490 13821
rect 8542 13789 8556 13821
rect 8608 13789 9044 13821
rect 9096 13789 9110 13821
rect 9162 13789 9598 13821
rect 9650 13789 9664 13821
rect 9716 13789 10152 13821
rect 7500 13774 7691 13789
rect 2950 13760 7691 13774
rect 3002 13708 3016 13760
rect 3068 13708 3504 13760
rect 3556 13708 3570 13760
rect 3622 13708 4058 13760
rect 4110 13708 4124 13760
rect 4176 13708 4612 13760
rect 4664 13708 4678 13760
rect 4730 13708 5166 13760
rect 5218 13708 5232 13760
rect 5284 13708 5720 13760
rect 5772 13708 5786 13760
rect 5838 13708 6274 13760
rect 6326 13708 6340 13760
rect 6392 13708 6828 13760
rect 6880 13708 6894 13760
rect 6946 13708 7382 13760
rect 7434 13708 7448 13760
rect 7500 13733 7691 13760
rect 7747 13733 7775 13789
rect 7831 13733 7858 13789
rect 7914 13774 7936 13789
rect 7997 13774 8002 13789
rect 7914 13760 7941 13774
rect 7997 13760 8024 13774
rect 7914 13733 7936 13760
rect 7997 13733 8002 13760
rect 8080 13733 8107 13789
rect 8163 13733 8190 13789
rect 8246 13733 8273 13789
rect 8329 13733 8356 13789
rect 8412 13733 8439 13789
rect 8495 13760 8522 13774
rect 8578 13760 8605 13774
rect 8661 13733 8688 13789
rect 8744 13733 8771 13789
rect 8827 13733 8854 13789
rect 8910 13733 8937 13789
rect 8993 13733 9020 13789
rect 9096 13774 9103 13789
rect 9162 13774 9186 13789
rect 9076 13760 9103 13774
rect 9159 13760 9186 13774
rect 9096 13733 9103 13760
rect 9162 13733 9186 13760
rect 9242 13733 9269 13789
rect 9325 13733 9352 13789
rect 9408 13733 9435 13789
rect 9491 13733 9518 13789
rect 9574 13774 9598 13789
rect 9657 13774 9664 13789
rect 9574 13760 9601 13774
rect 9657 13760 9684 13774
rect 9574 13733 9598 13760
rect 9657 13733 9664 13760
rect 9740 13733 9767 13789
rect 9823 13774 10152 13789
rect 10204 13774 10218 13826
rect 10270 13774 10706 13826
rect 10758 13774 10772 13826
rect 10824 13774 11260 13826
rect 11312 13774 11326 13826
rect 11378 13774 11814 13826
rect 11866 13774 11880 13826
rect 11932 13774 12368 13826
rect 12420 13774 12434 13826
rect 12486 13774 12922 13826
rect 12974 13774 12988 13826
rect 9823 13760 13040 13774
rect 9823 13733 10152 13760
rect 7500 13708 7936 13733
rect 7988 13708 8002 13733
rect 8054 13708 8490 13733
rect 8542 13708 8556 13733
rect 8608 13708 9044 13733
rect 9096 13708 9110 13733
rect 9162 13708 9598 13733
rect 9650 13708 9664 13733
rect 9716 13708 10152 13733
rect 10204 13708 10218 13760
rect 10270 13708 10706 13760
rect 10758 13708 10772 13760
rect 10824 13708 11260 13760
rect 11312 13708 11326 13760
rect 11378 13708 11814 13760
rect 11866 13708 11880 13760
rect 11932 13708 12368 13760
rect 12420 13708 12434 13760
rect 12486 13708 12922 13760
rect 12974 13708 12988 13760
rect 2950 13701 13040 13708
rect 2950 13694 7691 13701
rect 3002 13642 3016 13694
rect 3068 13642 3504 13694
rect 3556 13642 3570 13694
rect 3622 13642 4058 13694
rect 4110 13642 4124 13694
rect 4176 13642 4612 13694
rect 4664 13642 4678 13694
rect 4730 13642 5166 13694
rect 5218 13642 5232 13694
rect 5284 13642 5720 13694
rect 5772 13642 5786 13694
rect 5838 13642 6274 13694
rect 6326 13642 6340 13694
rect 6392 13642 6828 13694
rect 6880 13642 6894 13694
rect 6946 13642 7382 13694
rect 7434 13642 7448 13694
rect 7500 13645 7691 13694
rect 7747 13645 7775 13701
rect 7831 13645 7858 13701
rect 7914 13694 7941 13701
rect 7997 13694 8024 13701
rect 7914 13645 7936 13694
rect 7997 13645 8002 13694
rect 8080 13645 8107 13701
rect 8163 13645 8190 13701
rect 8246 13645 8273 13701
rect 8329 13645 8356 13701
rect 8412 13645 8439 13701
rect 8495 13694 8522 13701
rect 8578 13694 8605 13701
rect 8661 13645 8688 13701
rect 8744 13645 8771 13701
rect 8827 13645 8854 13701
rect 8910 13645 8937 13701
rect 8993 13645 9020 13701
rect 9076 13694 9103 13701
rect 9159 13694 9186 13701
rect 9096 13645 9103 13694
rect 9162 13645 9186 13694
rect 9242 13645 9269 13701
rect 9325 13645 9352 13701
rect 9408 13645 9435 13701
rect 9491 13645 9518 13701
rect 9574 13694 9601 13701
rect 9657 13694 9684 13701
rect 9574 13645 9598 13694
rect 9657 13645 9664 13694
rect 9740 13645 9767 13701
rect 9823 13694 13040 13701
rect 9823 13645 10152 13694
rect 7500 13642 7936 13645
rect 7988 13642 8002 13645
rect 8054 13642 8490 13645
rect 8542 13642 8556 13645
rect 8608 13642 9044 13645
rect 9096 13642 9110 13645
rect 9162 13642 9598 13645
rect 9650 13642 9664 13645
rect 9716 13642 10152 13645
rect 10204 13642 10218 13694
rect 10270 13642 10706 13694
rect 10758 13642 10772 13694
rect 10824 13642 11260 13694
rect 11312 13642 11326 13694
rect 11378 13642 11814 13694
rect 11866 13642 11880 13694
rect 11932 13642 12368 13694
rect 12420 13642 12434 13694
rect 12486 13642 12922 13694
rect 12974 13642 12988 13694
rect 2950 13628 13040 13642
rect 3002 13576 3016 13628
rect 3068 13576 3504 13628
rect 3556 13576 3570 13628
rect 3622 13576 4058 13628
rect 4110 13576 4124 13628
rect 4176 13576 4612 13628
rect 4664 13576 4678 13628
rect 4730 13576 5166 13628
rect 5218 13576 5232 13628
rect 5284 13576 5720 13628
rect 5772 13576 5786 13628
rect 5838 13576 6274 13628
rect 6326 13576 6340 13628
rect 6392 13576 6828 13628
rect 6880 13576 6894 13628
rect 6946 13576 7382 13628
rect 7434 13576 7448 13628
rect 7500 13613 7936 13628
rect 7988 13613 8002 13628
rect 8054 13613 8490 13628
rect 8542 13613 8556 13628
rect 8608 13613 9044 13628
rect 9096 13613 9110 13628
rect 9162 13613 9598 13628
rect 9650 13613 9664 13628
rect 9716 13613 10152 13628
rect 7500 13576 7691 13613
rect 2950 13562 7691 13576
rect 3002 13510 3016 13562
rect 3068 13510 3504 13562
rect 3556 13510 3570 13562
rect 3622 13510 4058 13562
rect 4110 13510 4124 13562
rect 4176 13510 4612 13562
rect 4664 13510 4678 13562
rect 4730 13510 5166 13562
rect 5218 13510 5232 13562
rect 5284 13510 5720 13562
rect 5772 13510 5786 13562
rect 5838 13510 6274 13562
rect 6326 13510 6340 13562
rect 6392 13510 6828 13562
rect 6880 13510 6894 13562
rect 6946 13510 7382 13562
rect 7434 13510 7448 13562
rect 7500 13557 7691 13562
rect 7747 13557 7775 13613
rect 7831 13557 7858 13613
rect 7914 13576 7936 13613
rect 7997 13576 8002 13613
rect 7914 13562 7941 13576
rect 7997 13562 8024 13576
rect 7914 13557 7936 13562
rect 7997 13557 8002 13562
rect 8080 13557 8107 13613
rect 8163 13557 8190 13613
rect 8246 13557 8273 13613
rect 8329 13557 8356 13613
rect 8412 13557 8439 13613
rect 8495 13562 8522 13576
rect 8578 13562 8605 13576
rect 8661 13557 8688 13613
rect 8744 13557 8771 13613
rect 8827 13557 8854 13613
rect 8910 13557 8937 13613
rect 8993 13557 9020 13613
rect 9096 13576 9103 13613
rect 9162 13576 9186 13613
rect 9076 13562 9103 13576
rect 9159 13562 9186 13576
rect 9096 13557 9103 13562
rect 9162 13557 9186 13562
rect 9242 13557 9269 13613
rect 9325 13557 9352 13613
rect 9408 13557 9435 13613
rect 9491 13557 9518 13613
rect 9574 13576 9598 13613
rect 9657 13576 9664 13613
rect 9574 13562 9601 13576
rect 9657 13562 9684 13576
rect 9574 13557 9598 13562
rect 9657 13557 9664 13562
rect 9740 13557 9767 13613
rect 9823 13576 10152 13613
rect 10204 13576 10218 13628
rect 10270 13576 10706 13628
rect 10758 13576 10772 13628
rect 10824 13576 11260 13628
rect 11312 13576 11326 13628
rect 11378 13576 11814 13628
rect 11866 13576 11880 13628
rect 11932 13576 12368 13628
rect 12420 13576 12434 13628
rect 12486 13576 12922 13628
rect 12974 13576 12988 13628
rect 9823 13562 13040 13576
rect 9823 13557 10152 13562
rect 7500 13525 7936 13557
rect 7988 13525 8002 13557
rect 8054 13525 8490 13557
rect 8542 13525 8556 13557
rect 8608 13525 9044 13557
rect 9096 13525 9110 13557
rect 9162 13525 9598 13557
rect 9650 13525 9664 13557
rect 9716 13525 10152 13557
rect 7500 13510 7691 13525
rect 2950 13495 7691 13510
rect 3002 13443 3016 13495
rect 3068 13443 3504 13495
rect 3556 13443 3570 13495
rect 3622 13443 4058 13495
rect 4110 13443 4124 13495
rect 4176 13443 4612 13495
rect 4664 13443 4678 13495
rect 4730 13443 5166 13495
rect 5218 13443 5232 13495
rect 5284 13443 5720 13495
rect 5772 13443 5786 13495
rect 5838 13443 6274 13495
rect 6326 13443 6340 13495
rect 6392 13443 6828 13495
rect 6880 13443 6894 13495
rect 6946 13443 7382 13495
rect 7434 13443 7448 13495
rect 7500 13469 7691 13495
rect 7747 13469 7775 13525
rect 7831 13469 7858 13525
rect 7914 13510 7936 13525
rect 7997 13510 8002 13525
rect 7914 13495 7941 13510
rect 7997 13495 8024 13510
rect 7914 13469 7936 13495
rect 7997 13469 8002 13495
rect 8080 13469 8107 13525
rect 8163 13469 8190 13525
rect 8246 13469 8273 13525
rect 8329 13469 8356 13525
rect 8412 13469 8439 13525
rect 8495 13495 8522 13510
rect 8578 13495 8605 13510
rect 8661 13469 8688 13525
rect 8744 13469 8771 13525
rect 8827 13469 8854 13525
rect 8910 13469 8937 13525
rect 8993 13469 9020 13525
rect 9096 13510 9103 13525
rect 9162 13510 9186 13525
rect 9076 13495 9103 13510
rect 9159 13495 9186 13510
rect 9096 13469 9103 13495
rect 9162 13469 9186 13495
rect 9242 13469 9269 13525
rect 9325 13469 9352 13525
rect 9408 13469 9435 13525
rect 9491 13469 9518 13525
rect 9574 13510 9598 13525
rect 9657 13510 9664 13525
rect 9574 13495 9601 13510
rect 9657 13495 9684 13510
rect 9574 13469 9598 13495
rect 9657 13469 9664 13495
rect 9740 13469 9767 13525
rect 9823 13510 10152 13525
rect 10204 13510 10218 13562
rect 10270 13510 10706 13562
rect 10758 13510 10772 13562
rect 10824 13510 11260 13562
rect 11312 13510 11326 13562
rect 11378 13510 11814 13562
rect 11866 13510 11880 13562
rect 11932 13510 12368 13562
rect 12420 13510 12434 13562
rect 12486 13510 12922 13562
rect 12974 13510 12988 13562
rect 9823 13495 13040 13510
rect 9823 13469 10152 13495
rect 7500 13443 7936 13469
rect 7988 13443 8002 13469
rect 8054 13443 8490 13469
rect 8542 13443 8556 13469
rect 8608 13443 9044 13469
rect 9096 13443 9110 13469
rect 9162 13443 9598 13469
rect 9650 13443 9664 13469
rect 9716 13443 10152 13469
rect 10204 13443 10218 13495
rect 10270 13443 10706 13495
rect 10758 13443 10772 13495
rect 10824 13443 11260 13495
rect 11312 13443 11326 13495
rect 11378 13443 11814 13495
rect 11866 13443 11880 13495
rect 11932 13443 12368 13495
rect 12420 13443 12434 13495
rect 12486 13443 12922 13495
rect 12974 13443 12988 13495
rect 2950 13437 13040 13443
rect 2950 13428 7691 13437
rect 3002 13376 3016 13428
rect 3068 13376 3504 13428
rect 3556 13376 3570 13428
rect 3622 13376 4058 13428
rect 4110 13376 4124 13428
rect 4176 13376 4612 13428
rect 4664 13376 4678 13428
rect 4730 13376 5166 13428
rect 5218 13376 5232 13428
rect 5284 13376 5720 13428
rect 5772 13376 5786 13428
rect 5838 13376 6274 13428
rect 6326 13376 6340 13428
rect 6392 13376 6828 13428
rect 6880 13376 6894 13428
rect 6946 13376 7382 13428
rect 7434 13376 7448 13428
rect 7500 13381 7691 13428
rect 7747 13381 7775 13437
rect 7831 13381 7858 13437
rect 7914 13428 7941 13437
rect 7997 13428 8024 13437
rect 7914 13381 7936 13428
rect 7997 13381 8002 13428
rect 8080 13381 8107 13437
rect 8163 13381 8190 13437
rect 8246 13381 8273 13437
rect 8329 13381 8356 13437
rect 8412 13381 8439 13437
rect 8495 13428 8522 13437
rect 8578 13428 8605 13437
rect 8661 13381 8688 13437
rect 8744 13381 8771 13437
rect 8827 13381 8854 13437
rect 8910 13381 8937 13437
rect 8993 13381 9020 13437
rect 9076 13428 9103 13437
rect 9159 13428 9186 13437
rect 9096 13381 9103 13428
rect 9162 13381 9186 13428
rect 9242 13381 9269 13437
rect 9325 13381 9352 13437
rect 9408 13381 9435 13437
rect 9491 13381 9518 13437
rect 9574 13428 9601 13437
rect 9657 13428 9684 13437
rect 9574 13381 9598 13428
rect 9657 13381 9664 13428
rect 9740 13381 9767 13437
rect 9823 13428 13040 13437
rect 9823 13381 10152 13428
rect 7500 13376 7936 13381
rect 7988 13376 8002 13381
rect 8054 13376 8490 13381
rect 8542 13376 8556 13381
rect 8608 13376 9044 13381
rect 9096 13376 9110 13381
rect 9162 13376 9598 13381
rect 9650 13376 9664 13381
rect 9716 13376 10152 13381
rect 10204 13376 10218 13428
rect 10270 13376 10706 13428
rect 10758 13376 10772 13428
rect 10824 13376 11260 13428
rect 11312 13376 11326 13428
rect 11378 13376 11814 13428
rect 11866 13376 11880 13428
rect 11932 13376 12368 13428
rect 12420 13376 12434 13428
rect 12486 13376 12922 13428
rect 12974 13376 12988 13428
rect 2950 13368 13040 13376
rect 13199 13894 13200 13946
rect 13252 13894 13270 13946
rect 13322 13894 13340 13946
rect 13392 13894 13410 13946
rect 13462 13894 13480 13946
rect 13532 13894 13550 13946
rect 13602 13894 14940 13946
rect 13199 13882 14940 13894
rect 13199 13830 13200 13882
rect 13252 13830 13270 13882
rect 13322 13830 13340 13882
rect 13392 13830 13410 13882
rect 13462 13830 13480 13882
rect 13532 13830 13550 13882
rect 13602 13830 14940 13882
rect 13199 13818 14940 13830
rect 13199 13766 13200 13818
rect 13252 13766 13270 13818
rect 13322 13766 13340 13818
rect 13392 13766 13410 13818
rect 13462 13766 13480 13818
rect 13532 13766 13550 13818
rect 13602 13766 14940 13818
rect 13199 13754 14940 13766
rect 13199 13702 13200 13754
rect 13252 13702 13270 13754
rect 13322 13702 13340 13754
rect 13392 13702 13410 13754
rect 13462 13702 13480 13754
rect 13532 13702 13550 13754
rect 13602 13702 14940 13754
rect 13199 13690 14940 13702
rect 13199 13638 13200 13690
rect 13252 13638 13270 13690
rect 13322 13638 13340 13690
rect 13392 13638 13410 13690
rect 13462 13638 13480 13690
rect 13532 13638 13550 13690
rect 13602 13638 14940 13690
rect 13199 13626 14940 13638
rect 13199 13574 13200 13626
rect 13252 13574 13270 13626
rect 13322 13574 13340 13626
rect 13392 13574 13410 13626
rect 13462 13574 13480 13626
rect 13532 13574 13550 13626
rect 13602 13574 14940 13626
rect 13199 13562 14940 13574
rect 13199 13510 13200 13562
rect 13252 13510 13270 13562
rect 13322 13510 13340 13562
rect 13392 13510 13410 13562
rect 13462 13510 13480 13562
rect 13532 13510 13550 13562
rect 13602 13510 14940 13562
rect 13199 13498 14940 13510
rect 13199 13446 13200 13498
rect 13252 13446 13270 13498
rect 13322 13446 13340 13498
rect 13392 13446 13410 13498
rect 13462 13446 13480 13498
rect 13532 13446 13550 13498
rect 13602 13446 14940 13498
rect 13199 13434 14940 13446
rect 13199 13382 13200 13434
rect 13252 13382 13270 13434
rect 13322 13382 13340 13434
rect 13392 13382 13410 13434
rect 13462 13382 13480 13434
rect 13532 13382 13550 13434
rect 13602 13382 14940 13434
rect 13199 13370 14940 13382
rect 13199 13318 13200 13370
rect 13252 13318 13270 13370
rect 13322 13318 13340 13370
rect 13392 13318 13410 13370
rect 13462 13318 13480 13370
rect 13532 13318 13550 13370
rect 13602 13318 14940 13370
rect 13199 13306 14940 13318
rect 13199 13254 13200 13306
rect 13252 13254 13270 13306
rect 13322 13254 13340 13306
rect 13392 13254 13410 13306
rect 13462 13254 13480 13306
rect 13532 13254 13550 13306
rect 13602 13254 14940 13306
rect 13199 13242 14940 13254
rect 13199 13190 13200 13242
rect 13252 13190 13270 13242
rect 13322 13190 13340 13242
rect 13392 13190 13410 13242
rect 13462 13190 13480 13242
rect 13532 13190 13550 13242
rect 13602 13190 14940 13242
rect 13199 13178 14940 13190
rect 13199 13126 13200 13178
rect 13252 13126 13270 13178
rect 13322 13126 13340 13178
rect 13392 13126 13410 13178
rect 13462 13126 13480 13178
rect 13532 13126 13550 13178
rect 13602 13126 14940 13178
rect 13199 13114 14940 13126
rect 13199 13062 13200 13114
rect 13252 13062 13270 13114
rect 13322 13062 13340 13114
rect 13392 13062 13410 13114
rect 13462 13062 13480 13114
rect 13532 13062 13550 13114
rect 13602 13062 14940 13114
rect 13199 13050 14940 13062
rect 13199 12998 13200 13050
rect 13252 12998 13270 13050
rect 13322 12998 13340 13050
rect 13392 12998 13410 13050
rect 13462 12998 13480 13050
rect 13532 12998 13550 13050
rect 13602 12998 14940 13050
rect 13199 12986 14940 12998
tri 13197 12934 13199 12936 se
rect 13199 12934 13200 12986
rect 13252 12934 13270 12986
rect 13322 12934 13340 12986
rect 13392 12934 13410 12986
rect 13462 12934 13480 12986
rect 13532 12934 13550 12986
rect 13602 12934 14940 12986
tri 13185 12922 13197 12934 se
rect 13197 12922 14940 12934
tri 13133 12870 13185 12922 se
rect 13185 12870 13200 12922
rect 13252 12870 13270 12922
rect 13322 12870 13340 12922
rect 13392 12870 13410 12922
rect 13462 12870 13480 12922
rect 13532 12870 13550 12922
rect 13602 12870 14940 12922
tri 13121 12858 13133 12870 se
rect 13133 12858 14940 12870
tri 13069 12806 13121 12858 se
rect 13121 12806 13200 12858
rect 13252 12806 13270 12858
rect 13322 12806 13340 12858
rect 13392 12806 13410 12858
rect 13462 12806 13480 12858
rect 13532 12806 13550 12858
rect 13602 12806 14940 12858
tri 13057 12794 13069 12806 se
rect 13069 12794 14940 12806
tri 13005 12742 13057 12794 se
rect 13057 12742 13200 12794
rect 13252 12742 13270 12794
rect 13322 12742 13340 12794
rect 13392 12742 13410 12794
rect 13462 12742 13480 12794
rect 13532 12742 13550 12794
rect 13602 12742 14940 12794
tri 12993 12730 13005 12742 se
rect 13005 12730 14940 12742
tri 12989 12726 12993 12730 se
rect 12993 12726 13200 12730
rect 3227 12720 13200 12726
rect 3279 12668 3293 12720
rect 3345 12668 3781 12720
rect 3833 12668 3847 12720
rect 3899 12668 4335 12720
rect 4387 12668 4401 12720
rect 4453 12668 4889 12720
rect 4941 12668 4955 12720
rect 5007 12668 5443 12720
rect 5495 12668 5509 12720
rect 5561 12668 5997 12720
rect 6049 12668 6063 12720
rect 6115 12668 6551 12720
rect 6603 12668 6617 12720
rect 6669 12668 7105 12720
rect 7157 12668 7171 12720
rect 7223 12668 7659 12720
rect 7711 12668 7725 12720
rect 7777 12668 8213 12720
rect 8265 12668 8279 12720
rect 8331 12668 8767 12720
rect 8819 12668 8833 12720
rect 8885 12668 9321 12720
rect 9373 12668 9387 12720
rect 9439 12668 9875 12720
rect 9927 12668 9941 12720
rect 9993 12668 10429 12720
rect 10481 12668 10495 12720
rect 10547 12668 10983 12720
rect 11035 12668 11049 12720
rect 11101 12668 11537 12720
rect 11589 12668 11603 12720
rect 11655 12668 12091 12720
rect 12143 12668 12157 12720
rect 12209 12668 12645 12720
rect 12697 12668 12711 12720
rect 12763 12678 13200 12720
rect 13252 12678 13270 12730
rect 13322 12678 13340 12730
rect 13392 12678 13410 12730
rect 13462 12678 13480 12730
rect 13532 12678 13550 12730
rect 13602 12678 14940 12730
rect 12763 12668 14940 12678
rect 3227 12666 14940 12668
rect 3227 12654 13200 12666
rect 3279 12602 3293 12654
rect 3345 12602 3781 12654
rect 3833 12602 3847 12654
rect 3899 12602 4335 12654
rect 4387 12602 4401 12654
rect 4453 12602 4889 12654
rect 4941 12602 4955 12654
rect 5007 12602 5443 12654
rect 5495 12602 5509 12654
rect 5561 12602 5997 12654
rect 6049 12602 6063 12654
rect 6115 12602 6551 12654
rect 6603 12602 6617 12654
rect 6669 12602 7105 12654
rect 7157 12602 7171 12654
rect 7223 12602 7659 12654
rect 7711 12602 7725 12654
rect 7777 12602 8213 12654
rect 8265 12602 8279 12654
rect 8331 12602 8767 12654
rect 8819 12602 8833 12654
rect 8885 12602 9321 12654
rect 9373 12602 9387 12654
rect 9439 12602 9875 12654
rect 9927 12602 9941 12654
rect 9993 12602 10429 12654
rect 10481 12602 10495 12654
rect 10547 12602 10983 12654
rect 11035 12602 11049 12654
rect 11101 12602 11537 12654
rect 11589 12602 11603 12654
rect 11655 12602 12091 12654
rect 12143 12602 12157 12654
rect 12209 12602 12645 12654
rect 12697 12602 12711 12654
rect 12763 12614 13200 12654
rect 13252 12614 13270 12666
rect 13322 12614 13340 12666
rect 13392 12614 13410 12666
rect 13462 12614 13480 12666
rect 13532 12614 13550 12666
rect 13602 12614 14940 12666
rect 12763 12602 14940 12614
rect 3227 12588 13200 12602
rect 3279 12536 3293 12588
rect 3345 12536 3781 12588
rect 3833 12536 3847 12588
rect 3899 12536 4335 12588
rect 4387 12536 4401 12588
rect 4453 12536 4889 12588
rect 4941 12536 4955 12588
rect 5007 12536 5443 12588
rect 5495 12536 5509 12588
rect 5561 12536 5997 12588
rect 6049 12536 6063 12588
rect 6115 12536 6551 12588
rect 6603 12536 6617 12588
rect 6669 12536 7105 12588
rect 7157 12536 7171 12588
rect 7223 12536 7659 12588
rect 7711 12536 7725 12588
rect 7777 12536 8213 12588
rect 8265 12536 8279 12588
rect 8331 12536 8767 12588
rect 8819 12536 8833 12588
rect 8885 12536 9321 12588
rect 9373 12536 9387 12588
rect 9439 12536 9875 12588
rect 9927 12536 9941 12588
rect 9993 12536 10429 12588
rect 10481 12536 10495 12588
rect 10547 12536 10983 12588
rect 11035 12536 11049 12588
rect 11101 12536 11537 12588
rect 11589 12536 11603 12588
rect 11655 12536 12091 12588
rect 12143 12536 12157 12588
rect 12209 12536 12645 12588
rect 12697 12536 12711 12588
rect 12763 12550 13200 12588
rect 13252 12550 13270 12602
rect 13322 12550 13340 12602
rect 13392 12550 13410 12602
rect 13462 12550 13480 12602
rect 13532 12550 13550 12602
rect 13602 12550 14940 12602
rect 12763 12538 14940 12550
rect 12763 12536 13200 12538
rect 3227 12522 13200 12536
rect 3279 12470 3293 12522
rect 3345 12470 3781 12522
rect 3833 12470 3847 12522
rect 3899 12470 4335 12522
rect 4387 12470 4401 12522
rect 4453 12470 4889 12522
rect 4941 12470 4955 12522
rect 5007 12470 5443 12522
rect 5495 12470 5509 12522
rect 5561 12470 5997 12522
rect 6049 12470 6063 12522
rect 6115 12470 6551 12522
rect 6603 12470 6617 12522
rect 6669 12470 7105 12522
rect 7157 12470 7171 12522
rect 7223 12470 7659 12522
rect 7711 12470 7725 12522
rect 7777 12470 8213 12522
rect 8265 12470 8279 12522
rect 8331 12470 8767 12522
rect 8819 12470 8833 12522
rect 8885 12470 9321 12522
rect 9373 12470 9387 12522
rect 9439 12470 9875 12522
rect 9927 12470 9941 12522
rect 9993 12470 10429 12522
rect 10481 12470 10495 12522
rect 10547 12470 10983 12522
rect 11035 12470 11049 12522
rect 11101 12470 11537 12522
rect 11589 12470 11603 12522
rect 11655 12470 12091 12522
rect 12143 12470 12157 12522
rect 12209 12470 12645 12522
rect 12697 12470 12711 12522
rect 12763 12486 13200 12522
rect 13252 12486 13270 12538
rect 13322 12486 13340 12538
rect 13392 12486 13410 12538
rect 13462 12486 13480 12538
rect 13532 12486 13550 12538
rect 13602 12486 14940 12538
rect 12763 12474 14940 12486
rect 12763 12470 13200 12474
rect 3227 12456 13200 12470
rect 3279 12404 3293 12456
rect 3345 12404 3781 12456
rect 3833 12404 3847 12456
rect 3899 12404 4335 12456
rect 4387 12404 4401 12456
rect 4453 12404 4889 12456
rect 4941 12404 4955 12456
rect 5007 12404 5443 12456
rect 5495 12404 5509 12456
rect 5561 12404 5997 12456
rect 6049 12404 6063 12456
rect 6115 12404 6551 12456
rect 6603 12404 6617 12456
rect 6669 12404 7105 12456
rect 7157 12404 7171 12456
rect 7223 12404 7659 12456
rect 7711 12404 7725 12456
rect 7777 12404 8213 12456
rect 8265 12404 8279 12456
rect 8331 12404 8767 12456
rect 8819 12404 8833 12456
rect 8885 12404 9321 12456
rect 9373 12404 9387 12456
rect 9439 12404 9875 12456
rect 9927 12404 9941 12456
rect 9993 12404 10429 12456
rect 10481 12404 10495 12456
rect 10547 12404 10983 12456
rect 11035 12404 11049 12456
rect 11101 12404 11537 12456
rect 11589 12404 11603 12456
rect 11655 12404 12091 12456
rect 12143 12404 12157 12456
rect 12209 12404 12645 12456
rect 12697 12404 12711 12456
rect 12763 12422 13200 12456
rect 13252 12422 13270 12474
rect 13322 12422 13340 12474
rect 13392 12422 13410 12474
rect 13462 12422 13480 12474
rect 13532 12422 13550 12474
rect 13602 12422 14940 12474
rect 12763 12410 14940 12422
rect 12763 12404 13200 12410
rect 3227 12390 13200 12404
rect 3279 12338 3293 12390
rect 3345 12338 3781 12390
rect 3833 12338 3847 12390
rect 3899 12338 4335 12390
rect 4387 12338 4401 12390
rect 4453 12338 4889 12390
rect 4941 12338 4955 12390
rect 5007 12338 5443 12390
rect 5495 12338 5509 12390
rect 5561 12338 5997 12390
rect 6049 12338 6063 12390
rect 6115 12338 6551 12390
rect 6603 12338 6617 12390
rect 6669 12338 7105 12390
rect 7157 12338 7171 12390
rect 7223 12338 7659 12390
rect 7711 12338 7725 12390
rect 7777 12338 8213 12390
rect 8265 12338 8279 12390
rect 8331 12338 8767 12390
rect 8819 12338 8833 12390
rect 8885 12338 9321 12390
rect 9373 12338 9387 12390
rect 9439 12338 9875 12390
rect 9927 12338 9941 12390
rect 9993 12338 10429 12390
rect 10481 12338 10495 12390
rect 10547 12338 10983 12390
rect 11035 12338 11049 12390
rect 11101 12338 11537 12390
rect 11589 12338 11603 12390
rect 11655 12338 12091 12390
rect 12143 12338 12157 12390
rect 12209 12338 12645 12390
rect 12697 12338 12711 12390
rect 12763 12358 13200 12390
rect 13252 12358 13270 12410
rect 13322 12358 13340 12410
rect 13392 12358 13410 12410
rect 13462 12358 13480 12410
rect 13532 12358 13550 12410
rect 13602 12358 14940 12410
rect 12763 12346 14940 12358
rect 12763 12338 13200 12346
rect 3227 12323 13200 12338
rect 3279 12271 3293 12323
rect 3345 12271 3781 12323
rect 3833 12271 3847 12323
rect 3899 12271 4335 12323
rect 4387 12271 4401 12323
rect 4453 12271 4889 12323
rect 4941 12271 4955 12323
rect 5007 12271 5443 12323
rect 5495 12271 5509 12323
rect 5561 12271 5997 12323
rect 6049 12271 6063 12323
rect 6115 12271 6551 12323
rect 6603 12271 6617 12323
rect 6669 12271 7105 12323
rect 7157 12271 7171 12323
rect 7223 12271 7659 12323
rect 7711 12271 7725 12323
rect 7777 12271 8213 12323
rect 8265 12271 8279 12323
rect 8331 12271 8767 12323
rect 8819 12271 8833 12323
rect 8885 12271 9321 12323
rect 9373 12271 9387 12323
rect 9439 12271 9875 12323
rect 9927 12271 9941 12323
rect 9993 12271 10429 12323
rect 10481 12271 10495 12323
rect 10547 12271 10983 12323
rect 11035 12271 11049 12323
rect 11101 12271 11537 12323
rect 11589 12271 11603 12323
rect 11655 12271 12091 12323
rect 12143 12271 12157 12323
rect 12209 12271 12645 12323
rect 12697 12271 12711 12323
rect 12763 12294 13200 12323
rect 13252 12294 13270 12346
rect 13322 12294 13340 12346
rect 13392 12294 13410 12346
rect 13462 12294 13480 12346
rect 13532 12294 13550 12346
rect 13602 12294 14940 12346
rect 12763 12282 14940 12294
rect 12763 12271 13200 12282
rect 3227 12256 13200 12271
rect 3279 12204 3293 12256
rect 3345 12204 3781 12256
rect 3833 12204 3847 12256
rect 3899 12204 4335 12256
rect 4387 12204 4401 12256
rect 4453 12204 4889 12256
rect 4941 12204 4955 12256
rect 5007 12204 5443 12256
rect 5495 12204 5509 12256
rect 5561 12204 5997 12256
rect 6049 12204 6063 12256
rect 6115 12204 6551 12256
rect 6603 12204 6617 12256
rect 6669 12204 7105 12256
rect 7157 12204 7171 12256
rect 7223 12204 7659 12256
rect 7711 12204 7725 12256
rect 7777 12204 8213 12256
rect 8265 12204 8279 12256
rect 8331 12204 8767 12256
rect 8819 12204 8833 12256
rect 8885 12204 9321 12256
rect 9373 12204 9387 12256
rect 9439 12204 9875 12256
rect 9927 12204 9941 12256
rect 9993 12204 10429 12256
rect 10481 12204 10495 12256
rect 10547 12204 10983 12256
rect 11035 12204 11049 12256
rect 11101 12204 11537 12256
rect 11589 12204 11603 12256
rect 11655 12204 12091 12256
rect 12143 12204 12157 12256
rect 12209 12204 12645 12256
rect 12697 12204 12711 12256
rect 12763 12230 13200 12256
rect 13252 12230 13270 12282
rect 13322 12230 13340 12282
rect 13392 12230 13410 12282
rect 13462 12230 13480 12282
rect 13532 12230 13550 12282
rect 13602 12230 14940 12282
rect 12763 12218 14940 12230
rect 12763 12204 13200 12218
rect 3227 12198 13200 12204
tri 12989 12166 13021 12198 ne
rect 13021 12166 13200 12198
rect 13252 12166 13270 12218
rect 13322 12166 13340 12218
rect 13392 12166 13410 12218
rect 13462 12166 13480 12218
rect 13532 12166 13550 12218
rect 13602 12166 14940 12218
tri 13021 12154 13033 12166 ne
rect 13033 12154 14940 12166
tri 13033 12102 13085 12154 ne
rect 13085 12102 13200 12154
rect 13252 12102 13270 12154
rect 13322 12102 13340 12154
rect 13392 12102 13410 12154
rect 13462 12102 13480 12154
rect 13532 12102 13550 12154
rect 13602 12102 14940 12154
tri 13085 12090 13097 12102 ne
rect 13097 12090 14940 12102
tri 13097 12038 13149 12090 ne
rect 13149 12038 13200 12090
rect 13252 12038 13270 12090
rect 13322 12038 13340 12090
rect 13392 12038 13410 12090
rect 13462 12038 13480 12090
rect 13532 12038 13550 12090
rect 13602 12038 14940 12090
tri 13149 12026 13161 12038 ne
rect 13161 12026 14940 12038
tri 13161 11988 13199 12026 ne
rect 13199 11974 13200 12026
rect 13252 11974 13270 12026
rect 13322 11974 13340 12026
rect 13392 11974 13410 12026
rect 13462 11974 13480 12026
rect 13532 11974 13550 12026
rect 13602 11974 14940 12026
rect 13199 11962 14940 11974
rect 13199 11910 13200 11962
rect 13252 11910 13270 11962
rect 13322 11910 13340 11962
rect 13392 11910 13410 11962
rect 13462 11910 13480 11962
rect 13532 11910 13550 11962
rect 13602 11910 14940 11962
rect 13199 11898 14940 11910
rect 2950 11892 13040 11898
rect 3002 11840 3016 11892
rect 3068 11840 3504 11892
rect 3556 11840 3570 11892
rect 3622 11840 4058 11892
rect 4110 11840 4124 11892
rect 4176 11840 4612 11892
rect 4664 11840 4678 11892
rect 4730 11840 5166 11892
rect 5218 11840 5232 11892
rect 5284 11840 5720 11892
rect 5772 11840 5786 11892
rect 5838 11840 6274 11892
rect 6326 11840 6340 11892
rect 6392 11840 6828 11892
rect 6880 11840 6894 11892
rect 6946 11840 7382 11892
rect 7434 11840 7448 11892
rect 7500 11882 7936 11892
rect 7988 11882 8002 11892
rect 8054 11882 8490 11892
rect 8542 11882 8556 11892
rect 8608 11882 9044 11892
rect 9096 11882 9110 11892
rect 9162 11882 9598 11892
rect 9650 11882 9664 11892
rect 9716 11882 10152 11892
rect 7500 11840 7691 11882
rect 2950 11826 7691 11840
rect 7747 11826 7775 11882
rect 7831 11826 7858 11882
rect 7914 11840 7936 11882
rect 7997 11840 8002 11882
rect 7914 11826 7941 11840
rect 7997 11826 8024 11840
rect 8080 11826 8107 11882
rect 8163 11826 8190 11882
rect 8246 11826 8273 11882
rect 8329 11826 8356 11882
rect 8412 11826 8439 11882
rect 8495 11826 8522 11840
rect 8578 11826 8605 11840
rect 8661 11826 8688 11882
rect 8744 11826 8771 11882
rect 8827 11826 8854 11882
rect 8910 11826 8937 11882
rect 8993 11826 9020 11882
rect 9096 11840 9103 11882
rect 9162 11840 9186 11882
rect 9076 11826 9103 11840
rect 9159 11826 9186 11840
rect 9242 11826 9269 11882
rect 9325 11826 9352 11882
rect 9408 11826 9435 11882
rect 9491 11826 9518 11882
rect 9574 11840 9598 11882
rect 9657 11840 9664 11882
rect 9574 11826 9601 11840
rect 9657 11826 9684 11840
rect 9740 11826 9767 11882
rect 9823 11840 10152 11882
rect 10204 11840 10218 11892
rect 10270 11840 10706 11892
rect 10758 11840 10772 11892
rect 10824 11840 11260 11892
rect 11312 11840 11326 11892
rect 11378 11840 11814 11892
rect 11866 11840 11880 11892
rect 11932 11840 12368 11892
rect 12420 11840 12434 11892
rect 12486 11840 12922 11892
rect 12974 11840 12988 11892
rect 9823 11826 13040 11840
rect 3002 11774 3016 11826
rect 3068 11774 3504 11826
rect 3556 11774 3570 11826
rect 3622 11774 4058 11826
rect 4110 11774 4124 11826
rect 4176 11774 4612 11826
rect 4664 11774 4678 11826
rect 4730 11774 5166 11826
rect 5218 11774 5232 11826
rect 5284 11774 5720 11826
rect 5772 11774 5786 11826
rect 5838 11774 6274 11826
rect 6326 11774 6340 11826
rect 6392 11774 6828 11826
rect 6880 11774 6894 11826
rect 6946 11774 7382 11826
rect 7434 11774 7448 11826
rect 7500 11794 7936 11826
rect 7988 11794 8002 11826
rect 8054 11794 8490 11826
rect 8542 11794 8556 11826
rect 8608 11794 9044 11826
rect 9096 11794 9110 11826
rect 9162 11794 9598 11826
rect 9650 11794 9664 11826
rect 9716 11794 10152 11826
rect 7500 11774 7691 11794
rect 2950 11760 7691 11774
rect 3002 11708 3016 11760
rect 3068 11708 3504 11760
rect 3556 11708 3570 11760
rect 3622 11708 4058 11760
rect 4110 11708 4124 11760
rect 4176 11708 4612 11760
rect 4664 11708 4678 11760
rect 4730 11708 5166 11760
rect 5218 11708 5232 11760
rect 5284 11708 5720 11760
rect 5772 11708 5786 11760
rect 5838 11708 6274 11760
rect 6326 11708 6340 11760
rect 6392 11708 6828 11760
rect 6880 11708 6894 11760
rect 6946 11708 7382 11760
rect 7434 11708 7448 11760
rect 7500 11738 7691 11760
rect 7747 11738 7775 11794
rect 7831 11738 7858 11794
rect 7914 11774 7936 11794
rect 7997 11774 8002 11794
rect 7914 11760 7941 11774
rect 7997 11760 8024 11774
rect 7914 11738 7936 11760
rect 7997 11738 8002 11760
rect 8080 11738 8107 11794
rect 8163 11738 8190 11794
rect 8246 11738 8273 11794
rect 8329 11738 8356 11794
rect 8412 11738 8439 11794
rect 8495 11760 8522 11774
rect 8578 11760 8605 11774
rect 8661 11738 8688 11794
rect 8744 11738 8771 11794
rect 8827 11738 8854 11794
rect 8910 11738 8937 11794
rect 8993 11738 9020 11794
rect 9096 11774 9103 11794
rect 9162 11774 9186 11794
rect 9076 11760 9103 11774
rect 9159 11760 9186 11774
rect 9096 11738 9103 11760
rect 9162 11738 9186 11760
rect 9242 11738 9269 11794
rect 9325 11738 9352 11794
rect 9408 11738 9435 11794
rect 9491 11738 9518 11794
rect 9574 11774 9598 11794
rect 9657 11774 9664 11794
rect 9574 11760 9601 11774
rect 9657 11760 9684 11774
rect 9574 11738 9598 11760
rect 9657 11738 9664 11760
rect 9740 11738 9767 11794
rect 9823 11774 10152 11794
rect 10204 11774 10218 11826
rect 10270 11774 10706 11826
rect 10758 11774 10772 11826
rect 10824 11774 11260 11826
rect 11312 11774 11326 11826
rect 11378 11774 11814 11826
rect 11866 11774 11880 11826
rect 11932 11774 12368 11826
rect 12420 11774 12434 11826
rect 12486 11774 12922 11826
rect 12974 11774 12988 11826
rect 9823 11760 13040 11774
rect 9823 11738 10152 11760
rect 7500 11708 7936 11738
rect 7988 11708 8002 11738
rect 8054 11708 8490 11738
rect 8542 11708 8556 11738
rect 8608 11708 9044 11738
rect 9096 11708 9110 11738
rect 9162 11708 9598 11738
rect 9650 11708 9664 11738
rect 9716 11708 10152 11738
rect 10204 11708 10218 11760
rect 10270 11708 10706 11760
rect 10758 11708 10772 11760
rect 10824 11708 11260 11760
rect 11312 11708 11326 11760
rect 11378 11708 11814 11760
rect 11866 11708 11880 11760
rect 11932 11708 12368 11760
rect 12420 11708 12434 11760
rect 12486 11708 12922 11760
rect 12974 11708 12988 11760
rect 2950 11706 13040 11708
rect 2950 11694 7691 11706
rect 3002 11642 3016 11694
rect 3068 11642 3504 11694
rect 3556 11642 3570 11694
rect 3622 11642 4058 11694
rect 4110 11642 4124 11694
rect 4176 11642 4612 11694
rect 4664 11642 4678 11694
rect 4730 11642 5166 11694
rect 5218 11642 5232 11694
rect 5284 11642 5720 11694
rect 5772 11642 5786 11694
rect 5838 11642 6274 11694
rect 6326 11642 6340 11694
rect 6392 11642 6828 11694
rect 6880 11642 6894 11694
rect 6946 11642 7382 11694
rect 7434 11642 7448 11694
rect 7500 11650 7691 11694
rect 7747 11650 7775 11706
rect 7831 11650 7858 11706
rect 7914 11694 7941 11706
rect 7997 11694 8024 11706
rect 7914 11650 7936 11694
rect 7997 11650 8002 11694
rect 8080 11650 8107 11706
rect 8163 11650 8190 11706
rect 8246 11650 8273 11706
rect 8329 11650 8356 11706
rect 8412 11650 8439 11706
rect 8495 11694 8522 11706
rect 8578 11694 8605 11706
rect 8661 11650 8688 11706
rect 8744 11650 8771 11706
rect 8827 11650 8854 11706
rect 8910 11650 8937 11706
rect 8993 11650 9020 11706
rect 9076 11694 9103 11706
rect 9159 11694 9186 11706
rect 9096 11650 9103 11694
rect 9162 11650 9186 11694
rect 9242 11650 9269 11706
rect 9325 11650 9352 11706
rect 9408 11650 9435 11706
rect 9491 11650 9518 11706
rect 9574 11694 9601 11706
rect 9657 11694 9684 11706
rect 9574 11650 9598 11694
rect 9657 11650 9664 11694
rect 9740 11650 9767 11706
rect 9823 11694 13040 11706
rect 9823 11650 10152 11694
rect 7500 11642 7936 11650
rect 7988 11642 8002 11650
rect 8054 11642 8490 11650
rect 8542 11642 8556 11650
rect 8608 11642 9044 11650
rect 9096 11642 9110 11650
rect 9162 11642 9598 11650
rect 9650 11642 9664 11650
rect 9716 11642 10152 11650
rect 10204 11642 10218 11694
rect 10270 11642 10706 11694
rect 10758 11642 10772 11694
rect 10824 11642 11260 11694
rect 11312 11642 11326 11694
rect 11378 11642 11814 11694
rect 11866 11642 11880 11694
rect 11932 11642 12368 11694
rect 12420 11642 12434 11694
rect 12486 11642 12922 11694
rect 12974 11642 12988 11694
rect 2950 11628 13040 11642
rect 3002 11576 3016 11628
rect 3068 11576 3504 11628
rect 3556 11576 3570 11628
rect 3622 11576 4058 11628
rect 4110 11576 4124 11628
rect 4176 11576 4612 11628
rect 4664 11576 4678 11628
rect 4730 11576 5166 11628
rect 5218 11576 5232 11628
rect 5284 11576 5720 11628
rect 5772 11576 5786 11628
rect 5838 11576 6274 11628
rect 6326 11576 6340 11628
rect 6392 11576 6828 11628
rect 6880 11576 6894 11628
rect 6946 11576 7382 11628
rect 7434 11576 7448 11628
rect 7500 11618 7936 11628
rect 7988 11618 8002 11628
rect 8054 11618 8490 11628
rect 8542 11618 8556 11628
rect 8608 11618 9044 11628
rect 9096 11618 9110 11628
rect 9162 11618 9598 11628
rect 9650 11618 9664 11628
rect 9716 11618 10152 11628
rect 7500 11576 7691 11618
rect 2950 11562 7691 11576
rect 7747 11562 7775 11618
rect 7831 11562 7858 11618
rect 7914 11576 7936 11618
rect 7997 11576 8002 11618
rect 7914 11562 7941 11576
rect 7997 11562 8024 11576
rect 8080 11562 8107 11618
rect 8163 11562 8190 11618
rect 8246 11562 8273 11618
rect 8329 11562 8356 11618
rect 8412 11562 8439 11618
rect 8495 11562 8522 11576
rect 8578 11562 8605 11576
rect 8661 11562 8688 11618
rect 8744 11562 8771 11618
rect 8827 11562 8854 11618
rect 8910 11562 8937 11618
rect 8993 11562 9020 11618
rect 9096 11576 9103 11618
rect 9162 11576 9186 11618
rect 9076 11562 9103 11576
rect 9159 11562 9186 11576
rect 9242 11562 9269 11618
rect 9325 11562 9352 11618
rect 9408 11562 9435 11618
rect 9491 11562 9518 11618
rect 9574 11576 9598 11618
rect 9657 11576 9664 11618
rect 9574 11562 9601 11576
rect 9657 11562 9684 11576
rect 9740 11562 9767 11618
rect 9823 11576 10152 11618
rect 10204 11576 10218 11628
rect 10270 11576 10706 11628
rect 10758 11576 10772 11628
rect 10824 11576 11260 11628
rect 11312 11576 11326 11628
rect 11378 11576 11814 11628
rect 11866 11576 11880 11628
rect 11932 11576 12368 11628
rect 12420 11576 12434 11628
rect 12486 11576 12922 11628
rect 12974 11576 12988 11628
rect 9823 11562 13040 11576
rect 3002 11510 3016 11562
rect 3068 11510 3504 11562
rect 3556 11510 3570 11562
rect 3622 11510 4058 11562
rect 4110 11510 4124 11562
rect 4176 11510 4612 11562
rect 4664 11510 4678 11562
rect 4730 11510 5166 11562
rect 5218 11510 5232 11562
rect 5284 11510 5720 11562
rect 5772 11510 5786 11562
rect 5838 11510 6274 11562
rect 6326 11510 6340 11562
rect 6392 11510 6828 11562
rect 6880 11510 6894 11562
rect 6946 11510 7382 11562
rect 7434 11510 7448 11562
rect 7500 11530 7936 11562
rect 7988 11530 8002 11562
rect 8054 11530 8490 11562
rect 8542 11530 8556 11562
rect 8608 11530 9044 11562
rect 9096 11530 9110 11562
rect 9162 11530 9598 11562
rect 9650 11530 9664 11562
rect 9716 11530 10152 11562
rect 7500 11510 7691 11530
rect 2950 11495 7691 11510
rect 3002 11443 3016 11495
rect 3068 11443 3504 11495
rect 3556 11443 3570 11495
rect 3622 11443 4058 11495
rect 4110 11443 4124 11495
rect 4176 11443 4612 11495
rect 4664 11443 4678 11495
rect 4730 11443 5166 11495
rect 5218 11443 5232 11495
rect 5284 11443 5720 11495
rect 5772 11443 5786 11495
rect 5838 11443 6274 11495
rect 6326 11443 6340 11495
rect 6392 11443 6828 11495
rect 6880 11443 6894 11495
rect 6946 11443 7382 11495
rect 7434 11443 7448 11495
rect 7500 11474 7691 11495
rect 7747 11474 7775 11530
rect 7831 11474 7858 11530
rect 7914 11510 7936 11530
rect 7997 11510 8002 11530
rect 7914 11495 7941 11510
rect 7997 11495 8024 11510
rect 7914 11474 7936 11495
rect 7997 11474 8002 11495
rect 8080 11474 8107 11530
rect 8163 11474 8190 11530
rect 8246 11474 8273 11530
rect 8329 11474 8356 11530
rect 8412 11474 8439 11530
rect 8495 11495 8522 11510
rect 8578 11495 8605 11510
rect 8661 11474 8688 11530
rect 8744 11474 8771 11530
rect 8827 11474 8854 11530
rect 8910 11474 8937 11530
rect 8993 11474 9020 11530
rect 9096 11510 9103 11530
rect 9162 11510 9186 11530
rect 9076 11495 9103 11510
rect 9159 11495 9186 11510
rect 9096 11474 9103 11495
rect 9162 11474 9186 11495
rect 9242 11474 9269 11530
rect 9325 11474 9352 11530
rect 9408 11474 9435 11530
rect 9491 11474 9518 11530
rect 9574 11510 9598 11530
rect 9657 11510 9664 11530
rect 9574 11495 9601 11510
rect 9657 11495 9684 11510
rect 9574 11474 9598 11495
rect 9657 11474 9664 11495
rect 9740 11474 9767 11530
rect 9823 11510 10152 11530
rect 10204 11510 10218 11562
rect 10270 11510 10706 11562
rect 10758 11510 10772 11562
rect 10824 11510 11260 11562
rect 11312 11510 11326 11562
rect 11378 11510 11814 11562
rect 11866 11510 11880 11562
rect 11932 11510 12368 11562
rect 12420 11510 12434 11562
rect 12486 11510 12922 11562
rect 12974 11510 12988 11562
rect 9823 11495 13040 11510
rect 9823 11474 10152 11495
rect 7500 11443 7936 11474
rect 7988 11443 8002 11474
rect 8054 11443 8490 11474
rect 8542 11443 8556 11474
rect 8608 11443 9044 11474
rect 9096 11443 9110 11474
rect 9162 11443 9598 11474
rect 9650 11443 9664 11474
rect 9716 11443 10152 11474
rect 10204 11443 10218 11495
rect 10270 11443 10706 11495
rect 10758 11443 10772 11495
rect 10824 11443 11260 11495
rect 11312 11443 11326 11495
rect 11378 11443 11814 11495
rect 11866 11443 11880 11495
rect 11932 11443 12368 11495
rect 12420 11443 12434 11495
rect 12486 11443 12922 11495
rect 12974 11443 12988 11495
rect 2950 11442 13040 11443
rect 2950 11428 7691 11442
rect 3002 11376 3016 11428
rect 3068 11376 3504 11428
rect 3556 11376 3570 11428
rect 3622 11376 4058 11428
rect 4110 11376 4124 11428
rect 4176 11376 4612 11428
rect 4664 11376 4678 11428
rect 4730 11376 5166 11428
rect 5218 11376 5232 11428
rect 5284 11376 5720 11428
rect 5772 11376 5786 11428
rect 5838 11376 6274 11428
rect 6326 11376 6340 11428
rect 6392 11376 6828 11428
rect 6880 11376 6894 11428
rect 6946 11376 7382 11428
rect 7434 11376 7448 11428
rect 7500 11386 7691 11428
rect 7747 11386 7775 11442
rect 7831 11386 7858 11442
rect 7914 11428 7941 11442
rect 7997 11428 8024 11442
rect 7914 11386 7936 11428
rect 7997 11386 8002 11428
rect 8080 11386 8107 11442
rect 8163 11386 8190 11442
rect 8246 11386 8273 11442
rect 8329 11386 8356 11442
rect 8412 11386 8439 11442
rect 8495 11428 8522 11442
rect 8578 11428 8605 11442
rect 8661 11386 8688 11442
rect 8744 11386 8771 11442
rect 8827 11386 8854 11442
rect 8910 11386 8937 11442
rect 8993 11386 9020 11442
rect 9076 11428 9103 11442
rect 9159 11428 9186 11442
rect 9096 11386 9103 11428
rect 9162 11386 9186 11428
rect 9242 11386 9269 11442
rect 9325 11386 9352 11442
rect 9408 11386 9435 11442
rect 9491 11386 9518 11442
rect 9574 11428 9601 11442
rect 9657 11428 9684 11442
rect 9574 11386 9598 11428
rect 9657 11386 9664 11428
rect 9740 11386 9767 11442
rect 9823 11428 13040 11442
rect 9823 11386 10152 11428
rect 7500 11376 7936 11386
rect 7988 11376 8002 11386
rect 8054 11376 8490 11386
rect 8542 11376 8556 11386
rect 8608 11376 9044 11386
rect 9096 11376 9110 11386
rect 9162 11376 9598 11386
rect 9650 11376 9664 11386
rect 9716 11376 10152 11386
rect 10204 11376 10218 11428
rect 10270 11376 10706 11428
rect 10758 11376 10772 11428
rect 10824 11376 11260 11428
rect 11312 11376 11326 11428
rect 11378 11376 11814 11428
rect 11866 11376 11880 11428
rect 11932 11376 12368 11428
rect 12420 11376 12434 11428
rect 12486 11376 12922 11428
rect 12974 11376 12988 11428
rect 2950 11368 13040 11376
rect 13199 11846 13200 11898
rect 13252 11846 13270 11898
rect 13322 11846 13340 11898
rect 13392 11846 13410 11898
rect 13462 11846 13480 11898
rect 13532 11846 13550 11898
rect 13602 11846 14940 11898
rect 13199 11834 14940 11846
rect 13199 11782 13200 11834
rect 13252 11782 13270 11834
rect 13322 11782 13340 11834
rect 13392 11782 13410 11834
rect 13462 11782 13480 11834
rect 13532 11782 13550 11834
rect 13602 11782 14940 11834
rect 13199 11770 14940 11782
rect 13199 11718 13200 11770
rect 13252 11718 13270 11770
rect 13322 11718 13340 11770
rect 13392 11718 13410 11770
rect 13462 11718 13480 11770
rect 13532 11718 13550 11770
rect 13602 11718 14940 11770
rect 13199 11706 14940 11718
rect 13199 11654 13200 11706
rect 13252 11654 13270 11706
rect 13322 11654 13340 11706
rect 13392 11654 13410 11706
rect 13462 11654 13480 11706
rect 13532 11654 13550 11706
rect 13602 11654 14940 11706
rect 13199 11642 14940 11654
rect 13199 11590 13200 11642
rect 13252 11590 13270 11642
rect 13322 11590 13340 11642
rect 13392 11590 13410 11642
rect 13462 11590 13480 11642
rect 13532 11590 13550 11642
rect 13602 11590 14940 11642
rect 13199 11578 14940 11590
rect 13199 11526 13200 11578
rect 13252 11526 13270 11578
rect 13322 11526 13340 11578
rect 13392 11526 13410 11578
rect 13462 11526 13480 11578
rect 13532 11526 13550 11578
rect 13602 11526 14940 11578
rect 13199 11514 14940 11526
rect 13199 11462 13200 11514
rect 13252 11462 13270 11514
rect 13322 11462 13340 11514
rect 13392 11462 13410 11514
rect 13462 11462 13480 11514
rect 13532 11462 13550 11514
rect 13602 11462 14940 11514
rect 13199 11450 14940 11462
rect 13199 11398 13200 11450
rect 13252 11398 13270 11450
rect 13322 11398 13340 11450
rect 13392 11398 13410 11450
rect 13462 11398 13480 11450
rect 13532 11398 13550 11450
rect 13602 11398 14940 11450
rect 13199 11386 14940 11398
rect 13199 11334 13200 11386
rect 13252 11334 13270 11386
rect 13322 11334 13340 11386
rect 13392 11334 13410 11386
rect 13462 11334 13480 11386
rect 13532 11334 13550 11386
rect 13602 11334 14940 11386
rect 13199 11322 14940 11334
rect 13199 11270 13200 11322
rect 13252 11270 13270 11322
rect 13322 11270 13340 11322
rect 13392 11270 13410 11322
rect 13462 11270 13480 11322
rect 13532 11270 13550 11322
rect 13602 11270 14940 11322
rect 13199 11258 14940 11270
rect 13199 11206 13200 11258
rect 13252 11206 13270 11258
rect 13322 11206 13340 11258
rect 13392 11206 13410 11258
rect 13462 11206 13480 11258
rect 13532 11206 13550 11258
rect 13602 11206 14940 11258
rect 13199 11194 14940 11206
rect 13199 11142 13200 11194
rect 13252 11142 13270 11194
rect 13322 11142 13340 11194
rect 13392 11142 13410 11194
rect 13462 11142 13480 11194
rect 13532 11142 13550 11194
rect 13602 11142 14940 11194
rect 13199 11130 14940 11142
rect 13199 11078 13200 11130
rect 13252 11078 13270 11130
rect 13322 11078 13340 11130
rect 13392 11078 13410 11130
rect 13462 11078 13480 11130
rect 13532 11078 13550 11130
rect 13602 11078 14940 11130
rect 13199 11066 14940 11078
rect 13199 11014 13200 11066
rect 13252 11014 13270 11066
rect 13322 11014 13340 11066
rect 13392 11014 13410 11066
rect 13462 11014 13480 11066
rect 13532 11014 13550 11066
rect 13602 11014 14940 11066
rect 13199 11002 14940 11014
rect 13199 10950 13200 11002
rect 13252 10950 13270 11002
rect 13322 10950 13340 11002
rect 13392 10950 13410 11002
rect 13462 10950 13480 11002
rect 13532 10950 13550 11002
rect 13602 10950 14940 11002
rect 13199 10938 14940 10950
tri 13148 10886 13199 10937 se
rect 13199 10886 13200 10938
rect 13252 10886 13270 10938
rect 13322 10886 13340 10938
rect 13392 10886 13410 10938
rect 13462 10886 13480 10938
rect 13532 10886 13550 10938
rect 13602 10886 14940 10938
tri 13136 10874 13148 10886 se
rect 13148 10874 14940 10886
tri 13084 10822 13136 10874 se
rect 13136 10822 13200 10874
rect 13252 10822 13270 10874
rect 13322 10822 13340 10874
rect 13392 10822 13410 10874
rect 13462 10822 13480 10874
rect 13532 10822 13550 10874
rect 13602 10822 14940 10874
tri 13072 10810 13084 10822 se
rect 13084 10810 14940 10822
tri 13020 10758 13072 10810 se
rect 13072 10758 13200 10810
rect 13252 10758 13270 10810
rect 13322 10758 13340 10810
rect 13392 10758 13410 10810
rect 13462 10758 13480 10810
rect 13532 10758 13550 10810
rect 13602 10758 14940 10810
tri 13008 10746 13020 10758 se
rect 13020 10746 14940 10758
tri 12992 10730 13008 10746 se
rect 13008 10730 13200 10746
rect 3227 10724 13200 10730
rect 3279 10672 3293 10724
rect 3345 10672 3781 10724
rect 3833 10672 3847 10724
rect 3899 10672 4335 10724
rect 4387 10672 4401 10724
rect 4453 10672 4889 10724
rect 4941 10672 4955 10724
rect 5007 10672 5443 10724
rect 5495 10672 5509 10724
rect 5561 10672 5997 10724
rect 6049 10672 6063 10724
rect 6115 10672 6551 10724
rect 6603 10672 6617 10724
rect 6669 10672 7105 10724
rect 7157 10672 7171 10724
rect 7223 10672 7659 10724
rect 7711 10672 7725 10724
rect 7777 10672 8213 10724
rect 8265 10672 8279 10724
rect 8331 10672 8767 10724
rect 8819 10672 8833 10724
rect 8885 10672 9321 10724
rect 9373 10672 9387 10724
rect 9439 10672 9875 10724
rect 9927 10672 9941 10724
rect 9993 10672 10429 10724
rect 10481 10672 10495 10724
rect 10547 10672 10983 10724
rect 11035 10672 11049 10724
rect 11101 10672 11537 10724
rect 11589 10672 11603 10724
rect 11655 10672 12091 10724
rect 12143 10672 12157 10724
rect 12209 10672 12645 10724
rect 12697 10672 12711 10724
rect 12763 10694 13200 10724
rect 13252 10694 13270 10746
rect 13322 10694 13340 10746
rect 13392 10694 13410 10746
rect 13462 10694 13480 10746
rect 13532 10694 13550 10746
rect 13602 10694 14940 10746
rect 12763 10682 14940 10694
rect 12763 10672 13200 10682
rect 3227 10658 13200 10672
rect 3279 10606 3293 10658
rect 3345 10606 3781 10658
rect 3833 10606 3847 10658
rect 3899 10606 4335 10658
rect 4387 10606 4401 10658
rect 4453 10606 4889 10658
rect 4941 10606 4955 10658
rect 5007 10606 5443 10658
rect 5495 10606 5509 10658
rect 5561 10606 5997 10658
rect 6049 10606 6063 10658
rect 6115 10606 6551 10658
rect 6603 10606 6617 10658
rect 6669 10606 7105 10658
rect 7157 10606 7171 10658
rect 7223 10606 7659 10658
rect 7711 10606 7725 10658
rect 7777 10606 8213 10658
rect 8265 10606 8279 10658
rect 8331 10606 8767 10658
rect 8819 10606 8833 10658
rect 8885 10606 9321 10658
rect 9373 10606 9387 10658
rect 9439 10606 9875 10658
rect 9927 10606 9941 10658
rect 9993 10606 10429 10658
rect 10481 10606 10495 10658
rect 10547 10606 10983 10658
rect 11035 10606 11049 10658
rect 11101 10606 11537 10658
rect 11589 10606 11603 10658
rect 11655 10606 12091 10658
rect 12143 10606 12157 10658
rect 12209 10606 12645 10658
rect 12697 10606 12711 10658
rect 12763 10630 13200 10658
rect 13252 10630 13270 10682
rect 13322 10630 13340 10682
rect 13392 10630 13410 10682
rect 13462 10630 13480 10682
rect 13532 10630 13550 10682
rect 13602 10630 14940 10682
rect 12763 10618 14940 10630
rect 12763 10606 13200 10618
rect 3227 10592 13200 10606
rect 3279 10540 3293 10592
rect 3345 10540 3781 10592
rect 3833 10540 3847 10592
rect 3899 10540 4335 10592
rect 4387 10540 4401 10592
rect 4453 10540 4889 10592
rect 4941 10540 4955 10592
rect 5007 10540 5443 10592
rect 5495 10540 5509 10592
rect 5561 10540 5997 10592
rect 6049 10540 6063 10592
rect 6115 10540 6551 10592
rect 6603 10540 6617 10592
rect 6669 10540 7105 10592
rect 7157 10540 7171 10592
rect 7223 10540 7659 10592
rect 7711 10540 7725 10592
rect 7777 10540 8213 10592
rect 8265 10540 8279 10592
rect 8331 10540 8767 10592
rect 8819 10540 8833 10592
rect 8885 10540 9321 10592
rect 9373 10540 9387 10592
rect 9439 10540 9875 10592
rect 9927 10540 9941 10592
rect 9993 10540 10429 10592
rect 10481 10540 10495 10592
rect 10547 10540 10983 10592
rect 11035 10540 11049 10592
rect 11101 10540 11537 10592
rect 11589 10540 11603 10592
rect 11655 10540 12091 10592
rect 12143 10540 12157 10592
rect 12209 10540 12645 10592
rect 12697 10540 12711 10592
rect 12763 10566 13200 10592
rect 13252 10566 13270 10618
rect 13322 10566 13340 10618
rect 13392 10566 13410 10618
rect 13462 10566 13480 10618
rect 13532 10566 13550 10618
rect 13602 10566 14940 10618
rect 12763 10554 14940 10566
rect 12763 10540 13200 10554
rect 3227 10526 13200 10540
rect 3279 10474 3293 10526
rect 3345 10474 3781 10526
rect 3833 10474 3847 10526
rect 3899 10474 4335 10526
rect 4387 10474 4401 10526
rect 4453 10474 4889 10526
rect 4941 10474 4955 10526
rect 5007 10474 5443 10526
rect 5495 10474 5509 10526
rect 5561 10474 5997 10526
rect 6049 10474 6063 10526
rect 6115 10474 6551 10526
rect 6603 10474 6617 10526
rect 6669 10474 7105 10526
rect 7157 10474 7171 10526
rect 7223 10474 7659 10526
rect 7711 10474 7725 10526
rect 7777 10474 8213 10526
rect 8265 10474 8279 10526
rect 8331 10474 8767 10526
rect 8819 10474 8833 10526
rect 8885 10474 9321 10526
rect 9373 10474 9387 10526
rect 9439 10474 9875 10526
rect 9927 10474 9941 10526
rect 9993 10474 10429 10526
rect 10481 10474 10495 10526
rect 10547 10474 10983 10526
rect 11035 10474 11049 10526
rect 11101 10474 11537 10526
rect 11589 10474 11603 10526
rect 11655 10474 12091 10526
rect 12143 10474 12157 10526
rect 12209 10474 12645 10526
rect 12697 10474 12711 10526
rect 12763 10502 13200 10526
rect 13252 10502 13270 10554
rect 13322 10502 13340 10554
rect 13392 10502 13410 10554
rect 13462 10502 13480 10554
rect 13532 10502 13550 10554
rect 13602 10502 14940 10554
rect 12763 10490 14940 10502
rect 12763 10474 13200 10490
rect 3227 10460 13200 10474
rect 3279 10408 3293 10460
rect 3345 10408 3781 10460
rect 3833 10408 3847 10460
rect 3899 10408 4335 10460
rect 4387 10408 4401 10460
rect 4453 10408 4889 10460
rect 4941 10408 4955 10460
rect 5007 10408 5443 10460
rect 5495 10408 5509 10460
rect 5561 10408 5997 10460
rect 6049 10408 6063 10460
rect 6115 10408 6551 10460
rect 6603 10408 6617 10460
rect 6669 10408 7105 10460
rect 7157 10408 7171 10460
rect 7223 10408 7659 10460
rect 7711 10408 7725 10460
rect 7777 10408 8213 10460
rect 8265 10408 8279 10460
rect 8331 10408 8767 10460
rect 8819 10408 8833 10460
rect 8885 10408 9321 10460
rect 9373 10408 9387 10460
rect 9439 10408 9875 10460
rect 9927 10408 9941 10460
rect 9993 10408 10429 10460
rect 10481 10408 10495 10460
rect 10547 10408 10983 10460
rect 11035 10408 11049 10460
rect 11101 10408 11537 10460
rect 11589 10408 11603 10460
rect 11655 10408 12091 10460
rect 12143 10408 12157 10460
rect 12209 10408 12645 10460
rect 12697 10408 12711 10460
rect 12763 10438 13200 10460
rect 13252 10438 13270 10490
rect 13322 10438 13340 10490
rect 13392 10438 13410 10490
rect 13462 10438 13480 10490
rect 13532 10438 13550 10490
rect 13602 10438 14940 10490
rect 12763 10426 14940 10438
rect 12763 10408 13200 10426
rect 3227 10394 13200 10408
rect 3279 10342 3293 10394
rect 3345 10342 3781 10394
rect 3833 10342 3847 10394
rect 3899 10342 4335 10394
rect 4387 10342 4401 10394
rect 4453 10342 4889 10394
rect 4941 10342 4955 10394
rect 5007 10342 5443 10394
rect 5495 10342 5509 10394
rect 5561 10342 5997 10394
rect 6049 10342 6063 10394
rect 6115 10342 6551 10394
rect 6603 10342 6617 10394
rect 6669 10342 7105 10394
rect 7157 10342 7171 10394
rect 7223 10342 7659 10394
rect 7711 10342 7725 10394
rect 7777 10342 8213 10394
rect 8265 10342 8279 10394
rect 8331 10342 8767 10394
rect 8819 10342 8833 10394
rect 8885 10342 9321 10394
rect 9373 10342 9387 10394
rect 9439 10342 9875 10394
rect 9927 10342 9941 10394
rect 9993 10342 10429 10394
rect 10481 10342 10495 10394
rect 10547 10342 10983 10394
rect 11035 10342 11049 10394
rect 11101 10342 11537 10394
rect 11589 10342 11603 10394
rect 11655 10342 12091 10394
rect 12143 10342 12157 10394
rect 12209 10342 12645 10394
rect 12697 10342 12711 10394
rect 12763 10374 13200 10394
rect 13252 10374 13270 10426
rect 13322 10374 13340 10426
rect 13392 10374 13410 10426
rect 13462 10374 13480 10426
rect 13532 10374 13550 10426
rect 13602 10374 14940 10426
rect 12763 10362 14940 10374
rect 12763 10342 13200 10362
rect 3227 10327 13200 10342
rect 3279 10275 3293 10327
rect 3345 10275 3781 10327
rect 3833 10275 3847 10327
rect 3899 10275 4335 10327
rect 4387 10275 4401 10327
rect 4453 10275 4889 10327
rect 4941 10275 4955 10327
rect 5007 10275 5443 10327
rect 5495 10275 5509 10327
rect 5561 10275 5997 10327
rect 6049 10275 6063 10327
rect 6115 10275 6551 10327
rect 6603 10275 6617 10327
rect 6669 10275 7105 10327
rect 7157 10275 7171 10327
rect 7223 10275 7659 10327
rect 7711 10275 7725 10327
rect 7777 10275 8213 10327
rect 8265 10275 8279 10327
rect 8331 10275 8767 10327
rect 8819 10275 8833 10327
rect 8885 10275 9321 10327
rect 9373 10275 9387 10327
rect 9439 10275 9875 10327
rect 9927 10275 9941 10327
rect 9993 10275 10429 10327
rect 10481 10275 10495 10327
rect 10547 10275 10983 10327
rect 11035 10275 11049 10327
rect 11101 10275 11537 10327
rect 11589 10275 11603 10327
rect 11655 10275 12091 10327
rect 12143 10275 12157 10327
rect 12209 10275 12645 10327
rect 12697 10275 12711 10327
rect 12763 10310 13200 10327
rect 13252 10310 13270 10362
rect 13322 10310 13340 10362
rect 13392 10310 13410 10362
rect 13462 10310 13480 10362
rect 13532 10310 13550 10362
rect 13602 10310 14940 10362
rect 12763 10298 14940 10310
rect 12763 10275 13200 10298
rect 3227 10260 13200 10275
rect 3279 10208 3293 10260
rect 3345 10208 3781 10260
rect 3833 10208 3847 10260
rect 3899 10208 4335 10260
rect 4387 10208 4401 10260
rect 4453 10208 4889 10260
rect 4941 10208 4955 10260
rect 5007 10208 5443 10260
rect 5495 10208 5509 10260
rect 5561 10208 5997 10260
rect 6049 10208 6063 10260
rect 6115 10208 6551 10260
rect 6603 10208 6617 10260
rect 6669 10208 7105 10260
rect 7157 10208 7171 10260
rect 7223 10208 7659 10260
rect 7711 10208 7725 10260
rect 7777 10208 8213 10260
rect 8265 10208 8279 10260
rect 8331 10208 8767 10260
rect 8819 10208 8833 10260
rect 8885 10208 9321 10260
rect 9373 10208 9387 10260
rect 9439 10208 9875 10260
rect 9927 10208 9941 10260
rect 9993 10208 10429 10260
rect 10481 10208 10495 10260
rect 10547 10208 10983 10260
rect 11035 10208 11049 10260
rect 11101 10208 11537 10260
rect 11589 10208 11603 10260
rect 11655 10208 12091 10260
rect 12143 10208 12157 10260
rect 12209 10208 12645 10260
rect 12697 10208 12711 10260
rect 12763 10246 13200 10260
rect 13252 10246 13270 10298
rect 13322 10246 13340 10298
rect 13392 10246 13410 10298
rect 13462 10246 13480 10298
rect 13532 10246 13550 10298
rect 13602 10246 14940 10298
rect 12763 10234 14940 10246
rect 12763 10208 13200 10234
rect 3227 10202 13200 10208
tri 12989 10182 13009 10202 ne
rect 13009 10182 13200 10202
rect 13252 10182 13270 10234
rect 13322 10182 13340 10234
rect 13392 10182 13410 10234
rect 13462 10182 13480 10234
rect 13532 10182 13550 10234
rect 13602 10182 14940 10234
tri 13009 10170 13021 10182 ne
rect 13021 10170 14940 10182
tri 13021 10118 13073 10170 ne
rect 13073 10118 13200 10170
rect 13252 10118 13270 10170
rect 13322 10118 13340 10170
rect 13392 10118 13410 10170
rect 13462 10118 13480 10170
rect 13532 10118 13550 10170
rect 13602 10118 14940 10170
tri 13073 10106 13085 10118 ne
rect 13085 10106 14940 10118
tri 13085 10054 13137 10106 ne
rect 13137 10054 13200 10106
rect 13252 10054 13270 10106
rect 13322 10054 13340 10106
rect 13392 10054 13410 10106
rect 13462 10054 13480 10106
rect 13532 10054 13550 10106
rect 13602 10054 14940 10106
tri 13137 10042 13149 10054 ne
rect 13149 10042 14940 10054
tri 13149 9991 13200 10042 ne
rect 13252 9990 13270 10042
rect 13322 9990 13340 10042
rect 13392 9990 13410 10042
rect 13462 9990 13480 10042
rect 13532 9990 13550 10042
rect 13602 9990 14940 10042
rect 13200 9978 14940 9990
rect 13252 9926 13270 9978
rect 13322 9926 13340 9978
rect 13392 9926 13410 9978
rect 13462 9926 13480 9978
rect 13532 9926 13550 9978
rect 13602 9926 14940 9978
rect 13200 9914 14940 9926
rect 2950 9896 13040 9902
rect 3002 9844 3016 9896
rect 3068 9844 3504 9896
rect 3556 9844 3570 9896
rect 3622 9844 4058 9896
rect 4110 9844 4124 9896
rect 4176 9844 4612 9896
rect 4664 9844 4678 9896
rect 4730 9844 5166 9896
rect 5218 9844 5232 9896
rect 5284 9844 5720 9896
rect 5772 9844 5786 9896
rect 5838 9844 6274 9896
rect 6326 9844 6340 9896
rect 6392 9844 6828 9896
rect 6880 9844 6894 9896
rect 6946 9844 7382 9896
rect 7434 9844 7448 9896
rect 7500 9877 7936 9896
rect 7988 9877 8002 9896
rect 8054 9877 8490 9896
rect 8542 9877 8556 9896
rect 8608 9877 9044 9896
rect 9096 9877 9110 9896
rect 9162 9877 9598 9896
rect 9650 9877 9664 9896
rect 9716 9877 10152 9896
rect 7500 9844 7691 9877
rect 2950 9830 7691 9844
rect 3002 9778 3016 9830
rect 3068 9778 3504 9830
rect 3556 9778 3570 9830
rect 3622 9778 4058 9830
rect 4110 9778 4124 9830
rect 4176 9778 4612 9830
rect 4664 9778 4678 9830
rect 4730 9778 5166 9830
rect 5218 9778 5232 9830
rect 5284 9778 5720 9830
rect 5772 9778 5786 9830
rect 5838 9778 6274 9830
rect 6326 9778 6340 9830
rect 6392 9778 6828 9830
rect 6880 9778 6894 9830
rect 6946 9778 7382 9830
rect 7434 9778 7448 9830
rect 7500 9821 7691 9830
rect 7747 9821 7775 9877
rect 7831 9821 7858 9877
rect 7914 9844 7936 9877
rect 7997 9844 8002 9877
rect 7914 9830 7941 9844
rect 7997 9830 8024 9844
rect 7914 9821 7936 9830
rect 7997 9821 8002 9830
rect 8080 9821 8107 9877
rect 8163 9821 8190 9877
rect 8246 9821 8273 9877
rect 8329 9821 8356 9877
rect 8412 9821 8439 9877
rect 8495 9830 8522 9844
rect 8578 9830 8605 9844
rect 8661 9821 8688 9877
rect 8744 9821 8771 9877
rect 8827 9821 8854 9877
rect 8910 9821 8937 9877
rect 8993 9821 9020 9877
rect 9096 9844 9103 9877
rect 9162 9844 9186 9877
rect 9076 9830 9103 9844
rect 9159 9830 9186 9844
rect 9096 9821 9103 9830
rect 9162 9821 9186 9830
rect 9242 9821 9269 9877
rect 9325 9821 9352 9877
rect 9408 9821 9435 9877
rect 9491 9821 9518 9877
rect 9574 9844 9598 9877
rect 9657 9844 9664 9877
rect 9574 9830 9601 9844
rect 9657 9830 9684 9844
rect 9574 9821 9598 9830
rect 9657 9821 9664 9830
rect 9740 9821 9767 9877
rect 9823 9844 10152 9877
rect 10204 9844 10218 9896
rect 10270 9844 10706 9896
rect 10758 9844 10772 9896
rect 10824 9844 11260 9896
rect 11312 9844 11326 9896
rect 11378 9844 11814 9896
rect 11866 9844 11880 9896
rect 11932 9844 12368 9896
rect 12420 9844 12434 9896
rect 12486 9844 12922 9896
rect 12974 9844 12988 9896
rect 9823 9830 13040 9844
rect 9823 9821 10152 9830
rect 7500 9789 7936 9821
rect 7988 9789 8002 9821
rect 8054 9789 8490 9821
rect 8542 9789 8556 9821
rect 8608 9789 9044 9821
rect 9096 9789 9110 9821
rect 9162 9789 9598 9821
rect 9650 9789 9664 9821
rect 9716 9789 10152 9821
rect 7500 9778 7691 9789
rect 2950 9764 7691 9778
rect 3002 9712 3016 9764
rect 3068 9712 3504 9764
rect 3556 9712 3570 9764
rect 3622 9712 4058 9764
rect 4110 9712 4124 9764
rect 4176 9712 4612 9764
rect 4664 9712 4678 9764
rect 4730 9712 5166 9764
rect 5218 9712 5232 9764
rect 5284 9712 5720 9764
rect 5772 9712 5786 9764
rect 5838 9712 6274 9764
rect 6326 9712 6340 9764
rect 6392 9712 6828 9764
rect 6880 9712 6894 9764
rect 6946 9712 7382 9764
rect 7434 9712 7448 9764
rect 7500 9733 7691 9764
rect 7747 9733 7775 9789
rect 7831 9733 7858 9789
rect 7914 9778 7936 9789
rect 7997 9778 8002 9789
rect 7914 9764 7941 9778
rect 7997 9764 8024 9778
rect 7914 9733 7936 9764
rect 7997 9733 8002 9764
rect 8080 9733 8107 9789
rect 8163 9733 8190 9789
rect 8246 9733 8273 9789
rect 8329 9733 8356 9789
rect 8412 9733 8439 9789
rect 8495 9764 8522 9778
rect 8578 9764 8605 9778
rect 8661 9733 8688 9789
rect 8744 9733 8771 9789
rect 8827 9733 8854 9789
rect 8910 9733 8937 9789
rect 8993 9733 9020 9789
rect 9096 9778 9103 9789
rect 9162 9778 9186 9789
rect 9076 9764 9103 9778
rect 9159 9764 9186 9778
rect 9096 9733 9103 9764
rect 9162 9733 9186 9764
rect 9242 9733 9269 9789
rect 9325 9733 9352 9789
rect 9408 9733 9435 9789
rect 9491 9733 9518 9789
rect 9574 9778 9598 9789
rect 9657 9778 9664 9789
rect 9574 9764 9601 9778
rect 9657 9764 9684 9778
rect 9574 9733 9598 9764
rect 9657 9733 9664 9764
rect 9740 9733 9767 9789
rect 9823 9778 10152 9789
rect 10204 9778 10218 9830
rect 10270 9778 10706 9830
rect 10758 9778 10772 9830
rect 10824 9778 11260 9830
rect 11312 9778 11326 9830
rect 11378 9778 11814 9830
rect 11866 9778 11880 9830
rect 11932 9778 12368 9830
rect 12420 9778 12434 9830
rect 12486 9778 12922 9830
rect 12974 9778 12988 9830
rect 9823 9764 13040 9778
rect 9823 9733 10152 9764
rect 7500 9712 7936 9733
rect 7988 9712 8002 9733
rect 8054 9712 8490 9733
rect 8542 9712 8556 9733
rect 8608 9712 9044 9733
rect 9096 9712 9110 9733
rect 9162 9712 9598 9733
rect 9650 9712 9664 9733
rect 9716 9712 10152 9733
rect 10204 9712 10218 9764
rect 10270 9712 10706 9764
rect 10758 9712 10772 9764
rect 10824 9712 11260 9764
rect 11312 9712 11326 9764
rect 11378 9712 11814 9764
rect 11866 9712 11880 9764
rect 11932 9712 12368 9764
rect 12420 9712 12434 9764
rect 12486 9712 12922 9764
rect 12974 9712 12988 9764
rect 2950 9701 13040 9712
rect 2950 9698 7691 9701
rect 3002 9646 3016 9698
rect 3068 9646 3504 9698
rect 3556 9646 3570 9698
rect 3622 9646 4058 9698
rect 4110 9646 4124 9698
rect 4176 9646 4612 9698
rect 4664 9646 4678 9698
rect 4730 9646 5166 9698
rect 5218 9646 5232 9698
rect 5284 9646 5720 9698
rect 5772 9646 5786 9698
rect 5838 9646 6274 9698
rect 6326 9646 6340 9698
rect 6392 9646 6828 9698
rect 6880 9646 6894 9698
rect 6946 9646 7382 9698
rect 7434 9646 7448 9698
rect 7500 9646 7691 9698
rect 2950 9645 7691 9646
rect 7747 9645 7775 9701
rect 7831 9645 7858 9701
rect 7914 9698 7941 9701
rect 7997 9698 8024 9701
rect 7914 9646 7936 9698
rect 7997 9646 8002 9698
rect 7914 9645 7941 9646
rect 7997 9645 8024 9646
rect 8080 9645 8107 9701
rect 8163 9645 8190 9701
rect 8246 9645 8273 9701
rect 8329 9645 8356 9701
rect 8412 9645 8439 9701
rect 8495 9698 8522 9701
rect 8578 9698 8605 9701
rect 8495 9645 8522 9646
rect 8578 9645 8605 9646
rect 8661 9645 8688 9701
rect 8744 9645 8771 9701
rect 8827 9645 8854 9701
rect 8910 9645 8937 9701
rect 8993 9645 9020 9701
rect 9076 9698 9103 9701
rect 9159 9698 9186 9701
rect 9096 9646 9103 9698
rect 9162 9646 9186 9698
rect 9076 9645 9103 9646
rect 9159 9645 9186 9646
rect 9242 9645 9269 9701
rect 9325 9645 9352 9701
rect 9408 9645 9435 9701
rect 9491 9645 9518 9701
rect 9574 9698 9601 9701
rect 9657 9698 9684 9701
rect 9574 9646 9598 9698
rect 9657 9646 9664 9698
rect 9574 9645 9601 9646
rect 9657 9645 9684 9646
rect 9740 9645 9767 9701
rect 9823 9698 13040 9701
rect 9823 9646 10152 9698
rect 10204 9646 10218 9698
rect 10270 9646 10706 9698
rect 10758 9646 10772 9698
rect 10824 9646 11260 9698
rect 11312 9646 11326 9698
rect 11378 9646 11814 9698
rect 11866 9646 11880 9698
rect 11932 9646 12368 9698
rect 12420 9646 12434 9698
rect 12486 9646 12922 9698
rect 12974 9646 12988 9698
rect 9823 9645 13040 9646
rect 2950 9632 13040 9645
rect 3002 9580 3016 9632
rect 3068 9580 3504 9632
rect 3556 9580 3570 9632
rect 3622 9580 4058 9632
rect 4110 9580 4124 9632
rect 4176 9580 4612 9632
rect 4664 9580 4678 9632
rect 4730 9580 5166 9632
rect 5218 9580 5232 9632
rect 5284 9580 5720 9632
rect 5772 9580 5786 9632
rect 5838 9580 6274 9632
rect 6326 9580 6340 9632
rect 6392 9580 6828 9632
rect 6880 9580 6894 9632
rect 6946 9580 7382 9632
rect 7434 9580 7448 9632
rect 7500 9613 7936 9632
rect 7988 9613 8002 9632
rect 8054 9613 8490 9632
rect 8542 9613 8556 9632
rect 8608 9613 9044 9632
rect 9096 9613 9110 9632
rect 9162 9613 9598 9632
rect 9650 9613 9664 9632
rect 9716 9613 10152 9632
rect 7500 9580 7691 9613
rect 2950 9566 7691 9580
rect 3002 9514 3016 9566
rect 3068 9514 3504 9566
rect 3556 9514 3570 9566
rect 3622 9514 4058 9566
rect 4110 9514 4124 9566
rect 4176 9514 4612 9566
rect 4664 9514 4678 9566
rect 4730 9514 5166 9566
rect 5218 9514 5232 9566
rect 5284 9514 5720 9566
rect 5772 9514 5786 9566
rect 5838 9514 6274 9566
rect 6326 9514 6340 9566
rect 6392 9514 6828 9566
rect 6880 9514 6894 9566
rect 6946 9514 7382 9566
rect 7434 9514 7448 9566
rect 7500 9557 7691 9566
rect 7747 9557 7775 9613
rect 7831 9557 7858 9613
rect 7914 9580 7936 9613
rect 7997 9580 8002 9613
rect 7914 9566 7941 9580
rect 7997 9566 8024 9580
rect 7914 9557 7936 9566
rect 7997 9557 8002 9566
rect 8080 9557 8107 9613
rect 8163 9557 8190 9613
rect 8246 9557 8273 9613
rect 8329 9557 8356 9613
rect 8412 9557 8439 9613
rect 8495 9566 8522 9580
rect 8578 9566 8605 9580
rect 8661 9557 8688 9613
rect 8744 9557 8771 9613
rect 8827 9557 8854 9613
rect 8910 9557 8937 9613
rect 8993 9557 9020 9613
rect 9096 9580 9103 9613
rect 9162 9580 9186 9613
rect 9076 9566 9103 9580
rect 9159 9566 9186 9580
rect 9096 9557 9103 9566
rect 9162 9557 9186 9566
rect 9242 9557 9269 9613
rect 9325 9557 9352 9613
rect 9408 9557 9435 9613
rect 9491 9557 9518 9613
rect 9574 9580 9598 9613
rect 9657 9580 9664 9613
rect 9574 9566 9601 9580
rect 9657 9566 9684 9580
rect 9574 9557 9598 9566
rect 9657 9557 9664 9566
rect 9740 9557 9767 9613
rect 9823 9580 10152 9613
rect 10204 9580 10218 9632
rect 10270 9580 10706 9632
rect 10758 9580 10772 9632
rect 10824 9580 11260 9632
rect 11312 9580 11326 9632
rect 11378 9580 11814 9632
rect 11866 9580 11880 9632
rect 11932 9580 12368 9632
rect 12420 9580 12434 9632
rect 12486 9580 12922 9632
rect 12974 9580 12988 9632
rect 9823 9566 13040 9580
rect 9823 9557 10152 9566
rect 7500 9525 7936 9557
rect 7988 9525 8002 9557
rect 8054 9525 8490 9557
rect 8542 9525 8556 9557
rect 8608 9525 9044 9557
rect 9096 9525 9110 9557
rect 9162 9525 9598 9557
rect 9650 9525 9664 9557
rect 9716 9525 10152 9557
rect 7500 9514 7691 9525
rect 2950 9499 7691 9514
rect 3002 9447 3016 9499
rect 3068 9447 3504 9499
rect 3556 9447 3570 9499
rect 3622 9447 4058 9499
rect 4110 9447 4124 9499
rect 4176 9447 4612 9499
rect 4664 9447 4678 9499
rect 4730 9447 5166 9499
rect 5218 9447 5232 9499
rect 5284 9447 5720 9499
rect 5772 9447 5786 9499
rect 5838 9447 6274 9499
rect 6326 9447 6340 9499
rect 6392 9447 6828 9499
rect 6880 9447 6894 9499
rect 6946 9447 7382 9499
rect 7434 9447 7448 9499
rect 7500 9469 7691 9499
rect 7747 9469 7775 9525
rect 7831 9469 7858 9525
rect 7914 9514 7936 9525
rect 7997 9514 8002 9525
rect 7914 9499 7941 9514
rect 7997 9499 8024 9514
rect 7914 9469 7936 9499
rect 7997 9469 8002 9499
rect 8080 9469 8107 9525
rect 8163 9469 8190 9525
rect 8246 9469 8273 9525
rect 8329 9469 8356 9525
rect 8412 9469 8439 9525
rect 8495 9499 8522 9514
rect 8578 9499 8605 9514
rect 8661 9469 8688 9525
rect 8744 9469 8771 9525
rect 8827 9469 8854 9525
rect 8910 9469 8937 9525
rect 8993 9469 9020 9525
rect 9096 9514 9103 9525
rect 9162 9514 9186 9525
rect 9076 9499 9103 9514
rect 9159 9499 9186 9514
rect 9096 9469 9103 9499
rect 9162 9469 9186 9499
rect 9242 9469 9269 9525
rect 9325 9469 9352 9525
rect 9408 9469 9435 9525
rect 9491 9469 9518 9525
rect 9574 9514 9598 9525
rect 9657 9514 9664 9525
rect 9574 9499 9601 9514
rect 9657 9499 9684 9514
rect 9574 9469 9598 9499
rect 9657 9469 9664 9499
rect 9740 9469 9767 9525
rect 9823 9514 10152 9525
rect 10204 9514 10218 9566
rect 10270 9514 10706 9566
rect 10758 9514 10772 9566
rect 10824 9514 11260 9566
rect 11312 9514 11326 9566
rect 11378 9514 11814 9566
rect 11866 9514 11880 9566
rect 11932 9514 12368 9566
rect 12420 9514 12434 9566
rect 12486 9514 12922 9566
rect 12974 9514 12988 9566
rect 9823 9499 13040 9514
rect 9823 9469 10152 9499
rect 7500 9447 7936 9469
rect 7988 9447 8002 9469
rect 8054 9447 8490 9469
rect 8542 9447 8556 9469
rect 8608 9447 9044 9469
rect 9096 9447 9110 9469
rect 9162 9447 9598 9469
rect 9650 9447 9664 9469
rect 9716 9447 10152 9469
rect 10204 9447 10218 9499
rect 10270 9447 10706 9499
rect 10758 9447 10772 9499
rect 10824 9447 11260 9499
rect 11312 9447 11326 9499
rect 11378 9447 11814 9499
rect 11866 9447 11880 9499
rect 11932 9447 12368 9499
rect 12420 9447 12434 9499
rect 12486 9447 12922 9499
rect 12974 9447 12988 9499
rect 2950 9437 13040 9447
rect 2950 9432 7691 9437
rect 3002 9380 3016 9432
rect 3068 9380 3504 9432
rect 3556 9380 3570 9432
rect 3622 9380 4058 9432
rect 4110 9380 4124 9432
rect 4176 9380 4612 9432
rect 4664 9380 4678 9432
rect 4730 9380 5166 9432
rect 5218 9380 5232 9432
rect 5284 9380 5720 9432
rect 5772 9380 5786 9432
rect 5838 9380 6274 9432
rect 6326 9380 6340 9432
rect 6392 9380 6828 9432
rect 6880 9380 6894 9432
rect 6946 9380 7382 9432
rect 7434 9380 7448 9432
rect 7500 9381 7691 9432
rect 7747 9381 7775 9437
rect 7831 9381 7858 9437
rect 7914 9432 7941 9437
rect 7997 9432 8024 9437
rect 7914 9381 7936 9432
rect 7997 9381 8002 9432
rect 8080 9381 8107 9437
rect 8163 9381 8190 9437
rect 8246 9381 8273 9437
rect 8329 9381 8356 9437
rect 8412 9381 8439 9437
rect 8495 9432 8522 9437
rect 8578 9432 8605 9437
rect 8661 9381 8688 9437
rect 8744 9381 8771 9437
rect 8827 9381 8854 9437
rect 8910 9381 8937 9437
rect 8993 9381 9020 9437
rect 9076 9432 9103 9437
rect 9159 9432 9186 9437
rect 9096 9381 9103 9432
rect 9162 9381 9186 9432
rect 9242 9381 9269 9437
rect 9325 9381 9352 9437
rect 9408 9381 9435 9437
rect 9491 9381 9518 9437
rect 9574 9432 9601 9437
rect 9657 9432 9684 9437
rect 9574 9381 9598 9432
rect 9657 9381 9664 9432
rect 9740 9381 9767 9437
rect 9823 9432 13040 9437
rect 9823 9381 10152 9432
rect 7500 9380 7936 9381
rect 7988 9380 8002 9381
rect 8054 9380 8490 9381
rect 8542 9380 8556 9381
rect 8608 9380 9044 9381
rect 9096 9380 9110 9381
rect 9162 9380 9598 9381
rect 9650 9380 9664 9381
rect 9716 9380 10152 9381
rect 10204 9380 10218 9432
rect 10270 9380 10706 9432
rect 10758 9380 10772 9432
rect 10824 9380 11260 9432
rect 11312 9380 11326 9432
rect 11378 9380 11814 9432
rect 11866 9380 11880 9432
rect 11932 9380 12368 9432
rect 12420 9380 12434 9432
rect 12486 9380 12922 9432
rect 12974 9380 12988 9432
rect 2950 9372 13040 9380
rect 13252 9862 13270 9914
rect 13322 9862 13340 9914
rect 13392 9862 13410 9914
rect 13462 9862 13480 9914
rect 13532 9862 13550 9914
rect 13602 9862 14940 9914
rect 13200 9850 14940 9862
rect 13252 9798 13270 9850
rect 13322 9798 13340 9850
rect 13392 9798 13410 9850
rect 13462 9798 13480 9850
rect 13532 9798 13550 9850
rect 13602 9798 14940 9850
rect 13200 9786 14940 9798
rect 13252 9734 13270 9786
rect 13322 9734 13340 9786
rect 13392 9734 13410 9786
rect 13462 9734 13480 9786
rect 13532 9734 13550 9786
rect 13602 9734 14940 9786
rect 13200 9722 14940 9734
rect 13252 9670 13270 9722
rect 13322 9670 13340 9722
rect 13392 9670 13410 9722
rect 13462 9670 13480 9722
rect 13532 9670 13550 9722
rect 13602 9670 14940 9722
rect 13200 9658 14940 9670
rect 13252 9606 13270 9658
rect 13322 9606 13340 9658
rect 13392 9606 13410 9658
rect 13462 9606 13480 9658
rect 13532 9606 13550 9658
rect 13602 9606 14940 9658
rect 13200 9594 14940 9606
rect 13252 9542 13270 9594
rect 13322 9542 13340 9594
rect 13392 9542 13410 9594
rect 13462 9542 13480 9594
rect 13532 9542 13550 9594
rect 13602 9542 14940 9594
rect 13200 9530 14940 9542
rect 13252 9478 13270 9530
rect 13322 9478 13340 9530
rect 13392 9478 13410 9530
rect 13462 9478 13480 9530
rect 13532 9478 13550 9530
rect 13602 9478 14940 9530
rect 13200 9466 14940 9478
rect 13252 9414 13270 9466
rect 13322 9414 13340 9466
rect 13392 9414 13410 9466
rect 13462 9414 13480 9466
rect 13532 9414 13550 9466
rect 13602 9414 14940 9466
rect 13200 9402 14940 9414
rect 13252 9350 13270 9402
rect 13322 9350 13340 9402
rect 13392 9350 13410 9402
rect 13462 9350 13480 9402
rect 13532 9350 13550 9402
rect 13602 9350 14940 9402
rect 13200 9338 14940 9350
rect 13252 9286 13270 9338
rect 13322 9286 13340 9338
rect 13392 9286 13410 9338
rect 13462 9286 13480 9338
rect 13532 9286 13550 9338
rect 13602 9286 14940 9338
rect 13200 9274 14940 9286
rect 13252 9222 13270 9274
rect 13322 9222 13340 9274
rect 13392 9222 13410 9274
rect 13462 9222 13480 9274
rect 13532 9222 13550 9274
rect 13602 9222 14940 9274
rect 13200 9210 14940 9222
rect 13252 9158 13270 9210
rect 13322 9158 13340 9210
rect 13392 9158 13410 9210
rect 13462 9158 13480 9210
rect 13532 9158 13550 9210
rect 13602 9158 14940 9210
rect 13200 9146 14940 9158
rect 13252 9094 13270 9146
rect 13322 9094 13340 9146
rect 13392 9094 13410 9146
rect 13462 9094 13480 9146
rect 13532 9094 13550 9146
rect 13602 9094 14940 9146
rect 13200 9082 14940 9094
rect 13252 9030 13270 9082
rect 13322 9030 13340 9082
rect 13392 9030 13410 9082
rect 13462 9030 13480 9082
rect 13532 9030 13550 9082
rect 13602 9030 14940 9082
rect 13200 9018 14940 9030
rect 13252 8966 13270 9018
rect 13322 8966 13340 9018
rect 13392 8966 13410 9018
rect 13462 8966 13480 9018
rect 13532 8966 13550 9018
rect 13602 8966 14940 9018
rect 13200 8954 14940 8966
tri 13168 8902 13200 8934 se
rect 13252 8902 13270 8954
rect 13322 8902 13340 8954
rect 13392 8902 13410 8954
rect 13462 8902 13480 8954
rect 13532 8902 13550 8954
rect 13602 8902 14940 8954
tri 13156 8890 13168 8902 se
rect 13168 8890 14940 8902
tri 13104 8838 13156 8890 se
rect 13156 8838 13200 8890
rect 13252 8838 13270 8890
rect 13322 8838 13340 8890
rect 13392 8838 13410 8890
rect 13462 8838 13480 8890
rect 13532 8838 13550 8890
rect 13602 8838 14940 8890
tri 13092 8826 13104 8838 se
rect 13104 8826 14940 8838
tri 13040 8774 13092 8826 se
rect 13092 8774 13200 8826
rect 13252 8774 13270 8826
rect 13322 8774 13340 8826
rect 13392 8774 13410 8826
rect 13462 8774 13480 8826
rect 13532 8774 13550 8826
rect 13602 8774 14940 8826
tri 13028 8762 13040 8774 se
rect 13040 8762 14940 8774
tri 12992 8726 13028 8762 se
rect 13028 8726 13200 8762
rect 3227 8720 13200 8726
rect 3279 8668 3293 8720
rect 3345 8668 3781 8720
rect 3833 8668 3847 8720
rect 3899 8668 4335 8720
rect 4387 8668 4401 8720
rect 4453 8668 4889 8720
rect 4941 8668 4955 8720
rect 5007 8668 5443 8720
rect 5495 8668 5509 8720
rect 5561 8668 5997 8720
rect 6049 8668 6063 8720
rect 6115 8668 6551 8720
rect 6603 8668 6617 8720
rect 6669 8668 7105 8720
rect 7157 8668 7171 8720
rect 7223 8668 7659 8720
rect 7711 8668 7725 8720
rect 7777 8668 8213 8720
rect 8265 8668 8279 8720
rect 8331 8668 8767 8720
rect 8819 8668 8833 8720
rect 8885 8668 9321 8720
rect 9373 8668 9387 8720
rect 9439 8668 9875 8720
rect 9927 8668 9941 8720
rect 9993 8668 10429 8720
rect 10481 8668 10495 8720
rect 10547 8668 10983 8720
rect 11035 8668 11049 8720
rect 11101 8668 11537 8720
rect 11589 8668 11603 8720
rect 11655 8668 12091 8720
rect 12143 8668 12157 8720
rect 12209 8668 12645 8720
rect 12697 8668 12711 8720
rect 12763 8710 13200 8720
rect 13252 8710 13270 8762
rect 13322 8710 13340 8762
rect 13392 8710 13410 8762
rect 13462 8710 13480 8762
rect 13532 8710 13550 8762
rect 13602 8710 14940 8762
rect 12763 8698 14940 8710
rect 12763 8668 13200 8698
rect 3227 8654 13200 8668
rect 3279 8602 3293 8654
rect 3345 8602 3781 8654
rect 3833 8602 3847 8654
rect 3899 8602 4335 8654
rect 4387 8602 4401 8654
rect 4453 8602 4889 8654
rect 4941 8602 4955 8654
rect 5007 8602 5443 8654
rect 5495 8602 5509 8654
rect 5561 8602 5997 8654
rect 6049 8602 6063 8654
rect 6115 8602 6551 8654
rect 6603 8602 6617 8654
rect 6669 8602 7105 8654
rect 7157 8602 7171 8654
rect 7223 8602 7659 8654
rect 7711 8602 7725 8654
rect 7777 8602 8213 8654
rect 8265 8602 8279 8654
rect 8331 8602 8767 8654
rect 8819 8602 8833 8654
rect 8885 8602 9321 8654
rect 9373 8602 9387 8654
rect 9439 8602 9875 8654
rect 9927 8602 9941 8654
rect 9993 8602 10429 8654
rect 10481 8602 10495 8654
rect 10547 8602 10983 8654
rect 11035 8602 11049 8654
rect 11101 8602 11537 8654
rect 11589 8602 11603 8654
rect 11655 8602 12091 8654
rect 12143 8602 12157 8654
rect 12209 8602 12645 8654
rect 12697 8602 12711 8654
rect 12763 8646 13200 8654
rect 13252 8646 13270 8698
rect 13322 8646 13340 8698
rect 13392 8646 13410 8698
rect 13462 8646 13480 8698
rect 13532 8646 13550 8698
rect 13602 8646 14940 8698
rect 12763 8634 14940 8646
rect 12763 8602 13200 8634
rect 3227 8588 13200 8602
rect 3279 8536 3293 8588
rect 3345 8536 3781 8588
rect 3833 8536 3847 8588
rect 3899 8536 4335 8588
rect 4387 8536 4401 8588
rect 4453 8536 4889 8588
rect 4941 8536 4955 8588
rect 5007 8536 5443 8588
rect 5495 8536 5509 8588
rect 5561 8536 5997 8588
rect 6049 8536 6063 8588
rect 6115 8536 6551 8588
rect 6603 8536 6617 8588
rect 6669 8536 7105 8588
rect 7157 8536 7171 8588
rect 7223 8536 7659 8588
rect 7711 8536 7725 8588
rect 7777 8536 8213 8588
rect 8265 8536 8279 8588
rect 8331 8536 8767 8588
rect 8819 8536 8833 8588
rect 8885 8536 9321 8588
rect 9373 8536 9387 8588
rect 9439 8536 9875 8588
rect 9927 8536 9941 8588
rect 9993 8536 10429 8588
rect 10481 8536 10495 8588
rect 10547 8536 10983 8588
rect 11035 8536 11049 8588
rect 11101 8536 11537 8588
rect 11589 8536 11603 8588
rect 11655 8536 12091 8588
rect 12143 8536 12157 8588
rect 12209 8536 12645 8588
rect 12697 8536 12711 8588
rect 12763 8582 13200 8588
rect 13252 8582 13270 8634
rect 13322 8582 13340 8634
rect 13392 8582 13410 8634
rect 13462 8582 13480 8634
rect 13532 8582 13550 8634
rect 13602 8582 14940 8634
rect 12763 8570 14940 8582
rect 12763 8536 13200 8570
rect 3227 8522 13200 8536
rect 3279 8470 3293 8522
rect 3345 8470 3781 8522
rect 3833 8470 3847 8522
rect 3899 8470 4335 8522
rect 4387 8470 4401 8522
rect 4453 8470 4889 8522
rect 4941 8470 4955 8522
rect 5007 8470 5443 8522
rect 5495 8470 5509 8522
rect 5561 8470 5997 8522
rect 6049 8470 6063 8522
rect 6115 8470 6551 8522
rect 6603 8470 6617 8522
rect 6669 8470 7105 8522
rect 7157 8470 7171 8522
rect 7223 8470 7659 8522
rect 7711 8470 7725 8522
rect 7777 8470 8213 8522
rect 8265 8470 8279 8522
rect 8331 8470 8767 8522
rect 8819 8470 8833 8522
rect 8885 8470 9321 8522
rect 9373 8470 9387 8522
rect 9439 8470 9875 8522
rect 9927 8470 9941 8522
rect 9993 8470 10429 8522
rect 10481 8470 10495 8522
rect 10547 8470 10983 8522
rect 11035 8470 11049 8522
rect 11101 8470 11537 8522
rect 11589 8470 11603 8522
rect 11655 8470 12091 8522
rect 12143 8470 12157 8522
rect 12209 8470 12645 8522
rect 12697 8470 12711 8522
rect 12763 8518 13200 8522
rect 13252 8518 13270 8570
rect 13322 8518 13340 8570
rect 13392 8518 13410 8570
rect 13462 8518 13480 8570
rect 13532 8518 13550 8570
rect 13602 8518 14940 8570
rect 12763 8506 14940 8518
rect 12763 8470 13200 8506
rect 3227 8456 13200 8470
rect 3279 8404 3293 8456
rect 3345 8404 3781 8456
rect 3833 8404 3847 8456
rect 3899 8404 4335 8456
rect 4387 8404 4401 8456
rect 4453 8404 4889 8456
rect 4941 8404 4955 8456
rect 5007 8404 5443 8456
rect 5495 8404 5509 8456
rect 5561 8404 5997 8456
rect 6049 8404 6063 8456
rect 6115 8404 6551 8456
rect 6603 8404 6617 8456
rect 6669 8404 7105 8456
rect 7157 8404 7171 8456
rect 7223 8404 7659 8456
rect 7711 8404 7725 8456
rect 7777 8404 8213 8456
rect 8265 8404 8279 8456
rect 8331 8404 8767 8456
rect 8819 8404 8833 8456
rect 8885 8404 9321 8456
rect 9373 8404 9387 8456
rect 9439 8404 9875 8456
rect 9927 8404 9941 8456
rect 9993 8404 10429 8456
rect 10481 8404 10495 8456
rect 10547 8404 10983 8456
rect 11035 8404 11049 8456
rect 11101 8404 11537 8456
rect 11589 8404 11603 8456
rect 11655 8404 12091 8456
rect 12143 8404 12157 8456
rect 12209 8404 12645 8456
rect 12697 8404 12711 8456
rect 12763 8454 13200 8456
rect 13252 8454 13270 8506
rect 13322 8454 13340 8506
rect 13392 8454 13410 8506
rect 13462 8454 13480 8506
rect 13532 8454 13550 8506
rect 13602 8454 14940 8506
rect 12763 8442 14940 8454
rect 12763 8404 13200 8442
rect 3227 8390 13200 8404
rect 13252 8390 13270 8442
rect 13322 8390 13340 8442
rect 13392 8390 13410 8442
rect 13462 8390 13480 8442
rect 13532 8390 13550 8442
rect 13602 8390 14940 8442
rect 3279 8338 3293 8390
rect 3345 8338 3781 8390
rect 3833 8338 3847 8390
rect 3899 8338 4335 8390
rect 4387 8338 4401 8390
rect 4453 8338 4889 8390
rect 4941 8338 4955 8390
rect 5007 8338 5443 8390
rect 5495 8338 5509 8390
rect 5561 8338 5997 8390
rect 6049 8338 6063 8390
rect 6115 8338 6551 8390
rect 6603 8338 6617 8390
rect 6669 8338 7105 8390
rect 7157 8338 7171 8390
rect 7223 8338 7659 8390
rect 7711 8338 7725 8390
rect 7777 8338 8213 8390
rect 8265 8338 8279 8390
rect 8331 8338 8767 8390
rect 8819 8338 8833 8390
rect 8885 8338 9321 8390
rect 9373 8338 9387 8390
rect 9439 8338 9875 8390
rect 9927 8338 9941 8390
rect 9993 8338 10429 8390
rect 10481 8338 10495 8390
rect 10547 8338 10983 8390
rect 11035 8338 11049 8390
rect 11101 8338 11537 8390
rect 11589 8338 11603 8390
rect 11655 8338 12091 8390
rect 12143 8338 12157 8390
rect 12209 8338 12645 8390
rect 12697 8338 12711 8390
rect 12763 8378 14940 8390
rect 12763 8338 13200 8378
rect 3227 8326 13200 8338
rect 13252 8326 13270 8378
rect 13322 8326 13340 8378
rect 13392 8326 13410 8378
rect 13462 8326 13480 8378
rect 13532 8326 13550 8378
rect 13602 8326 14940 8378
rect 3227 8323 14940 8326
rect 3279 8271 3293 8323
rect 3345 8271 3781 8323
rect 3833 8271 3847 8323
rect 3899 8271 4335 8323
rect 4387 8271 4401 8323
rect 4453 8271 4889 8323
rect 4941 8271 4955 8323
rect 5007 8271 5443 8323
rect 5495 8271 5509 8323
rect 5561 8271 5997 8323
rect 6049 8271 6063 8323
rect 6115 8271 6551 8323
rect 6603 8271 6617 8323
rect 6669 8271 7105 8323
rect 7157 8271 7171 8323
rect 7223 8271 7659 8323
rect 7711 8271 7725 8323
rect 7777 8271 8213 8323
rect 8265 8271 8279 8323
rect 8331 8271 8767 8323
rect 8819 8271 8833 8323
rect 8885 8271 9321 8323
rect 9373 8271 9387 8323
rect 9439 8271 9875 8323
rect 9927 8271 9941 8323
rect 9993 8271 10429 8323
rect 10481 8271 10495 8323
rect 10547 8271 10983 8323
rect 11035 8271 11049 8323
rect 11101 8271 11537 8323
rect 11589 8271 11603 8323
rect 11655 8271 12091 8323
rect 12143 8271 12157 8323
rect 12209 8271 12645 8323
rect 12697 8271 12711 8323
rect 12763 8314 14940 8323
rect 12763 8271 13200 8314
rect 3227 8262 13200 8271
rect 13252 8262 13270 8314
rect 13322 8262 13340 8314
rect 13392 8262 13410 8314
rect 13462 8262 13480 8314
rect 13532 8262 13550 8314
rect 13602 8262 14940 8314
rect 3227 8256 14940 8262
rect 3279 8204 3293 8256
rect 3345 8204 3781 8256
rect 3833 8204 3847 8256
rect 3899 8204 4335 8256
rect 4387 8204 4401 8256
rect 4453 8204 4889 8256
rect 4941 8204 4955 8256
rect 5007 8204 5443 8256
rect 5495 8204 5509 8256
rect 5561 8204 5997 8256
rect 6049 8204 6063 8256
rect 6115 8204 6551 8256
rect 6603 8204 6617 8256
rect 6669 8204 7105 8256
rect 7157 8204 7171 8256
rect 7223 8204 7659 8256
rect 7711 8204 7725 8256
rect 7777 8204 8213 8256
rect 8265 8204 8279 8256
rect 8331 8204 8767 8256
rect 8819 8204 8833 8256
rect 8885 8204 9321 8256
rect 9373 8204 9387 8256
rect 9439 8204 9875 8256
rect 9927 8204 9941 8256
rect 9993 8204 10429 8256
rect 10481 8204 10495 8256
rect 10547 8204 10983 8256
rect 11035 8204 11049 8256
rect 11101 8204 11537 8256
rect 11589 8204 11603 8256
rect 11655 8204 12091 8256
rect 12143 8204 12157 8256
rect 12209 8204 12645 8256
rect 12697 8204 12711 8256
rect 12763 8250 14940 8256
rect 12763 8204 13200 8250
rect 3227 8198 13200 8204
rect 13252 8198 13270 8250
rect 13322 8198 13340 8250
rect 13392 8198 13410 8250
rect 13462 8198 13480 8250
rect 13532 8198 13550 8250
rect 13602 8198 14940 8250
tri 12989 8186 13001 8198 ne
rect 13001 8186 14940 8198
tri 13001 8134 13053 8186 ne
rect 13053 8134 13200 8186
rect 13252 8134 13270 8186
rect 13322 8134 13340 8186
rect 13392 8134 13410 8186
rect 13462 8134 13480 8186
rect 13532 8134 13550 8186
rect 13602 8134 14940 8186
tri 13053 8122 13065 8134 ne
rect 13065 8122 14940 8134
tri 13065 8070 13117 8122 ne
rect 13117 8070 13200 8122
rect 13252 8070 13270 8122
rect 13322 8070 13340 8122
rect 13392 8070 13410 8122
rect 13462 8070 13480 8122
rect 13532 8070 13550 8122
rect 13602 8070 14940 8122
tri 13117 8058 13129 8070 ne
rect 13129 8058 14940 8070
tri 13129 8006 13181 8058 ne
rect 13181 8006 13200 8058
rect 13252 8006 13270 8058
rect 13322 8006 13340 8058
rect 13392 8006 13410 8058
rect 13462 8006 13480 8058
rect 13532 8006 13550 8058
rect 13602 8006 14940 8058
tri 13181 7994 13193 8006 ne
rect 13193 7994 14940 8006
tri 13193 7987 13200 7994 ne
rect 13252 7942 13270 7994
rect 13322 7942 13340 7994
rect 13392 7942 13410 7994
rect 13462 7942 13480 7994
rect 13532 7942 13550 7994
rect 13602 7942 14940 7994
rect 13200 7930 14940 7942
rect 2950 7892 13040 7898
rect 3002 7840 3016 7892
rect 3068 7840 3504 7892
rect 3556 7840 3570 7892
rect 3622 7840 4058 7892
rect 4110 7840 4124 7892
rect 4176 7840 4612 7892
rect 4664 7840 4678 7892
rect 4730 7840 5166 7892
rect 5218 7840 5232 7892
rect 5284 7840 5720 7892
rect 5772 7840 5786 7892
rect 5838 7840 6274 7892
rect 6326 7840 6340 7892
rect 6392 7840 6828 7892
rect 6880 7840 6894 7892
rect 6946 7840 7382 7892
rect 7434 7840 7448 7892
rect 7500 7882 7936 7892
rect 7988 7882 8002 7892
rect 8054 7882 8490 7892
rect 8542 7882 8556 7892
rect 8608 7882 9044 7892
rect 9096 7882 9110 7892
rect 9162 7882 9598 7892
rect 9650 7882 9664 7892
rect 9716 7882 10152 7892
rect 7500 7840 7691 7882
rect 2950 7826 7691 7840
rect 7747 7826 7775 7882
rect 7831 7826 7858 7882
rect 7914 7840 7936 7882
rect 7997 7840 8002 7882
rect 7914 7826 7941 7840
rect 7997 7826 8024 7840
rect 8080 7826 8107 7882
rect 8163 7826 8190 7882
rect 8246 7826 8273 7882
rect 8329 7826 8356 7882
rect 8412 7826 8439 7882
rect 8495 7826 8522 7840
rect 8578 7826 8605 7840
rect 8661 7826 8688 7882
rect 8744 7826 8771 7882
rect 8827 7826 8854 7882
rect 8910 7826 8937 7882
rect 8993 7826 9020 7882
rect 9096 7840 9103 7882
rect 9162 7840 9186 7882
rect 9076 7826 9103 7840
rect 9159 7826 9186 7840
rect 9242 7826 9269 7882
rect 9325 7826 9352 7882
rect 9408 7826 9435 7882
rect 9491 7826 9518 7882
rect 9574 7840 9598 7882
rect 9657 7840 9664 7882
rect 9574 7826 9601 7840
rect 9657 7826 9684 7840
rect 9740 7826 9767 7882
rect 9823 7840 10152 7882
rect 10204 7840 10218 7892
rect 10270 7840 10706 7892
rect 10758 7840 10772 7892
rect 10824 7840 11260 7892
rect 11312 7840 11326 7892
rect 11378 7840 11814 7892
rect 11866 7840 11880 7892
rect 11932 7891 13040 7892
rect 11932 7840 12368 7891
rect 9823 7839 12368 7840
rect 12420 7839 12434 7891
rect 12486 7839 12922 7891
rect 12974 7839 12988 7891
rect 9823 7826 13040 7839
rect 3002 7774 3016 7826
rect 3068 7774 3504 7826
rect 3556 7774 3570 7826
rect 3622 7774 4058 7826
rect 4110 7774 4124 7826
rect 4176 7774 4612 7826
rect 4664 7774 4678 7826
rect 4730 7774 5166 7826
rect 5218 7774 5232 7826
rect 5284 7774 5720 7826
rect 5772 7774 5786 7826
rect 5838 7774 6274 7826
rect 6326 7774 6340 7826
rect 6392 7774 6828 7826
rect 6880 7774 6894 7826
rect 6946 7774 7382 7826
rect 7434 7774 7448 7826
rect 7500 7794 7936 7826
rect 7988 7794 8002 7826
rect 8054 7794 8490 7826
rect 8542 7794 8556 7826
rect 8608 7794 9044 7826
rect 9096 7794 9110 7826
rect 9162 7794 9598 7826
rect 9650 7794 9664 7826
rect 9716 7794 10152 7826
rect 7500 7774 7691 7794
rect 2950 7760 7691 7774
rect 3002 7708 3016 7760
rect 3068 7708 3504 7760
rect 3556 7708 3570 7760
rect 3622 7708 4058 7760
rect 4110 7708 4124 7760
rect 4176 7708 4612 7760
rect 4664 7708 4678 7760
rect 4730 7708 5166 7760
rect 5218 7708 5232 7760
rect 5284 7708 5720 7760
rect 5772 7708 5786 7760
rect 5838 7708 6274 7760
rect 6326 7708 6340 7760
rect 6392 7708 6828 7760
rect 6880 7708 6894 7760
rect 6946 7708 7382 7760
rect 7434 7708 7448 7760
rect 7500 7738 7691 7760
rect 7747 7738 7775 7794
rect 7831 7738 7858 7794
rect 7914 7774 7936 7794
rect 7997 7774 8002 7794
rect 7914 7760 7941 7774
rect 7997 7760 8024 7774
rect 7914 7738 7936 7760
rect 7997 7738 8002 7760
rect 8080 7738 8107 7794
rect 8163 7738 8190 7794
rect 8246 7738 8273 7794
rect 8329 7738 8356 7794
rect 8412 7738 8439 7794
rect 8495 7760 8522 7774
rect 8578 7760 8605 7774
rect 8661 7738 8688 7794
rect 8744 7738 8771 7794
rect 8827 7738 8854 7794
rect 8910 7738 8937 7794
rect 8993 7738 9020 7794
rect 9096 7774 9103 7794
rect 9162 7774 9186 7794
rect 9076 7760 9103 7774
rect 9159 7760 9186 7774
rect 9096 7738 9103 7760
rect 9162 7738 9186 7760
rect 9242 7738 9269 7794
rect 9325 7738 9352 7794
rect 9408 7738 9435 7794
rect 9491 7738 9518 7794
rect 9574 7774 9598 7794
rect 9657 7774 9664 7794
rect 9574 7760 9601 7774
rect 9657 7760 9684 7774
rect 9574 7738 9598 7760
rect 9657 7738 9664 7760
rect 9740 7738 9767 7794
rect 9823 7774 10152 7794
rect 10204 7774 10218 7826
rect 10270 7774 10706 7826
rect 10758 7774 10772 7826
rect 10824 7774 11260 7826
rect 11312 7774 11326 7826
rect 11378 7774 11814 7826
rect 11866 7774 11880 7826
rect 11932 7825 13040 7826
rect 11932 7774 12368 7825
rect 9823 7773 12368 7774
rect 12420 7773 12434 7825
rect 12486 7773 12922 7825
rect 12974 7773 12988 7825
rect 9823 7760 13040 7773
rect 9823 7738 10152 7760
rect 7500 7708 7936 7738
rect 7988 7708 8002 7738
rect 8054 7708 8490 7738
rect 8542 7708 8556 7738
rect 8608 7708 9044 7738
rect 9096 7708 9110 7738
rect 9162 7708 9598 7738
rect 9650 7708 9664 7738
rect 9716 7708 10152 7738
rect 10204 7708 10218 7760
rect 10270 7708 10706 7760
rect 10758 7708 10772 7760
rect 10824 7708 11260 7760
rect 11312 7708 11326 7760
rect 11378 7708 11814 7760
rect 11866 7708 11880 7760
rect 11932 7759 13040 7760
rect 11932 7708 12368 7759
rect 2950 7707 12368 7708
rect 12420 7707 12434 7759
rect 12486 7707 12922 7759
rect 12974 7707 12988 7759
rect 2950 7706 13040 7707
rect 2950 7694 7691 7706
rect 3002 7642 3016 7694
rect 3068 7642 3504 7694
rect 3556 7642 3570 7694
rect 3622 7642 4058 7694
rect 4110 7642 4124 7694
rect 4176 7642 4612 7694
rect 4664 7642 4678 7694
rect 4730 7642 5166 7694
rect 5218 7642 5232 7694
rect 5284 7642 5720 7694
rect 5772 7642 5786 7694
rect 5838 7642 6274 7694
rect 6326 7642 6340 7694
rect 6392 7642 6828 7694
rect 6880 7642 6894 7694
rect 6946 7642 7382 7694
rect 7434 7642 7448 7694
rect 7500 7650 7691 7694
rect 7747 7650 7775 7706
rect 7831 7650 7858 7706
rect 7914 7694 7941 7706
rect 7997 7694 8024 7706
rect 7914 7650 7936 7694
rect 7997 7650 8002 7694
rect 8080 7650 8107 7706
rect 8163 7650 8190 7706
rect 8246 7650 8273 7706
rect 8329 7650 8356 7706
rect 8412 7650 8439 7706
rect 8495 7694 8522 7706
rect 8578 7694 8605 7706
rect 8661 7650 8688 7706
rect 8744 7650 8771 7706
rect 8827 7650 8854 7706
rect 8910 7650 8937 7706
rect 8993 7650 9020 7706
rect 9076 7694 9103 7706
rect 9159 7694 9186 7706
rect 9096 7650 9103 7694
rect 9162 7650 9186 7694
rect 9242 7650 9269 7706
rect 9325 7650 9352 7706
rect 9408 7650 9435 7706
rect 9491 7650 9518 7706
rect 9574 7694 9601 7706
rect 9657 7694 9684 7706
rect 9574 7650 9598 7694
rect 9657 7650 9664 7694
rect 9740 7650 9767 7706
rect 9823 7694 13040 7706
rect 9823 7650 10152 7694
rect 7500 7642 7936 7650
rect 7988 7642 8002 7650
rect 8054 7642 8490 7650
rect 8542 7642 8556 7650
rect 8608 7642 9044 7650
rect 9096 7642 9110 7650
rect 9162 7642 9598 7650
rect 9650 7642 9664 7650
rect 9716 7642 10152 7650
rect 10204 7642 10218 7694
rect 10270 7642 10706 7694
rect 10758 7642 10772 7694
rect 10824 7642 11260 7694
rect 11312 7642 11326 7694
rect 11378 7642 11814 7694
rect 11866 7642 11880 7694
rect 11932 7693 13040 7694
rect 11932 7642 12368 7693
rect 2950 7641 12368 7642
rect 12420 7641 12434 7693
rect 12486 7641 12922 7693
rect 12974 7641 12988 7693
rect 2950 7628 13040 7641
rect 3002 7576 3016 7628
rect 3068 7576 3504 7628
rect 3556 7576 3570 7628
rect 3622 7576 4058 7628
rect 4110 7576 4124 7628
rect 4176 7576 4612 7628
rect 4664 7576 4678 7628
rect 4730 7576 5166 7628
rect 5218 7576 5232 7628
rect 5284 7576 5720 7628
rect 5772 7576 5786 7628
rect 5838 7576 6274 7628
rect 6326 7576 6340 7628
rect 6392 7576 6828 7628
rect 6880 7576 6894 7628
rect 6946 7576 7382 7628
rect 7434 7576 7448 7628
rect 7500 7618 7936 7628
rect 7988 7618 8002 7628
rect 8054 7618 8490 7628
rect 8542 7618 8556 7628
rect 8608 7618 9044 7628
rect 9096 7618 9110 7628
rect 9162 7618 9598 7628
rect 9650 7618 9664 7628
rect 9716 7618 10152 7628
rect 7500 7576 7691 7618
rect 2950 7562 7691 7576
rect 7747 7562 7775 7618
rect 7831 7562 7858 7618
rect 7914 7576 7936 7618
rect 7997 7576 8002 7618
rect 7914 7562 7941 7576
rect 7997 7562 8024 7576
rect 8080 7562 8107 7618
rect 8163 7562 8190 7618
rect 8246 7562 8273 7618
rect 8329 7562 8356 7618
rect 8412 7562 8439 7618
rect 8495 7562 8522 7576
rect 8578 7562 8605 7576
rect 8661 7562 8688 7618
rect 8744 7562 8771 7618
rect 8827 7562 8854 7618
rect 8910 7562 8937 7618
rect 8993 7562 9020 7618
rect 9096 7576 9103 7618
rect 9162 7576 9186 7618
rect 9076 7562 9103 7576
rect 9159 7562 9186 7576
rect 9242 7562 9269 7618
rect 9325 7562 9352 7618
rect 9408 7562 9435 7618
rect 9491 7562 9518 7618
rect 9574 7576 9598 7618
rect 9657 7576 9664 7618
rect 9574 7562 9601 7576
rect 9657 7562 9684 7576
rect 9740 7562 9767 7618
rect 9823 7576 10152 7618
rect 10204 7576 10218 7628
rect 10270 7576 10706 7628
rect 10758 7576 10772 7628
rect 10824 7576 11260 7628
rect 11312 7576 11326 7628
rect 11378 7576 11814 7628
rect 11866 7576 11880 7628
rect 11932 7627 13040 7628
rect 11932 7576 12368 7627
rect 9823 7575 12368 7576
rect 12420 7575 12434 7627
rect 12486 7575 12922 7627
rect 12974 7575 12988 7627
rect 9823 7562 13040 7575
rect 3002 7510 3016 7562
rect 3068 7510 3504 7562
rect 3556 7510 3570 7562
rect 3622 7510 4058 7562
rect 4110 7510 4124 7562
rect 4176 7510 4612 7562
rect 4664 7510 4678 7562
rect 4730 7510 5166 7562
rect 5218 7510 5232 7562
rect 5284 7510 5720 7562
rect 5772 7510 5786 7562
rect 5838 7510 6274 7562
rect 6326 7510 6340 7562
rect 6392 7510 6828 7562
rect 6880 7510 6894 7562
rect 6946 7510 7382 7562
rect 7434 7510 7448 7562
rect 7500 7530 7936 7562
rect 7988 7530 8002 7562
rect 8054 7530 8490 7562
rect 8542 7530 8556 7562
rect 8608 7530 9044 7562
rect 9096 7530 9110 7562
rect 9162 7530 9598 7562
rect 9650 7530 9664 7562
rect 9716 7530 10152 7562
rect 7500 7510 7691 7530
rect 2950 7495 7691 7510
rect 3002 7443 3016 7495
rect 3068 7443 3504 7495
rect 3556 7443 3570 7495
rect 3622 7443 4058 7495
rect 4110 7443 4124 7495
rect 4176 7443 4612 7495
rect 4664 7443 4678 7495
rect 4730 7443 5166 7495
rect 5218 7443 5232 7495
rect 5284 7443 5720 7495
rect 5772 7443 5786 7495
rect 5838 7443 6274 7495
rect 6326 7443 6340 7495
rect 6392 7443 6828 7495
rect 6880 7443 6894 7495
rect 6946 7443 7382 7495
rect 7434 7443 7448 7495
rect 7500 7474 7691 7495
rect 7747 7474 7775 7530
rect 7831 7474 7858 7530
rect 7914 7510 7936 7530
rect 7997 7510 8002 7530
rect 7914 7495 7941 7510
rect 7997 7495 8024 7510
rect 7914 7474 7936 7495
rect 7997 7474 8002 7495
rect 8080 7474 8107 7530
rect 8163 7474 8190 7530
rect 8246 7474 8273 7530
rect 8329 7474 8356 7530
rect 8412 7474 8439 7530
rect 8495 7495 8522 7510
rect 8578 7495 8605 7510
rect 8661 7474 8688 7530
rect 8744 7474 8771 7530
rect 8827 7474 8854 7530
rect 8910 7474 8937 7530
rect 8993 7474 9020 7530
rect 9096 7510 9103 7530
rect 9162 7510 9186 7530
rect 9076 7495 9103 7510
rect 9159 7495 9186 7510
rect 9096 7474 9103 7495
rect 9162 7474 9186 7495
rect 9242 7474 9269 7530
rect 9325 7474 9352 7530
rect 9408 7474 9435 7530
rect 9491 7474 9518 7530
rect 9574 7510 9598 7530
rect 9657 7510 9664 7530
rect 9574 7495 9601 7510
rect 9657 7495 9684 7510
rect 9574 7474 9598 7495
rect 9657 7474 9664 7495
rect 9740 7474 9767 7530
rect 9823 7510 10152 7530
rect 10204 7510 10218 7562
rect 10270 7510 10706 7562
rect 10758 7510 10772 7562
rect 10824 7510 11260 7562
rect 11312 7510 11326 7562
rect 11378 7510 11814 7562
rect 11866 7510 11880 7562
rect 11932 7561 13040 7562
rect 11932 7510 12368 7561
rect 9823 7509 12368 7510
rect 12420 7509 12434 7561
rect 12486 7509 12922 7561
rect 12974 7509 12988 7561
rect 9823 7495 13040 7509
rect 9823 7474 10152 7495
rect 7500 7443 7936 7474
rect 7988 7443 8002 7474
rect 8054 7443 8490 7474
rect 8542 7443 8556 7474
rect 8608 7443 9044 7474
rect 9096 7443 9110 7474
rect 9162 7443 9598 7474
rect 9650 7443 9664 7474
rect 9716 7443 10152 7474
rect 10204 7443 10218 7495
rect 10270 7443 10706 7495
rect 10758 7443 10772 7495
rect 10824 7443 11260 7495
rect 11312 7443 11326 7495
rect 11378 7443 11814 7495
rect 11866 7443 11880 7495
rect 11932 7494 13040 7495
rect 11932 7443 12368 7494
rect 2950 7442 12368 7443
rect 12420 7442 12434 7494
rect 12486 7442 12922 7494
rect 12974 7442 12988 7494
rect 2950 7428 7691 7442
rect 3002 7376 3016 7428
rect 3068 7376 3504 7428
rect 3556 7376 3570 7428
rect 3622 7376 4058 7428
rect 4110 7376 4124 7428
rect 4176 7376 4612 7428
rect 4664 7376 4678 7428
rect 4730 7376 5166 7428
rect 5218 7376 5232 7428
rect 5284 7376 5720 7428
rect 5772 7376 5786 7428
rect 5838 7376 6274 7428
rect 6326 7376 6340 7428
rect 6392 7376 6828 7428
rect 6880 7376 6894 7428
rect 6946 7376 7382 7428
rect 7434 7376 7448 7428
rect 7500 7386 7691 7428
rect 7747 7386 7775 7442
rect 7831 7386 7858 7442
rect 7914 7428 7941 7442
rect 7997 7428 8024 7442
rect 7914 7386 7936 7428
rect 7997 7386 8002 7428
rect 8080 7386 8107 7442
rect 8163 7386 8190 7442
rect 8246 7386 8273 7442
rect 8329 7386 8356 7442
rect 8412 7386 8439 7442
rect 8495 7428 8522 7442
rect 8578 7428 8605 7442
rect 8661 7386 8688 7442
rect 8744 7386 8771 7442
rect 8827 7386 8854 7442
rect 8910 7386 8937 7442
rect 8993 7386 9020 7442
rect 9076 7428 9103 7442
rect 9159 7428 9186 7442
rect 9096 7386 9103 7428
rect 9162 7386 9186 7428
rect 9242 7386 9269 7442
rect 9325 7386 9352 7442
rect 9408 7386 9435 7442
rect 9491 7386 9518 7442
rect 9574 7428 9601 7442
rect 9657 7428 9684 7442
rect 9574 7386 9598 7428
rect 9657 7386 9664 7428
rect 9740 7386 9767 7442
rect 9823 7428 13040 7442
rect 9823 7386 10152 7428
rect 7500 7376 7936 7386
rect 7988 7376 8002 7386
rect 8054 7376 8490 7386
rect 8542 7376 8556 7386
rect 8608 7376 9044 7386
rect 9096 7376 9110 7386
rect 9162 7376 9598 7386
rect 9650 7376 9664 7386
rect 9716 7376 10152 7386
rect 10204 7376 10218 7428
rect 10270 7376 10706 7428
rect 10758 7376 10772 7428
rect 10824 7376 11260 7428
rect 11312 7376 11326 7428
rect 11378 7376 11814 7428
rect 11866 7376 11880 7428
rect 11932 7427 13040 7428
rect 11932 7376 12368 7427
rect 2950 7375 12368 7376
rect 12420 7375 12434 7427
rect 12486 7375 12922 7427
rect 12974 7375 12988 7427
rect 2950 7368 13040 7375
rect 13252 7878 13270 7930
rect 13322 7878 13340 7930
rect 13392 7878 13410 7930
rect 13462 7878 13480 7930
rect 13532 7878 13550 7930
rect 13602 7878 14940 7930
rect 13200 7866 14940 7878
rect 13252 7814 13270 7866
rect 13322 7814 13340 7866
rect 13392 7814 13410 7866
rect 13462 7814 13480 7866
rect 13532 7814 13550 7866
rect 13602 7814 14940 7866
rect 13200 7802 14940 7814
rect 13252 7750 13270 7802
rect 13322 7750 13340 7802
rect 13392 7750 13410 7802
rect 13462 7750 13480 7802
rect 13532 7750 13550 7802
rect 13602 7750 14940 7802
rect 13200 7738 14940 7750
rect 13252 7686 13270 7738
rect 13322 7686 13340 7738
rect 13392 7686 13410 7738
rect 13462 7686 13480 7738
rect 13532 7686 13550 7738
rect 13602 7686 14940 7738
rect 13200 7674 14940 7686
rect 13252 7622 13270 7674
rect 13322 7622 13340 7674
rect 13392 7622 13410 7674
rect 13462 7622 13480 7674
rect 13532 7622 13550 7674
rect 13602 7622 14940 7674
rect 13200 7610 14940 7622
rect 13252 7558 13270 7610
rect 13322 7558 13340 7610
rect 13392 7558 13410 7610
rect 13462 7558 13480 7610
rect 13532 7558 13550 7610
rect 13602 7558 14940 7610
rect 13200 7546 14940 7558
rect 13252 7494 13270 7546
rect 13322 7494 13340 7546
rect 13392 7494 13410 7546
rect 13462 7494 13480 7546
rect 13532 7494 13550 7546
rect 13602 7494 14940 7546
rect 13200 7482 14940 7494
rect 13252 7430 13270 7482
rect 13322 7430 13340 7482
rect 13392 7430 13410 7482
rect 13462 7430 13480 7482
rect 13532 7430 13550 7482
rect 13602 7430 14940 7482
rect 13200 7418 14940 7430
rect 13252 7366 13270 7418
rect 13322 7366 13340 7418
rect 13392 7366 13410 7418
rect 13462 7366 13480 7418
rect 13532 7366 13550 7418
rect 13602 7366 14940 7418
rect 13200 7354 14940 7366
rect 13252 7302 13270 7354
rect 13322 7302 13340 7354
rect 13392 7302 13410 7354
rect 13462 7302 13480 7354
rect 13532 7302 13550 7354
rect 13602 7302 14940 7354
rect 13200 7290 14940 7302
rect 13252 7238 13270 7290
rect 13322 7238 13340 7290
rect 13392 7238 13410 7290
rect 13462 7238 13480 7290
rect 13532 7238 13550 7290
rect 13602 7238 14940 7290
rect 13200 7226 14940 7238
rect 13252 7174 13270 7226
rect 13322 7174 13340 7226
rect 13392 7174 13410 7226
rect 13462 7174 13480 7226
rect 13532 7174 13550 7226
rect 13602 7174 14940 7226
rect 13200 7162 14940 7174
rect 13252 7110 13270 7162
rect 13322 7110 13340 7162
rect 13392 7110 13410 7162
rect 13462 7110 13480 7162
rect 13532 7110 13550 7162
rect 13602 7110 14940 7162
rect 13200 7098 14940 7110
rect 13252 7046 13270 7098
rect 13322 7046 13340 7098
rect 13392 7046 13410 7098
rect 13462 7046 13480 7098
rect 13532 7046 13550 7098
rect 13602 7046 14940 7098
rect 13200 7034 14940 7046
rect 13252 6982 13270 7034
rect 13322 6982 13340 7034
rect 13392 6982 13410 7034
rect 13462 6982 13480 7034
rect 13532 6982 13550 7034
rect 13602 6982 14940 7034
rect 13200 6970 14940 6982
tri 13180 6918 13200 6938 se
rect 13252 6918 13270 6970
rect 13322 6918 13340 6970
rect 13392 6918 13410 6970
rect 13462 6918 13480 6970
rect 13532 6918 13550 6970
rect 13602 6918 14940 6970
tri 13168 6906 13180 6918 se
rect 13180 6906 14940 6918
tri 13116 6854 13168 6906 se
rect 13168 6854 13200 6906
rect 13252 6854 13270 6906
rect 13322 6854 13340 6906
rect 13392 6854 13410 6906
rect 13462 6854 13480 6906
rect 13532 6854 13550 6906
rect 13602 6854 14940 6906
tri 13104 6842 13116 6854 se
rect 13116 6842 14940 6854
tri 13052 6790 13104 6842 se
rect 13104 6790 13200 6842
rect 13252 6790 13270 6842
rect 13322 6790 13340 6842
rect 13392 6790 13410 6842
rect 13462 6790 13480 6842
rect 13532 6790 13550 6842
rect 13602 6790 14940 6842
tri 13040 6778 13052 6790 se
rect 13052 6778 14940 6790
tri 12992 6730 13040 6778 se
rect 13040 6730 13200 6778
rect 3227 6726 13200 6730
rect 13252 6726 13270 6778
rect 13322 6726 13340 6778
rect 13392 6726 13410 6778
rect 13462 6726 13480 6778
rect 13532 6726 13550 6778
rect 13602 6726 14940 6778
rect 3227 6724 14940 6726
rect 3279 6672 3293 6724
rect 3345 6672 3781 6724
rect 3833 6672 3847 6724
rect 3899 6672 4335 6724
rect 4387 6672 4401 6724
rect 4453 6672 4889 6724
rect 4941 6672 4955 6724
rect 5007 6672 5443 6724
rect 5495 6672 5509 6724
rect 5561 6672 5997 6724
rect 6049 6672 6063 6724
rect 6115 6672 6551 6724
rect 6603 6672 6617 6724
rect 6669 6672 7105 6724
rect 7157 6672 7171 6724
rect 7223 6672 7659 6724
rect 7711 6672 7725 6724
rect 7777 6672 8213 6724
rect 8265 6672 8279 6724
rect 8331 6672 8767 6724
rect 8819 6672 8833 6724
rect 8885 6672 9321 6724
rect 9373 6672 9387 6724
rect 9439 6672 9875 6724
rect 9927 6672 9941 6724
rect 9993 6672 10429 6724
rect 10481 6672 10495 6724
rect 10547 6672 10983 6724
rect 11035 6672 11049 6724
rect 11101 6672 11537 6724
rect 11589 6672 11603 6724
rect 11655 6672 12091 6724
rect 12143 6672 12157 6724
rect 12209 6672 12645 6724
rect 12697 6672 12711 6724
rect 12763 6714 14940 6724
rect 12763 6672 13200 6714
rect 3227 6662 13200 6672
rect 13252 6662 13270 6714
rect 13322 6662 13340 6714
rect 13392 6662 13410 6714
rect 13462 6662 13480 6714
rect 13532 6662 13550 6714
rect 13602 6662 14940 6714
rect 3227 6658 14940 6662
rect 3279 6606 3293 6658
rect 3345 6606 3781 6658
rect 3833 6606 3847 6658
rect 3899 6606 4335 6658
rect 4387 6606 4401 6658
rect 4453 6606 4889 6658
rect 4941 6606 4955 6658
rect 5007 6606 5443 6658
rect 5495 6606 5509 6658
rect 5561 6606 5997 6658
rect 6049 6606 6063 6658
rect 6115 6606 6551 6658
rect 6603 6606 6617 6658
rect 6669 6606 7105 6658
rect 7157 6606 7171 6658
rect 7223 6606 7659 6658
rect 7711 6606 7725 6658
rect 7777 6606 8213 6658
rect 8265 6606 8279 6658
rect 8331 6606 8767 6658
rect 8819 6606 8833 6658
rect 8885 6606 9321 6658
rect 9373 6606 9387 6658
rect 9439 6606 9875 6658
rect 9927 6606 9941 6658
rect 9993 6606 10429 6658
rect 10481 6606 10495 6658
rect 10547 6606 10983 6658
rect 11035 6606 11049 6658
rect 11101 6606 11537 6658
rect 11589 6606 11603 6658
rect 11655 6606 12091 6658
rect 12143 6606 12157 6658
rect 12209 6606 12645 6658
rect 12697 6606 12711 6658
rect 12763 6650 14940 6658
rect 12763 6606 13200 6650
rect 3227 6598 13200 6606
rect 13252 6598 13270 6650
rect 13322 6598 13340 6650
rect 13392 6598 13410 6650
rect 13462 6598 13480 6650
rect 13532 6598 13550 6650
rect 13602 6598 14940 6650
rect 3227 6592 14940 6598
rect 3279 6540 3293 6592
rect 3345 6540 3781 6592
rect 3833 6540 3847 6592
rect 3899 6540 4335 6592
rect 4387 6540 4401 6592
rect 4453 6540 4889 6592
rect 4941 6540 4955 6592
rect 5007 6540 5443 6592
rect 5495 6540 5509 6592
rect 5561 6540 5997 6592
rect 6049 6540 6063 6592
rect 6115 6540 6551 6592
rect 6603 6540 6617 6592
rect 6669 6540 7105 6592
rect 7157 6540 7171 6592
rect 7223 6540 7659 6592
rect 7711 6540 7725 6592
rect 7777 6540 8213 6592
rect 8265 6540 8279 6592
rect 8331 6540 8767 6592
rect 8819 6540 8833 6592
rect 8885 6540 9321 6592
rect 9373 6540 9387 6592
rect 9439 6540 9875 6592
rect 9927 6540 9941 6592
rect 9993 6540 10429 6592
rect 10481 6540 10495 6592
rect 10547 6540 10983 6592
rect 11035 6540 11049 6592
rect 11101 6540 11537 6592
rect 11589 6540 11603 6592
rect 11655 6540 12091 6592
rect 12143 6540 12157 6592
rect 12209 6540 12645 6592
rect 12697 6540 12711 6592
rect 12763 6586 14940 6592
rect 12763 6540 13200 6586
rect 3227 6534 13200 6540
rect 13252 6534 13270 6586
rect 13322 6534 13340 6586
rect 13392 6534 13410 6586
rect 13462 6534 13480 6586
rect 13532 6534 13550 6586
rect 13602 6534 14940 6586
rect 3227 6526 14940 6534
rect 3279 6474 3293 6526
rect 3345 6474 3781 6526
rect 3833 6474 3847 6526
rect 3899 6474 4335 6526
rect 4387 6474 4401 6526
rect 4453 6474 4889 6526
rect 4941 6474 4955 6526
rect 5007 6474 5443 6526
rect 5495 6474 5509 6526
rect 5561 6474 5997 6526
rect 6049 6474 6063 6526
rect 6115 6474 6551 6526
rect 6603 6474 6617 6526
rect 6669 6474 7105 6526
rect 7157 6474 7171 6526
rect 7223 6474 7659 6526
rect 7711 6474 7725 6526
rect 7777 6474 8213 6526
rect 8265 6474 8279 6526
rect 8331 6474 8767 6526
rect 8819 6474 8833 6526
rect 8885 6474 9321 6526
rect 9373 6474 9387 6526
rect 9439 6474 9875 6526
rect 9927 6474 9941 6526
rect 9993 6474 10429 6526
rect 10481 6474 10495 6526
rect 10547 6474 10983 6526
rect 11035 6474 11049 6526
rect 11101 6474 11537 6526
rect 11589 6474 11603 6526
rect 11655 6474 12091 6526
rect 12143 6474 12157 6526
rect 12209 6474 12645 6526
rect 12697 6474 12711 6526
rect 12763 6522 14940 6526
rect 12763 6474 13200 6522
rect 3227 6470 13200 6474
rect 13252 6470 13270 6522
rect 13322 6470 13340 6522
rect 13392 6470 13410 6522
rect 13462 6470 13480 6522
rect 13532 6470 13550 6522
rect 13602 6470 14940 6522
rect 3227 6460 14940 6470
rect 3279 6408 3293 6460
rect 3345 6408 3781 6460
rect 3833 6408 3847 6460
rect 3899 6408 4335 6460
rect 4387 6408 4401 6460
rect 4453 6408 4889 6460
rect 4941 6408 4955 6460
rect 5007 6408 5443 6460
rect 5495 6408 5509 6460
rect 5561 6408 5997 6460
rect 6049 6408 6063 6460
rect 6115 6408 6551 6460
rect 6603 6408 6617 6460
rect 6669 6408 7105 6460
rect 7157 6408 7171 6460
rect 7223 6408 7659 6460
rect 7711 6408 7725 6460
rect 7777 6408 8213 6460
rect 8265 6408 8279 6460
rect 8331 6408 8767 6460
rect 8819 6408 8833 6460
rect 8885 6408 9321 6460
rect 9373 6408 9387 6460
rect 9439 6408 9875 6460
rect 9927 6408 9941 6460
rect 9993 6408 10429 6460
rect 10481 6408 10495 6460
rect 10547 6408 10983 6460
rect 11035 6408 11049 6460
rect 11101 6408 11537 6460
rect 11589 6408 11603 6460
rect 11655 6408 12091 6460
rect 12143 6408 12157 6460
rect 12209 6408 12645 6460
rect 12697 6408 12711 6460
rect 12763 6458 14940 6460
rect 12763 6408 13200 6458
rect 3227 6406 13200 6408
rect 13252 6406 13270 6458
rect 13322 6406 13340 6458
rect 13392 6406 13410 6458
rect 13462 6406 13480 6458
rect 13532 6406 13550 6458
rect 13602 6406 14940 6458
rect 3227 6394 14940 6406
rect 3279 6342 3293 6394
rect 3345 6342 3781 6394
rect 3833 6342 3847 6394
rect 3899 6342 4335 6394
rect 4387 6342 4401 6394
rect 4453 6342 4889 6394
rect 4941 6342 4955 6394
rect 5007 6342 5443 6394
rect 5495 6342 5509 6394
rect 5561 6342 5997 6394
rect 6049 6342 6063 6394
rect 6115 6342 6551 6394
rect 6603 6342 6617 6394
rect 6669 6342 7105 6394
rect 7157 6342 7171 6394
rect 7223 6342 7659 6394
rect 7711 6342 7725 6394
rect 7777 6342 8213 6394
rect 8265 6342 8279 6394
rect 8331 6342 8767 6394
rect 8819 6342 8833 6394
rect 8885 6342 9321 6394
rect 9373 6342 9387 6394
rect 9439 6342 9875 6394
rect 9927 6342 9941 6394
rect 9993 6342 10429 6394
rect 10481 6342 10495 6394
rect 10547 6342 10983 6394
rect 11035 6342 11049 6394
rect 11101 6342 11537 6394
rect 11589 6342 11603 6394
rect 11655 6342 12091 6394
rect 12143 6342 12157 6394
rect 12209 6342 12645 6394
rect 12697 6342 12711 6394
rect 12763 6342 13200 6394
rect 13252 6342 13270 6394
rect 13322 6342 13340 6394
rect 13392 6342 13410 6394
rect 13462 6342 13480 6394
rect 13532 6342 13550 6394
rect 13602 6342 14940 6394
rect 3227 6330 14940 6342
rect 3227 6327 13200 6330
rect 3279 6275 3293 6327
rect 3345 6275 3781 6327
rect 3833 6275 3847 6327
rect 3899 6275 4335 6327
rect 4387 6275 4401 6327
rect 4453 6275 4889 6327
rect 4941 6275 4955 6327
rect 5007 6275 5443 6327
rect 5495 6275 5509 6327
rect 5561 6275 5997 6327
rect 6049 6275 6063 6327
rect 6115 6275 6551 6327
rect 6603 6275 6617 6327
rect 6669 6275 7105 6327
rect 7157 6275 7171 6327
rect 7223 6275 7659 6327
rect 7711 6275 7725 6327
rect 7777 6275 8213 6327
rect 8265 6275 8279 6327
rect 8331 6275 8767 6327
rect 8819 6275 8833 6327
rect 8885 6275 9321 6327
rect 9373 6275 9387 6327
rect 9439 6275 9875 6327
rect 9927 6275 9941 6327
rect 9993 6275 10429 6327
rect 10481 6275 10495 6327
rect 10547 6275 10983 6327
rect 11035 6275 11049 6327
rect 11101 6275 11537 6327
rect 11589 6275 11603 6327
rect 11655 6275 12091 6327
rect 12143 6275 12157 6327
rect 12209 6275 12645 6327
rect 12697 6275 12711 6327
rect 12763 6278 13200 6327
rect 13252 6278 13270 6330
rect 13322 6278 13340 6330
rect 13392 6278 13410 6330
rect 13462 6278 13480 6330
rect 13532 6278 13550 6330
rect 13602 6278 14940 6330
rect 12763 6275 14940 6278
rect 3227 6266 14940 6275
rect 3227 6260 13200 6266
rect 3279 6208 3293 6260
rect 3345 6208 3781 6260
rect 3833 6208 3847 6260
rect 3899 6208 4335 6260
rect 4387 6208 4401 6260
rect 4453 6208 4889 6260
rect 4941 6208 4955 6260
rect 5007 6208 5443 6260
rect 5495 6208 5509 6260
rect 5561 6208 5997 6260
rect 6049 6208 6063 6260
rect 6115 6208 6551 6260
rect 6603 6208 6617 6260
rect 6669 6208 7105 6260
rect 7157 6208 7171 6260
rect 7223 6208 7659 6260
rect 7711 6208 7725 6260
rect 7777 6208 8213 6260
rect 8265 6208 8279 6260
rect 8331 6208 8767 6260
rect 8819 6208 8833 6260
rect 8885 6208 9321 6260
rect 9373 6208 9387 6260
rect 9439 6208 9875 6260
rect 9927 6208 9941 6260
rect 9993 6208 10429 6260
rect 10481 6208 10495 6260
rect 10547 6208 10983 6260
rect 11035 6208 11049 6260
rect 11101 6208 11537 6260
rect 11589 6208 11603 6260
rect 11655 6208 12091 6260
rect 12143 6208 12157 6260
rect 12209 6208 12645 6260
rect 12697 6208 12711 6260
rect 12763 6214 13200 6260
rect 13252 6214 13270 6266
rect 13322 6214 13340 6266
rect 13392 6214 13410 6266
rect 13462 6214 13480 6266
rect 13532 6214 13550 6266
rect 13602 6214 14940 6266
rect 12763 6208 14940 6214
rect 3227 6202 14940 6208
tri 12974 6150 13026 6202 ne
rect 13026 6150 13200 6202
rect 13252 6150 13270 6202
rect 13322 6150 13340 6202
rect 13392 6150 13410 6202
rect 13462 6150 13480 6202
rect 13532 6150 13550 6202
rect 13602 6150 14940 6202
tri 13026 6138 13038 6150 ne
rect 13038 6138 14940 6150
tri 13038 6086 13090 6138 ne
rect 13090 6086 13200 6138
rect 13252 6086 13270 6138
rect 13322 6086 13340 6138
rect 13392 6086 13410 6138
rect 13462 6086 13480 6138
rect 13532 6086 13550 6138
rect 13602 6086 14940 6138
tri 13090 6074 13102 6086 ne
rect 13102 6074 14940 6086
tri 13102 6022 13154 6074 ne
rect 13154 6022 13200 6074
rect 13252 6022 13270 6074
rect 13322 6022 13340 6074
rect 13392 6022 13410 6074
rect 13462 6022 13480 6074
rect 13532 6022 13550 6074
rect 13602 6022 14940 6074
tri 13154 6010 13166 6022 ne
rect 13166 6010 14940 6022
tri 13166 5976 13200 6010 ne
rect 13252 5958 13270 6010
rect 13322 5958 13340 6010
rect 13392 5958 13410 6010
rect 13462 5958 13480 6010
rect 13532 5958 13550 6010
rect 13602 5958 14940 6010
rect 13200 5946 14940 5958
rect 2950 5896 13040 5902
rect 3002 5844 3016 5896
rect 3068 5844 3504 5896
rect 3556 5844 3570 5896
rect 3622 5844 4058 5896
rect 4110 5844 4124 5896
rect 4176 5844 4612 5896
rect 4664 5844 4678 5896
rect 4730 5844 5166 5896
rect 5218 5844 5232 5896
rect 5284 5844 5720 5896
rect 5772 5844 5786 5896
rect 5838 5844 6274 5896
rect 6326 5844 6340 5896
rect 6392 5844 6828 5896
rect 6880 5844 6894 5896
rect 6946 5844 7382 5896
rect 7434 5844 7448 5896
rect 7500 5877 7936 5896
rect 7988 5877 8002 5896
rect 8054 5877 8490 5896
rect 8542 5877 8556 5896
rect 8608 5877 9044 5896
rect 9096 5877 9110 5896
rect 9162 5877 9598 5896
rect 9650 5877 9664 5896
rect 9716 5877 10152 5896
rect 7500 5844 7691 5877
rect 2950 5830 7691 5844
rect 3002 5778 3016 5830
rect 3068 5778 3504 5830
rect 3556 5778 3570 5830
rect 3622 5778 4058 5830
rect 4110 5778 4124 5830
rect 4176 5778 4612 5830
rect 4664 5778 4678 5830
rect 4730 5778 5166 5830
rect 5218 5778 5232 5830
rect 5284 5778 5720 5830
rect 5772 5778 5786 5830
rect 5838 5778 6274 5830
rect 6326 5778 6340 5830
rect 6392 5778 6828 5830
rect 6880 5778 6894 5830
rect 6946 5778 7382 5830
rect 7434 5778 7448 5830
rect 7500 5821 7691 5830
rect 7747 5821 7775 5877
rect 7831 5821 7858 5877
rect 7914 5844 7936 5877
rect 7997 5844 8002 5877
rect 7914 5830 7941 5844
rect 7997 5830 8024 5844
rect 7914 5821 7936 5830
rect 7997 5821 8002 5830
rect 8080 5821 8107 5877
rect 8163 5821 8190 5877
rect 8246 5821 8273 5877
rect 8329 5821 8356 5877
rect 8412 5821 8439 5877
rect 8495 5830 8522 5844
rect 8578 5830 8605 5844
rect 8661 5821 8688 5877
rect 8744 5821 8771 5877
rect 8827 5821 8854 5877
rect 8910 5821 8937 5877
rect 8993 5821 9020 5877
rect 9096 5844 9103 5877
rect 9162 5844 9186 5877
rect 9076 5830 9103 5844
rect 9159 5830 9186 5844
rect 9096 5821 9103 5830
rect 9162 5821 9186 5830
rect 9242 5821 9269 5877
rect 9325 5821 9352 5877
rect 9408 5821 9435 5877
rect 9491 5821 9518 5877
rect 9574 5844 9598 5877
rect 9657 5844 9664 5877
rect 9574 5830 9601 5844
rect 9657 5830 9684 5844
rect 9574 5821 9598 5830
rect 9657 5821 9664 5830
rect 9740 5821 9767 5877
rect 9823 5844 10152 5877
rect 10204 5844 10218 5896
rect 10270 5844 10706 5896
rect 10758 5844 10772 5896
rect 10824 5844 11260 5896
rect 11312 5844 11326 5896
rect 11378 5844 11814 5896
rect 11866 5844 11880 5896
rect 11932 5894 13040 5896
rect 11932 5844 12368 5894
rect 9823 5842 12368 5844
rect 12420 5842 12434 5894
rect 12486 5842 12922 5894
rect 12974 5842 12988 5894
rect 9823 5830 13040 5842
rect 9823 5821 10152 5830
rect 7500 5789 7936 5821
rect 7988 5789 8002 5821
rect 8054 5789 8490 5821
rect 8542 5789 8556 5821
rect 8608 5789 9044 5821
rect 9096 5789 9110 5821
rect 9162 5789 9598 5821
rect 9650 5789 9664 5821
rect 9716 5789 10152 5821
rect 7500 5778 7691 5789
rect 2950 5764 7691 5778
rect 3002 5712 3016 5764
rect 3068 5712 3504 5764
rect 3556 5712 3570 5764
rect 3622 5712 4058 5764
rect 4110 5712 4124 5764
rect 4176 5712 4612 5764
rect 4664 5712 4678 5764
rect 4730 5712 5166 5764
rect 5218 5712 5232 5764
rect 5284 5712 5720 5764
rect 5772 5712 5786 5764
rect 5838 5712 6274 5764
rect 6326 5712 6340 5764
rect 6392 5712 6828 5764
rect 6880 5712 6894 5764
rect 6946 5712 7382 5764
rect 7434 5712 7448 5764
rect 7500 5733 7691 5764
rect 7747 5733 7775 5789
rect 7831 5733 7858 5789
rect 7914 5778 7936 5789
rect 7997 5778 8002 5789
rect 7914 5764 7941 5778
rect 7997 5764 8024 5778
rect 7914 5733 7936 5764
rect 7997 5733 8002 5764
rect 8080 5733 8107 5789
rect 8163 5733 8190 5789
rect 8246 5733 8273 5789
rect 8329 5733 8356 5789
rect 8412 5733 8439 5789
rect 8495 5764 8522 5778
rect 8578 5764 8605 5778
rect 8661 5733 8688 5789
rect 8744 5733 8771 5789
rect 8827 5733 8854 5789
rect 8910 5733 8937 5789
rect 8993 5733 9020 5789
rect 9096 5778 9103 5789
rect 9162 5778 9186 5789
rect 9076 5764 9103 5778
rect 9159 5764 9186 5778
rect 9096 5733 9103 5764
rect 9162 5733 9186 5764
rect 9242 5733 9269 5789
rect 9325 5733 9352 5789
rect 9408 5733 9435 5789
rect 9491 5733 9518 5789
rect 9574 5778 9598 5789
rect 9657 5778 9664 5789
rect 9574 5764 9601 5778
rect 9657 5764 9684 5778
rect 9574 5733 9598 5764
rect 9657 5733 9664 5764
rect 9740 5733 9767 5789
rect 9823 5778 10152 5789
rect 10204 5778 10218 5830
rect 10270 5778 10706 5830
rect 10758 5778 10772 5830
rect 10824 5778 11260 5830
rect 11312 5778 11326 5830
rect 11378 5778 11814 5830
rect 11866 5778 11880 5830
rect 11932 5828 13040 5830
rect 11932 5778 12368 5828
rect 9823 5776 12368 5778
rect 12420 5776 12434 5828
rect 12486 5776 12922 5828
rect 12974 5776 12988 5828
rect 9823 5764 13040 5776
rect 9823 5733 10152 5764
rect 7500 5712 7936 5733
rect 7988 5712 8002 5733
rect 8054 5712 8490 5733
rect 8542 5712 8556 5733
rect 8608 5712 9044 5733
rect 9096 5712 9110 5733
rect 9162 5712 9598 5733
rect 9650 5712 9664 5733
rect 9716 5712 10152 5733
rect 10204 5712 10218 5764
rect 10270 5712 10706 5764
rect 10758 5712 10772 5764
rect 10824 5712 11260 5764
rect 11312 5712 11326 5764
rect 11378 5712 11814 5764
rect 11866 5712 11880 5764
rect 11932 5762 13040 5764
rect 11932 5712 12368 5762
rect 2950 5710 12368 5712
rect 12420 5710 12434 5762
rect 12486 5710 12922 5762
rect 12974 5710 12988 5762
rect 2950 5701 13040 5710
rect 2950 5698 7691 5701
rect 3002 5646 3016 5698
rect 3068 5646 3504 5698
rect 3556 5646 3570 5698
rect 3622 5646 4058 5698
rect 4110 5646 4124 5698
rect 4176 5646 4612 5698
rect 4664 5646 4678 5698
rect 4730 5646 5166 5698
rect 5218 5646 5232 5698
rect 5284 5646 5720 5698
rect 5772 5646 5786 5698
rect 5838 5646 6274 5698
rect 6326 5646 6340 5698
rect 6392 5646 6828 5698
rect 6880 5646 6894 5698
rect 6946 5646 7382 5698
rect 7434 5646 7448 5698
rect 7500 5646 7691 5698
rect 2950 5645 7691 5646
rect 7747 5645 7775 5701
rect 7831 5645 7858 5701
rect 7914 5698 7941 5701
rect 7997 5698 8024 5701
rect 7914 5646 7936 5698
rect 7997 5646 8002 5698
rect 7914 5645 7941 5646
rect 7997 5645 8024 5646
rect 8080 5645 8107 5701
rect 8163 5645 8190 5701
rect 8246 5645 8273 5701
rect 8329 5645 8356 5701
rect 8412 5645 8439 5701
rect 8495 5698 8522 5701
rect 8578 5698 8605 5701
rect 8495 5645 8522 5646
rect 8578 5645 8605 5646
rect 8661 5645 8688 5701
rect 8744 5645 8771 5701
rect 8827 5645 8854 5701
rect 8910 5645 8937 5701
rect 8993 5645 9020 5701
rect 9076 5698 9103 5701
rect 9159 5698 9186 5701
rect 9096 5646 9103 5698
rect 9162 5646 9186 5698
rect 9076 5645 9103 5646
rect 9159 5645 9186 5646
rect 9242 5645 9269 5701
rect 9325 5645 9352 5701
rect 9408 5645 9435 5701
rect 9491 5645 9518 5701
rect 9574 5698 9601 5701
rect 9657 5698 9684 5701
rect 9574 5646 9598 5698
rect 9657 5646 9664 5698
rect 9574 5645 9601 5646
rect 9657 5645 9684 5646
rect 9740 5645 9767 5701
rect 9823 5698 13040 5701
rect 9823 5646 10152 5698
rect 10204 5646 10218 5698
rect 10270 5646 10706 5698
rect 10758 5646 10772 5698
rect 10824 5646 11260 5698
rect 11312 5646 11326 5698
rect 11378 5646 11814 5698
rect 11866 5646 11880 5698
rect 11932 5696 13040 5698
rect 11932 5646 12368 5696
rect 9823 5645 12368 5646
rect 2950 5644 12368 5645
rect 12420 5644 12434 5696
rect 12486 5644 12922 5696
rect 12974 5644 12988 5696
rect 2950 5632 13040 5644
rect 3002 5580 3016 5632
rect 3068 5580 3504 5632
rect 3556 5580 3570 5632
rect 3622 5580 4058 5632
rect 4110 5580 4124 5632
rect 4176 5580 4612 5632
rect 4664 5580 4678 5632
rect 4730 5580 5166 5632
rect 5218 5580 5232 5632
rect 5284 5580 5720 5632
rect 5772 5580 5786 5632
rect 5838 5580 6274 5632
rect 6326 5580 6340 5632
rect 6392 5580 6828 5632
rect 6880 5580 6894 5632
rect 6946 5580 7382 5632
rect 7434 5580 7448 5632
rect 7500 5613 7936 5632
rect 7988 5613 8002 5632
rect 8054 5613 8490 5632
rect 8542 5613 8556 5632
rect 8608 5613 9044 5632
rect 9096 5613 9110 5632
rect 9162 5613 9598 5632
rect 9650 5613 9664 5632
rect 9716 5613 10152 5632
rect 7500 5580 7691 5613
rect 2950 5566 7691 5580
rect 3002 5514 3016 5566
rect 3068 5514 3504 5566
rect 3556 5514 3570 5566
rect 3622 5514 4058 5566
rect 4110 5514 4124 5566
rect 4176 5514 4612 5566
rect 4664 5514 4678 5566
rect 4730 5514 5166 5566
rect 5218 5514 5232 5566
rect 5284 5514 5720 5566
rect 5772 5514 5786 5566
rect 5838 5514 6274 5566
rect 6326 5514 6340 5566
rect 6392 5514 6828 5566
rect 6880 5514 6894 5566
rect 6946 5514 7382 5566
rect 7434 5514 7448 5566
rect 7500 5557 7691 5566
rect 7747 5557 7775 5613
rect 7831 5557 7858 5613
rect 7914 5580 7936 5613
rect 7997 5580 8002 5613
rect 7914 5566 7941 5580
rect 7997 5566 8024 5580
rect 7914 5557 7936 5566
rect 7997 5557 8002 5566
rect 8080 5557 8107 5613
rect 8163 5557 8190 5613
rect 8246 5557 8273 5613
rect 8329 5557 8356 5613
rect 8412 5557 8439 5613
rect 8495 5566 8522 5580
rect 8578 5566 8605 5580
rect 8661 5557 8688 5613
rect 8744 5557 8771 5613
rect 8827 5557 8854 5613
rect 8910 5557 8937 5613
rect 8993 5557 9020 5613
rect 9096 5580 9103 5613
rect 9162 5580 9186 5613
rect 9076 5566 9103 5580
rect 9159 5566 9186 5580
rect 9096 5557 9103 5566
rect 9162 5557 9186 5566
rect 9242 5557 9269 5613
rect 9325 5557 9352 5613
rect 9408 5557 9435 5613
rect 9491 5557 9518 5613
rect 9574 5580 9598 5613
rect 9657 5580 9664 5613
rect 9574 5566 9601 5580
rect 9657 5566 9684 5580
rect 9574 5557 9598 5566
rect 9657 5557 9664 5566
rect 9740 5557 9767 5613
rect 9823 5580 10152 5613
rect 10204 5580 10218 5632
rect 10270 5580 10706 5632
rect 10758 5580 10772 5632
rect 10824 5580 11260 5632
rect 11312 5580 11326 5632
rect 11378 5580 11814 5632
rect 11866 5580 11880 5632
rect 11932 5630 13040 5632
rect 11932 5580 12368 5630
rect 9823 5578 12368 5580
rect 12420 5578 12434 5630
rect 12486 5578 12922 5630
rect 12974 5578 12988 5630
rect 9823 5566 13040 5578
rect 9823 5557 10152 5566
rect 7500 5525 7936 5557
rect 7988 5525 8002 5557
rect 8054 5525 8490 5557
rect 8542 5525 8556 5557
rect 8608 5525 9044 5557
rect 9096 5525 9110 5557
rect 9162 5525 9598 5557
rect 9650 5525 9664 5557
rect 9716 5525 10152 5557
rect 7500 5514 7691 5525
rect 2950 5499 7691 5514
rect 3002 5447 3016 5499
rect 3068 5447 3504 5499
rect 3556 5447 3570 5499
rect 3622 5447 4058 5499
rect 4110 5447 4124 5499
rect 4176 5447 4612 5499
rect 4664 5447 4678 5499
rect 4730 5447 5166 5499
rect 5218 5447 5232 5499
rect 5284 5447 5720 5499
rect 5772 5447 5786 5499
rect 5838 5447 6274 5499
rect 6326 5447 6340 5499
rect 6392 5447 6828 5499
rect 6880 5447 6894 5499
rect 6946 5447 7382 5499
rect 7434 5447 7448 5499
rect 7500 5469 7691 5499
rect 7747 5469 7775 5525
rect 7831 5469 7858 5525
rect 7914 5514 7936 5525
rect 7997 5514 8002 5525
rect 7914 5499 7941 5514
rect 7997 5499 8024 5514
rect 7914 5469 7936 5499
rect 7997 5469 8002 5499
rect 8080 5469 8107 5525
rect 8163 5469 8190 5525
rect 8246 5469 8273 5525
rect 8329 5469 8356 5525
rect 8412 5469 8439 5525
rect 8495 5499 8522 5514
rect 8578 5499 8605 5514
rect 8661 5469 8688 5525
rect 8744 5469 8771 5525
rect 8827 5469 8854 5525
rect 8910 5469 8937 5525
rect 8993 5469 9020 5525
rect 9096 5514 9103 5525
rect 9162 5514 9186 5525
rect 9076 5499 9103 5514
rect 9159 5499 9186 5514
rect 9096 5469 9103 5499
rect 9162 5469 9186 5499
rect 9242 5469 9269 5525
rect 9325 5469 9352 5525
rect 9408 5469 9435 5525
rect 9491 5469 9518 5525
rect 9574 5514 9598 5525
rect 9657 5514 9664 5525
rect 9574 5499 9601 5514
rect 9657 5499 9684 5514
rect 9574 5469 9598 5499
rect 9657 5469 9664 5499
rect 9740 5469 9767 5525
rect 9823 5514 10152 5525
rect 10204 5514 10218 5566
rect 10270 5514 10706 5566
rect 10758 5514 10772 5566
rect 10824 5514 11260 5566
rect 11312 5514 11326 5566
rect 11378 5514 11814 5566
rect 11866 5514 11880 5566
rect 11932 5564 13040 5566
rect 11932 5514 12368 5564
rect 9823 5512 12368 5514
rect 12420 5512 12434 5564
rect 12486 5512 12922 5564
rect 12974 5512 12988 5564
rect 9823 5499 13040 5512
rect 9823 5469 10152 5499
rect 7500 5447 7936 5469
rect 7988 5447 8002 5469
rect 8054 5447 8490 5469
rect 8542 5447 8556 5469
rect 8608 5447 9044 5469
rect 9096 5447 9110 5469
rect 9162 5447 9598 5469
rect 9650 5447 9664 5469
rect 9716 5447 10152 5469
rect 10204 5447 10218 5499
rect 10270 5447 10706 5499
rect 10758 5447 10772 5499
rect 10824 5447 11260 5499
rect 11312 5447 11326 5499
rect 11378 5447 11814 5499
rect 11866 5447 11880 5499
rect 11932 5497 13040 5499
rect 11932 5447 12368 5497
rect 2950 5445 12368 5447
rect 12420 5445 12434 5497
rect 12486 5445 12922 5497
rect 12974 5445 12988 5497
rect 2950 5437 13040 5445
rect 2950 5432 7691 5437
rect 3002 5380 3016 5432
rect 3068 5380 3504 5432
rect 3556 5380 3570 5432
rect 3622 5380 4058 5432
rect 4110 5380 4124 5432
rect 4176 5380 4612 5432
rect 4664 5380 4678 5432
rect 4730 5380 5166 5432
rect 5218 5380 5232 5432
rect 5284 5380 5720 5432
rect 5772 5380 5786 5432
rect 5838 5380 6274 5432
rect 6326 5380 6340 5432
rect 6392 5380 6828 5432
rect 6880 5380 6894 5432
rect 6946 5380 7382 5432
rect 7434 5380 7448 5432
rect 7500 5381 7691 5432
rect 7747 5381 7775 5437
rect 7831 5381 7858 5437
rect 7914 5432 7941 5437
rect 7997 5432 8024 5437
rect 7914 5381 7936 5432
rect 7997 5381 8002 5432
rect 8080 5381 8107 5437
rect 8163 5381 8190 5437
rect 8246 5381 8273 5437
rect 8329 5381 8356 5437
rect 8412 5381 8439 5437
rect 8495 5432 8522 5437
rect 8578 5432 8605 5437
rect 8661 5381 8688 5437
rect 8744 5381 8771 5437
rect 8827 5381 8854 5437
rect 8910 5381 8937 5437
rect 8993 5381 9020 5437
rect 9076 5432 9103 5437
rect 9159 5432 9186 5437
rect 9096 5381 9103 5432
rect 9162 5381 9186 5432
rect 9242 5381 9269 5437
rect 9325 5381 9352 5437
rect 9408 5381 9435 5437
rect 9491 5381 9518 5437
rect 9574 5432 9601 5437
rect 9657 5432 9684 5437
rect 9574 5381 9598 5432
rect 9657 5381 9664 5432
rect 9740 5381 9767 5437
rect 9823 5432 13040 5437
rect 9823 5381 10152 5432
rect 7500 5380 7936 5381
rect 7988 5380 8002 5381
rect 8054 5380 8490 5381
rect 8542 5380 8556 5381
rect 8608 5380 9044 5381
rect 9096 5380 9110 5381
rect 9162 5380 9598 5381
rect 9650 5380 9664 5381
rect 9716 5380 10152 5381
rect 10204 5380 10218 5432
rect 10270 5380 10706 5432
rect 10758 5380 10772 5432
rect 10824 5380 11260 5432
rect 11312 5380 11326 5432
rect 11378 5380 11814 5432
rect 11866 5380 11880 5432
rect 11932 5430 13040 5432
rect 11932 5380 12368 5430
rect 2950 5378 12368 5380
rect 12420 5378 12434 5430
rect 12486 5378 12922 5430
rect 12974 5378 12988 5430
rect 2950 5372 13040 5378
rect 13252 5894 13270 5946
rect 13322 5894 13340 5946
rect 13392 5894 13410 5946
rect 13462 5894 13480 5946
rect 13532 5894 13550 5946
rect 13602 5894 14940 5946
rect 13200 5882 14940 5894
rect 13252 5830 13270 5882
rect 13322 5830 13340 5882
rect 13392 5830 13410 5882
rect 13462 5830 13480 5882
rect 13532 5830 13550 5882
rect 13602 5830 14940 5882
rect 13200 5818 14940 5830
rect 13252 5766 13270 5818
rect 13322 5766 13340 5818
rect 13392 5766 13410 5818
rect 13462 5766 13480 5818
rect 13532 5766 13550 5818
rect 13602 5766 14940 5818
rect 13200 5754 14940 5766
rect 13252 5702 13270 5754
rect 13322 5702 13340 5754
rect 13392 5702 13410 5754
rect 13462 5702 13480 5754
rect 13532 5702 13550 5754
rect 13602 5702 14940 5754
rect 13200 5690 14940 5702
rect 13252 5638 13270 5690
rect 13322 5638 13340 5690
rect 13392 5638 13410 5690
rect 13462 5638 13480 5690
rect 13532 5638 13550 5690
rect 13602 5638 14940 5690
rect 13200 5626 14940 5638
rect 13252 5574 13270 5626
rect 13322 5574 13340 5626
rect 13392 5574 13410 5626
rect 13462 5574 13480 5626
rect 13532 5574 13550 5626
rect 13602 5574 14940 5626
rect 13200 5562 14940 5574
rect 13252 5510 13270 5562
rect 13322 5510 13340 5562
rect 13392 5510 13410 5562
rect 13462 5510 13480 5562
rect 13532 5510 13550 5562
rect 13602 5510 14940 5562
rect 13200 5498 14940 5510
rect 13252 5446 13270 5498
rect 13322 5446 13340 5498
rect 13392 5446 13410 5498
rect 13462 5446 13480 5498
rect 13532 5446 13550 5498
rect 13602 5446 14940 5498
rect 13200 5434 14940 5446
rect 13252 5382 13270 5434
rect 13322 5382 13340 5434
rect 13392 5382 13410 5434
rect 13462 5382 13480 5434
rect 13532 5382 13550 5434
rect 13602 5382 14940 5434
rect 13200 5370 14940 5382
rect 13252 5318 13270 5370
rect 13322 5318 13340 5370
rect 13392 5318 13410 5370
rect 13462 5318 13480 5370
rect 13532 5318 13550 5370
rect 13602 5318 14940 5370
rect 13200 5306 14940 5318
rect 13252 5254 13270 5306
rect 13322 5254 13340 5306
rect 13392 5254 13410 5306
rect 13462 5254 13480 5306
rect 13532 5254 13550 5306
rect 13602 5254 14940 5306
rect 13200 5242 14940 5254
rect 5013 5201 6356 5210
rect 5069 5145 6356 5201
rect 5013 5121 6356 5145
rect 5069 5065 6356 5121
rect 13252 5190 13270 5242
rect 13322 5190 13340 5242
rect 13392 5190 13410 5242
rect 13462 5190 13480 5242
rect 13532 5190 13550 5242
rect 13602 5190 14940 5242
rect 13200 5178 14940 5190
rect 13252 5126 13270 5178
rect 13322 5126 13340 5178
rect 13392 5126 13410 5178
rect 13462 5126 13480 5178
rect 13532 5126 13550 5178
rect 13602 5126 14940 5178
rect 13200 5114 14940 5126
rect 5013 5056 6356 5065
tri 13174 5062 13200 5088 se
rect 13252 5062 13270 5114
rect 13322 5062 13340 5114
rect 13392 5062 13410 5114
rect 13462 5062 13480 5114
rect 13532 5062 13550 5114
rect 13602 5062 14940 5114
tri 13168 5056 13174 5062 se
rect 13174 5056 14940 5062
tri 6050 5049 6057 5056 ne
rect 6057 5049 6356 5056
tri 13161 5049 13168 5056 se
rect 13168 5049 14940 5056
tri 6057 5037 6069 5049 ne
rect 6069 5037 6356 5049
tri 2750 4997 2790 5037 sw
tri 6069 4997 6109 5037 ne
rect 6109 4997 6356 5037
tri 13109 4997 13161 5049 se
rect 13161 4997 13200 5049
rect 13252 4997 13270 5049
rect 13322 4997 13340 5049
rect 13392 4997 13410 5049
rect 13462 4997 13480 5049
rect 13532 4997 13550 5049
rect 13602 4997 14940 5049
rect 100 4877 2790 4997
tri 2790 4877 2910 4997 sw
tri 6109 4922 6184 4997 ne
rect 100 4825 2910 4877
tri 2910 4825 2962 4877 sw
rect 4962 4825 4968 4877
rect 5020 4867 5085 4877
rect 5020 4825 5022 4867
rect 100 4811 2962 4825
tri 2962 4811 2976 4825 sw
rect 4962 4811 5022 4825
rect 5078 4825 5085 4867
rect 5137 4825 5202 4877
rect 5254 4825 5260 4877
rect 5078 4811 5260 4825
rect 100 4759 2976 4811
tri 2976 4759 3028 4811 sw
rect 4962 4759 4968 4811
rect 5020 4785 5085 4811
rect 5020 4759 5022 4785
rect 100 4724 3028 4759
tri 3028 4724 3063 4759 sw
tri 4981 4724 5016 4759 ne
rect 5016 4729 5022 4759
rect 5078 4759 5085 4785
rect 5137 4759 5202 4811
rect 5254 4759 5260 4811
rect 5078 4729 5084 4759
rect 100 4721 3063 4724
tri 3063 4721 3066 4724 sw
rect 100 4669 3066 4721
tri 3066 4669 3118 4721 sw
rect 5016 4702 5084 4729
tri 5084 4722 5121 4759 nw
rect 100 4637 3118 4669
tri 3118 4637 3150 4669 sw
rect 5016 4646 5022 4702
rect 5078 4646 5084 4702
rect 5016 4637 5084 4646
rect 100 4635 3150 4637
tri 3150 4635 3152 4637 sw
rect 100 4583 3152 4635
tri 3152 4583 3204 4635 sw
rect 100 4577 3204 4583
tri 3204 4577 3210 4583 sw
rect 100 4339 3210 4577
tri 3210 4339 3448 4577 sw
rect 100 4220 3448 4339
tri 3448 4220 3567 4339 sw
rect 100 4168 3567 4220
tri 3567 4168 3619 4220 sw
rect 5203 4168 5209 4220
rect 5268 4168 5278 4220
rect 5330 4168 5346 4220
rect 5403 4168 5414 4220
rect 5466 4168 5481 4220
rect 5537 4168 5550 4220
rect 5602 4168 5615 4220
rect 5671 4168 5686 4220
rect 5738 4168 5749 4220
rect 5806 4168 5822 4220
rect 5874 4168 5883 4220
rect 5942 4168 5948 4220
rect 100 4096 3619 4168
tri 3619 4096 3691 4168 sw
rect 5203 4164 5212 4168
rect 5268 4164 5347 4168
rect 5403 4164 5481 4168
rect 5537 4164 5615 4168
rect 5671 4164 5749 4168
rect 5805 4164 5883 4168
rect 5939 4164 5948 4168
rect 5203 4100 5948 4164
rect 5203 4096 5212 4100
rect 5268 4096 5347 4100
rect 5403 4096 5481 4100
rect 5537 4096 5615 4100
rect 5671 4096 5749 4100
rect 5805 4096 5883 4100
rect 5939 4096 5948 4100
rect 100 4044 3691 4096
tri 3691 4044 3743 4096 sw
rect 5203 4044 5209 4096
rect 5268 4044 5278 4096
rect 5330 4044 5346 4096
rect 5403 4044 5414 4096
rect 5466 4044 5481 4096
rect 5537 4044 5550 4096
rect 5602 4044 5615 4096
rect 5671 4044 5686 4096
rect 5738 4044 5749 4096
rect 5806 4044 5822 4096
rect 5874 4044 5883 4096
rect 5942 4044 5948 4096
rect 100 3666 3743 4044
tri 3743 3666 4121 4044 sw
tri 6091 3666 6184 3759 se
rect 6184 3666 6356 4997
tri 12989 4877 13109 4997 se
rect 13109 4877 14940 4997
tri 12871 4759 12989 4877 se
rect 12989 4759 14940 4877
tri 12839 4727 12871 4759 se
rect 12871 4727 14940 4759
rect 7676 4724 10501 4727
rect 7676 4668 7692 4724
rect 7748 4668 7853 4724
rect 7909 4668 8014 4724
rect 8070 4668 8175 4724
rect 8231 4668 8336 4724
rect 8392 4668 8497 4724
rect 8553 4668 8658 4724
rect 8714 4668 8819 4724
rect 8875 4668 8980 4724
rect 9036 4668 9141 4724
rect 9197 4668 9302 4724
rect 9358 4668 9462 4724
rect 9518 4668 9622 4724
rect 9678 4668 9782 4724
rect 9838 4721 10501 4724
tri 12834 4722 12839 4727 se
rect 12839 4722 14940 4727
rect 9838 4669 10369 4721
rect 10421 4669 10445 4721
rect 10497 4669 10501 4721
rect 9838 4668 10501 4669
rect 7676 4636 10501 4668
tri 12749 4637 12834 4722 se
rect 12834 4637 14940 4722
rect 7676 4580 7692 4636
rect 7748 4580 7853 4636
rect 7909 4580 8014 4636
rect 8070 4580 8175 4636
rect 8231 4580 8336 4636
rect 8392 4580 8497 4636
rect 8553 4580 8658 4636
rect 8714 4580 8819 4636
rect 8875 4580 8980 4636
rect 9036 4580 9141 4636
rect 9197 4580 9302 4636
rect 9358 4580 9462 4636
rect 9518 4580 9622 4636
rect 9678 4580 9782 4636
rect 9838 4635 10501 4636
rect 9838 4583 10369 4635
rect 10421 4583 10445 4635
rect 10497 4583 10501 4635
rect 9838 4580 10501 4583
rect 7676 4577 10501 4580
tri 12689 4577 12749 4637 se
rect 12749 4577 14940 4637
tri 12451 4339 12689 4577 se
rect 12689 4339 14940 4577
rect 10819 3998 14940 4339
tri 10819 3759 11058 3998 ne
rect 11058 3759 14940 3998
tri 6356 3666 6449 3759 sw
tri 11058 3666 11151 3759 ne
rect 11151 3666 14940 3759
rect 100 3614 4121 3666
tri 4121 3614 4173 3666 sw
rect 4814 3614 4820 3666
rect 4872 3614 4885 3666
rect 4937 3614 4950 3666
rect 5002 3614 5015 3666
rect 5067 3614 5080 3666
rect 5132 3614 5145 3666
rect 5197 3614 5210 3666
rect 5262 3614 5275 3666
rect 5327 3614 5340 3666
rect 5392 3614 5405 3666
rect 5457 3614 5470 3666
rect 5522 3614 5535 3666
rect 5587 3614 5600 3666
rect 5652 3614 5665 3666
rect 5717 3614 5730 3666
rect 5782 3614 5795 3666
rect 5847 3614 5860 3666
rect 5912 3614 5925 3666
rect 5977 3614 5990 3666
rect 6042 3614 6055 3666
rect 6107 3614 6120 3666
rect 6172 3614 6185 3666
rect 6237 3614 6250 3666
rect 6302 3614 6315 3666
rect 6367 3614 6380 3666
rect 6432 3614 6445 3666
rect 6497 3614 6510 3666
rect 6562 3614 6575 3666
rect 6627 3614 6640 3666
rect 6692 3614 6705 3666
rect 6757 3614 6770 3666
rect 6822 3614 6835 3666
rect 6887 3614 6900 3666
rect 6952 3614 6965 3666
rect 7017 3614 7030 3666
rect 7082 3614 7095 3666
rect 7147 3614 7160 3666
rect 7212 3614 7225 3666
rect 7277 3614 7290 3666
rect 7342 3614 7355 3666
rect 7407 3614 7419 3666
rect 7471 3614 7483 3666
rect 7535 3614 7547 3666
rect 7599 3614 7611 3666
rect 7663 3614 7675 3666
rect 7727 3614 7739 3666
rect 7791 3614 7803 3666
rect 7855 3614 7867 3666
rect 7919 3614 7931 3666
rect 7983 3614 7995 3666
rect 8047 3614 8059 3666
rect 8111 3614 8123 3666
rect 8175 3614 8187 3666
rect 8239 3614 8251 3666
rect 8303 3614 8315 3666
rect 8367 3614 8379 3666
rect 8431 3614 8443 3666
rect 8495 3614 8507 3666
rect 8559 3614 8571 3666
rect 8623 3614 8635 3666
rect 8687 3614 8699 3666
rect 8751 3614 8763 3666
rect 8815 3614 8827 3666
rect 8879 3614 8891 3666
rect 8943 3614 8955 3666
rect 9007 3614 9019 3666
rect 9071 3614 9083 3666
rect 9135 3614 9147 3666
rect 9199 3614 9211 3666
rect 9263 3614 9275 3666
rect 9327 3614 9339 3666
rect 9391 3614 9403 3666
rect 9455 3614 9467 3666
rect 9519 3614 9531 3666
rect 9583 3614 9595 3666
rect 9647 3614 9659 3666
rect 9711 3614 9723 3666
rect 9775 3614 9787 3666
rect 9839 3614 9851 3666
rect 9903 3614 9915 3666
rect 9967 3614 9979 3666
rect 10031 3614 10043 3666
rect 10095 3614 10107 3666
rect 10159 3614 10171 3666
rect 10223 3614 10235 3666
rect 10287 3614 10299 3666
rect 10351 3614 10363 3666
rect 10415 3614 10427 3666
rect 10479 3614 10491 3666
rect 10543 3614 10555 3666
rect 10607 3614 10619 3666
rect 10671 3614 10683 3666
rect 10735 3614 10747 3666
rect 10799 3614 10811 3666
rect 10863 3614 10869 3666
rect 100 3578 4173 3614
tri 4173 3578 4209 3614 sw
rect 4814 3578 10869 3614
rect 100 3526 4209 3578
tri 4209 3526 4261 3578 sw
rect 4814 3526 4820 3578
rect 4872 3526 4885 3578
rect 4937 3526 4950 3578
rect 5002 3526 5015 3578
rect 5067 3526 5080 3578
rect 5132 3526 5145 3578
rect 5197 3526 5210 3578
rect 5262 3526 5275 3578
rect 5327 3526 5340 3578
rect 5392 3526 5405 3578
rect 5457 3526 5470 3578
rect 5522 3526 5535 3578
rect 5587 3526 5600 3578
rect 5652 3526 5665 3578
rect 5717 3526 5730 3578
rect 5782 3526 5795 3578
rect 5847 3526 5860 3578
rect 5912 3526 5925 3578
rect 5977 3526 5990 3578
rect 6042 3526 6055 3578
rect 6107 3526 6120 3578
rect 6172 3526 6185 3578
rect 6237 3526 6250 3578
rect 6302 3526 6315 3578
rect 6367 3526 6380 3578
rect 6432 3526 6445 3578
rect 6497 3526 6510 3578
rect 6562 3526 6575 3578
rect 6627 3526 6640 3578
rect 6692 3526 6705 3578
rect 6757 3526 6770 3578
rect 6822 3526 6835 3578
rect 6887 3526 6900 3578
rect 6952 3526 6965 3578
rect 7017 3526 7030 3578
rect 7082 3526 7095 3578
rect 7147 3526 7160 3578
rect 7212 3526 7225 3578
rect 7277 3526 7290 3578
rect 7342 3526 7355 3578
rect 7407 3526 7419 3578
rect 7471 3526 7483 3578
rect 7535 3526 7547 3578
rect 7599 3526 7611 3578
rect 7663 3526 7675 3578
rect 7727 3526 7739 3578
rect 7791 3526 7803 3578
rect 7855 3526 7867 3578
rect 7919 3526 7931 3578
rect 7983 3526 7995 3578
rect 8047 3526 8059 3578
rect 8111 3526 8123 3578
rect 8175 3526 8187 3578
rect 8239 3526 8251 3578
rect 8303 3526 8315 3578
rect 8367 3526 8379 3578
rect 8431 3526 8443 3578
rect 8495 3526 8507 3578
rect 8559 3526 8571 3578
rect 8623 3526 8635 3578
rect 8687 3526 8699 3578
rect 8751 3526 8763 3578
rect 8815 3526 8827 3578
rect 8879 3526 8891 3578
rect 8943 3526 8955 3578
rect 9007 3526 9019 3578
rect 9071 3526 9083 3578
rect 9135 3526 9147 3578
rect 9199 3526 9211 3578
rect 9263 3526 9275 3578
rect 9327 3526 9339 3578
rect 9391 3526 9403 3578
rect 9455 3526 9467 3578
rect 9519 3526 9531 3578
rect 9583 3526 9595 3578
rect 9647 3526 9659 3578
rect 9711 3526 9723 3578
rect 9775 3526 9787 3578
rect 9839 3526 9851 3578
rect 9903 3526 9915 3578
rect 9967 3526 9979 3578
rect 10031 3526 10043 3578
rect 10095 3526 10107 3578
rect 10159 3526 10171 3578
rect 10223 3526 10235 3578
rect 10287 3526 10299 3578
rect 10351 3526 10363 3578
rect 10415 3526 10427 3578
rect 10479 3526 10491 3578
rect 10543 3526 10555 3578
rect 10607 3526 10619 3578
rect 10671 3526 10683 3578
rect 10735 3526 10747 3578
rect 10799 3526 10811 3578
rect 10863 3526 10869 3578
tri 11151 3567 11250 3666 ne
rect 100 3416 4261 3526
tri 4261 3416 4371 3526 sw
rect 100 3410 11119 3416
rect 100 3358 3938 3410
rect 3990 3358 4020 3410
rect 4072 3358 4102 3410
rect 4154 3358 4184 3410
rect 4236 3358 4762 3410
rect 4814 3358 4844 3410
rect 4896 3358 4926 3410
rect 4978 3358 5008 3410
rect 5060 3358 5586 3410
rect 5638 3358 5668 3410
rect 5720 3358 5750 3410
rect 5802 3358 5832 3410
rect 5884 3358 6410 3410
rect 6462 3358 6492 3410
rect 6544 3358 6574 3410
rect 6626 3358 6656 3410
rect 6708 3358 7524 3410
rect 7576 3358 7606 3410
rect 7658 3358 7688 3410
rect 7740 3358 7770 3410
rect 7822 3358 8348 3410
rect 8400 3358 8430 3410
rect 8482 3358 8512 3410
rect 8564 3358 8594 3410
rect 8646 3358 9172 3410
rect 9224 3358 9254 3410
rect 9306 3358 9336 3410
rect 9388 3358 9418 3410
rect 9470 3358 9996 3410
rect 10048 3358 10078 3410
rect 10130 3358 10160 3410
rect 10212 3358 10242 3410
rect 10294 3358 10820 3410
rect 10872 3358 10902 3410
rect 10954 3358 10984 3410
rect 11036 3358 11066 3410
rect 11118 3358 11119 3410
rect 100 3344 11119 3358
rect 100 3292 3938 3344
rect 3990 3292 4020 3344
rect 4072 3292 4102 3344
rect 4154 3292 4184 3344
rect 4236 3292 4762 3344
rect 4814 3292 4844 3344
rect 4896 3292 4926 3344
rect 4978 3292 5008 3344
rect 5060 3292 5586 3344
rect 5638 3292 5668 3344
rect 5720 3292 5750 3344
rect 5802 3292 5832 3344
rect 5884 3292 6410 3344
rect 6462 3292 6492 3344
rect 6544 3292 6574 3344
rect 6626 3292 6656 3344
rect 6708 3292 7524 3344
rect 7576 3292 7606 3344
rect 7658 3292 7688 3344
rect 7740 3292 7770 3344
rect 7822 3292 8348 3344
rect 8400 3292 8430 3344
rect 8482 3292 8512 3344
rect 8564 3292 8594 3344
rect 8646 3292 9172 3344
rect 9224 3292 9254 3344
rect 9306 3292 9336 3344
rect 9388 3292 9418 3344
rect 9470 3292 9996 3344
rect 10048 3292 10078 3344
rect 10130 3292 10160 3344
rect 10212 3292 10242 3344
rect 10294 3292 10820 3344
rect 10872 3292 10902 3344
rect 10954 3292 10984 3344
rect 11036 3292 11066 3344
rect 11118 3292 11119 3344
rect 100 3278 11119 3292
rect 100 3226 3938 3278
rect 3990 3226 4020 3278
rect 4072 3226 4102 3278
rect 4154 3226 4184 3278
rect 4236 3226 4762 3278
rect 4814 3226 4844 3278
rect 4896 3226 4926 3278
rect 4978 3226 5008 3278
rect 5060 3226 5586 3278
rect 5638 3226 5668 3278
rect 5720 3226 5750 3278
rect 5802 3226 5832 3278
rect 5884 3226 6410 3278
rect 6462 3226 6492 3278
rect 6544 3226 6574 3278
rect 6626 3226 6656 3278
rect 6708 3226 7524 3278
rect 7576 3226 7606 3278
rect 7658 3226 7688 3278
rect 7740 3226 7770 3278
rect 7822 3226 8348 3278
rect 8400 3226 8430 3278
rect 8482 3226 8512 3278
rect 8564 3226 8594 3278
rect 8646 3226 9172 3278
rect 9224 3226 9254 3278
rect 9306 3226 9336 3278
rect 9388 3226 9418 3278
rect 9470 3226 9996 3278
rect 10048 3226 10078 3278
rect 10130 3226 10160 3278
rect 10212 3226 10242 3278
rect 10294 3226 10820 3278
rect 10872 3226 10902 3278
rect 10954 3226 10984 3278
rect 11036 3226 11066 3278
rect 11118 3226 11119 3278
rect 100 3212 11119 3226
rect 100 3160 3938 3212
rect 3990 3160 4020 3212
rect 4072 3160 4102 3212
rect 4154 3160 4184 3212
rect 4236 3160 4762 3212
rect 4814 3160 4844 3212
rect 4896 3160 4926 3212
rect 4978 3160 5008 3212
rect 5060 3160 5586 3212
rect 5638 3160 5668 3212
rect 5720 3160 5750 3212
rect 5802 3160 5832 3212
rect 5884 3160 6410 3212
rect 6462 3160 6492 3212
rect 6544 3160 6574 3212
rect 6626 3160 6656 3212
rect 6708 3160 7524 3212
rect 7576 3160 7606 3212
rect 7658 3160 7688 3212
rect 7740 3160 7770 3212
rect 7822 3160 8348 3212
rect 8400 3160 8430 3212
rect 8482 3160 8512 3212
rect 8564 3160 8594 3212
rect 8646 3160 9172 3212
rect 9224 3160 9254 3212
rect 9306 3160 9336 3212
rect 9388 3160 9418 3212
rect 9470 3160 9996 3212
rect 10048 3160 10078 3212
rect 10130 3160 10160 3212
rect 10212 3160 10242 3212
rect 10294 3160 10820 3212
rect 10872 3160 10902 3212
rect 10954 3160 10984 3212
rect 11036 3160 11066 3212
rect 11118 3160 11119 3212
rect 100 3146 11119 3160
rect 100 3094 3938 3146
rect 3990 3094 4020 3146
rect 4072 3094 4102 3146
rect 4154 3094 4184 3146
rect 4236 3094 4762 3146
rect 4814 3094 4844 3146
rect 4896 3094 4926 3146
rect 4978 3094 5008 3146
rect 5060 3094 5586 3146
rect 5638 3094 5668 3146
rect 5720 3094 5750 3146
rect 5802 3094 5832 3146
rect 5884 3094 6410 3146
rect 6462 3094 6492 3146
rect 6544 3094 6574 3146
rect 6626 3094 6656 3146
rect 6708 3094 7524 3146
rect 7576 3094 7606 3146
rect 7658 3094 7688 3146
rect 7740 3094 7770 3146
rect 7822 3094 8348 3146
rect 8400 3094 8430 3146
rect 8482 3094 8512 3146
rect 8564 3094 8594 3146
rect 8646 3094 9172 3146
rect 9224 3094 9254 3146
rect 9306 3094 9336 3146
rect 9388 3094 9418 3146
rect 9470 3094 9996 3146
rect 10048 3094 10078 3146
rect 10130 3094 10160 3146
rect 10212 3094 10242 3146
rect 10294 3094 10820 3146
rect 10872 3094 10902 3146
rect 10954 3094 10984 3146
rect 11036 3094 11066 3146
rect 11118 3094 11119 3146
rect 100 3079 11119 3094
rect 100 3042 3938 3079
rect 100 2862 1939 3042
rect 2119 2990 2132 3042
rect 2184 2990 2197 3042
rect 2249 2990 2262 3042
rect 2314 2990 2327 3042
rect 2379 2990 2392 3042
rect 2444 2990 2457 3042
rect 2509 2990 2522 3042
rect 2574 2990 2587 3042
rect 2639 2990 2652 3042
rect 2704 2990 2717 3042
rect 2769 2990 2782 3042
rect 2834 2990 2847 3042
rect 2899 2990 2912 3042
rect 2964 2990 2977 3042
rect 3029 2990 3042 3042
rect 3094 2990 3107 3042
rect 3159 3027 3938 3042
rect 3990 3027 4020 3079
rect 4072 3027 4102 3079
rect 4154 3027 4184 3079
rect 4236 3027 4762 3079
rect 4814 3027 4844 3079
rect 4896 3027 4926 3079
rect 4978 3027 5008 3079
rect 5060 3027 5586 3079
rect 5638 3027 5668 3079
rect 5720 3027 5750 3079
rect 5802 3027 5832 3079
rect 5884 3027 6410 3079
rect 6462 3027 6492 3079
rect 6544 3027 6574 3079
rect 6626 3027 6656 3079
rect 6708 3027 7524 3079
rect 7576 3027 7606 3079
rect 7658 3027 7688 3079
rect 7740 3027 7770 3079
rect 7822 3027 8348 3079
rect 8400 3027 8430 3079
rect 8482 3027 8512 3079
rect 8564 3027 8594 3079
rect 8646 3027 9172 3079
rect 9224 3027 9254 3079
rect 9306 3027 9336 3079
rect 9388 3027 9418 3079
rect 9470 3027 9996 3079
rect 10048 3027 10078 3079
rect 10130 3027 10160 3079
rect 10212 3027 10242 3079
rect 10294 3027 10820 3079
rect 10872 3027 10902 3079
rect 10954 3027 10984 3079
rect 11036 3027 11066 3079
rect 11118 3027 11119 3079
rect 3159 3012 11119 3027
rect 3159 2990 3938 3012
rect 2119 2978 3938 2990
rect 2119 2926 2132 2978
rect 2184 2926 2197 2978
rect 2249 2926 2262 2978
rect 2314 2926 2327 2978
rect 2379 2926 2392 2978
rect 2444 2926 2457 2978
rect 2509 2926 2522 2978
rect 2574 2926 2587 2978
rect 2639 2926 2652 2978
rect 2704 2926 2717 2978
rect 2769 2926 2782 2978
rect 2834 2926 2847 2978
rect 2899 2926 2912 2978
rect 2964 2926 2977 2978
rect 3029 2926 3042 2978
rect 3094 2926 3107 2978
rect 2055 2914 3107 2926
rect 3223 2960 3938 2978
rect 3990 2960 4020 3012
rect 4072 2960 4102 3012
rect 4154 2960 4184 3012
rect 4236 2960 4762 3012
rect 4814 2960 4844 3012
rect 4896 2960 4926 3012
rect 4978 2960 5008 3012
rect 5060 2960 5586 3012
rect 5638 2960 5668 3012
rect 5720 2960 5750 3012
rect 5802 2960 5832 3012
rect 5884 2960 6410 3012
rect 6462 2960 6492 3012
rect 6544 2960 6574 3012
rect 6626 2960 6656 3012
rect 6708 2960 7524 3012
rect 7576 2960 7606 3012
rect 7658 2960 7688 3012
rect 7740 2960 7770 3012
rect 7822 2960 8348 3012
rect 8400 2960 8430 3012
rect 8482 2960 8512 3012
rect 8564 2960 8594 3012
rect 8646 2960 9172 3012
rect 9224 2960 9254 3012
rect 9306 2960 9336 3012
rect 9388 2960 9418 3012
rect 9470 2960 9996 3012
rect 10048 2960 10078 3012
rect 10130 2960 10160 3012
rect 10212 2960 10242 3012
rect 10294 2960 10820 3012
rect 10872 2960 10902 3012
rect 10954 2960 10984 3012
rect 11036 2960 11066 3012
rect 11118 2960 11119 3012
rect 3223 2945 11119 2960
rect 2055 2862 2068 2914
rect 2120 2862 2133 2914
rect 2185 2862 2198 2914
rect 2250 2862 2263 2914
rect 2315 2862 2328 2914
rect 2380 2862 2393 2914
rect 2445 2862 2458 2914
rect 2510 2862 2523 2914
rect 2575 2862 2588 2914
rect 2640 2862 2653 2914
rect 2705 2862 2718 2914
rect 2770 2862 2783 2914
rect 2835 2862 2848 2914
rect 2900 2862 2913 2914
rect 2965 2862 2978 2914
rect 3030 2862 3043 2914
rect 100 2850 3043 2862
rect 3223 2893 3938 2945
rect 3990 2893 4020 2945
rect 4072 2893 4102 2945
rect 4154 2893 4184 2945
rect 4236 2893 4762 2945
rect 4814 2893 4844 2945
rect 4896 2893 4926 2945
rect 4978 2893 5008 2945
rect 5060 2893 5586 2945
rect 5638 2893 5668 2945
rect 5720 2893 5750 2945
rect 5802 2893 5832 2945
rect 5884 2893 6410 2945
rect 6462 2893 6492 2945
rect 6544 2893 6574 2945
rect 6626 2893 6656 2945
rect 6708 2893 7524 2945
rect 7576 2893 7606 2945
rect 7658 2893 7688 2945
rect 7740 2893 7770 2945
rect 7822 2893 8348 2945
rect 8400 2893 8430 2945
rect 8482 2893 8512 2945
rect 8564 2893 8594 2945
rect 8646 2893 9172 2945
rect 9224 2893 9254 2945
rect 9306 2893 9336 2945
rect 9388 2893 9418 2945
rect 9470 2893 9996 2945
rect 10048 2893 10078 2945
rect 10130 2893 10160 2945
rect 10212 2893 10242 2945
rect 10294 2893 10820 2945
rect 10872 2893 10902 2945
rect 10954 2893 10984 2945
rect 11036 2893 11066 2945
rect 11118 2893 11119 2945
rect 3223 2878 11119 2893
rect 100 2798 1939 2850
rect 1991 2798 2004 2850
rect 2056 2798 2069 2850
rect 2121 2798 2134 2850
rect 2186 2798 2199 2850
rect 2251 2798 2264 2850
rect 2316 2798 2329 2850
rect 2381 2798 2394 2850
rect 2446 2798 2459 2850
rect 2511 2798 2524 2850
rect 2576 2798 2589 2850
rect 2641 2798 2654 2850
rect 2706 2798 2719 2850
rect 2771 2798 2784 2850
rect 2836 2798 2849 2850
rect 2901 2798 2914 2850
rect 2966 2798 2979 2850
rect 100 2786 2979 2798
rect 3223 2826 3938 2878
rect 3990 2826 4020 2878
rect 4072 2826 4102 2878
rect 4154 2826 4184 2878
rect 4236 2826 4762 2878
rect 4814 2826 4844 2878
rect 4896 2826 4926 2878
rect 4978 2826 5008 2878
rect 5060 2826 5586 2878
rect 5638 2826 5668 2878
rect 5720 2826 5750 2878
rect 5802 2826 5832 2878
rect 5884 2826 6410 2878
rect 6462 2826 6492 2878
rect 6544 2826 6574 2878
rect 6626 2826 6656 2878
rect 6708 2826 7524 2878
rect 7576 2826 7606 2878
rect 7658 2826 7688 2878
rect 7740 2826 7770 2878
rect 7822 2826 8348 2878
rect 8400 2826 8430 2878
rect 8482 2826 8512 2878
rect 8564 2826 8594 2878
rect 8646 2826 9172 2878
rect 9224 2826 9254 2878
rect 9306 2826 9336 2878
rect 9388 2826 9418 2878
rect 9470 2826 9996 2878
rect 10048 2826 10078 2878
rect 10130 2826 10160 2878
rect 10212 2826 10242 2878
rect 10294 2826 10820 2878
rect 10872 2826 10902 2878
rect 10954 2826 10984 2878
rect 11036 2826 11066 2878
rect 11118 2826 11119 2878
rect 3223 2811 11119 2826
rect 100 2734 1939 2786
rect 1991 2734 2004 2786
rect 2056 2734 2069 2786
rect 2121 2734 2134 2786
rect 2186 2734 2199 2786
rect 2251 2734 2264 2786
rect 2316 2734 2329 2786
rect 2381 2734 2394 2786
rect 2446 2734 2459 2786
rect 2511 2734 2524 2786
rect 2576 2734 2589 2786
rect 2641 2734 2654 2786
rect 2706 2734 2719 2786
rect 2771 2734 2784 2786
rect 2836 2734 2849 2786
rect 2901 2734 2915 2786
rect 100 2722 2915 2734
rect 3223 2759 3938 2811
rect 3990 2759 4020 2811
rect 4072 2759 4102 2811
rect 4154 2759 4184 2811
rect 4236 2759 4762 2811
rect 4814 2759 4844 2811
rect 4896 2759 4926 2811
rect 4978 2759 5008 2811
rect 5060 2759 5586 2811
rect 5638 2759 5668 2811
rect 5720 2759 5750 2811
rect 5802 2759 5832 2811
rect 5884 2759 6410 2811
rect 6462 2759 6492 2811
rect 6544 2759 6574 2811
rect 6626 2759 6656 2811
rect 6708 2759 7524 2811
rect 7576 2759 7606 2811
rect 7658 2759 7688 2811
rect 7740 2759 7770 2811
rect 7822 2759 8348 2811
rect 8400 2759 8430 2811
rect 8482 2759 8512 2811
rect 8564 2759 8594 2811
rect 8646 2759 9172 2811
rect 9224 2759 9254 2811
rect 9306 2759 9336 2811
rect 9388 2759 9418 2811
rect 9470 2759 9996 2811
rect 10048 2759 10078 2811
rect 10130 2759 10160 2811
rect 10212 2759 10242 2811
rect 10294 2759 10820 2811
rect 10872 2759 10902 2811
rect 10954 2759 10984 2811
rect 11036 2759 11066 2811
rect 11118 2759 11119 2811
rect 3223 2744 11119 2759
rect 100 2670 1939 2722
rect 1991 2670 2004 2722
rect 2056 2670 2069 2722
rect 2121 2670 2134 2722
rect 2186 2670 2199 2722
rect 2251 2670 2264 2722
rect 2316 2670 2329 2722
rect 2381 2670 2394 2722
rect 2446 2670 2459 2722
rect 2511 2670 2524 2722
rect 2576 2670 2589 2722
rect 2641 2670 2654 2722
rect 2706 2670 2719 2722
rect 2771 2670 2785 2722
rect 2837 2670 2851 2722
rect 100 2658 2851 2670
rect 3223 2692 3938 2744
rect 3990 2692 4020 2744
rect 4072 2692 4102 2744
rect 4154 2692 4184 2744
rect 4236 2692 4762 2744
rect 4814 2692 4844 2744
rect 4896 2692 4926 2744
rect 4978 2692 5008 2744
rect 5060 2692 5586 2744
rect 5638 2692 5668 2744
rect 5720 2692 5750 2744
rect 5802 2692 5832 2744
rect 5884 2692 6410 2744
rect 6462 2692 6492 2744
rect 6544 2692 6574 2744
rect 6626 2692 6656 2744
rect 6708 2692 7524 2744
rect 7576 2692 7606 2744
rect 7658 2692 7688 2744
rect 7740 2692 7770 2744
rect 7822 2692 8348 2744
rect 8400 2692 8430 2744
rect 8482 2692 8512 2744
rect 8564 2692 8594 2744
rect 8646 2692 9172 2744
rect 9224 2692 9254 2744
rect 9306 2692 9336 2744
rect 9388 2692 9418 2744
rect 9470 2692 9996 2744
rect 10048 2692 10078 2744
rect 10130 2692 10160 2744
rect 10212 2692 10242 2744
rect 10294 2692 10820 2744
rect 10872 2692 10902 2744
rect 10954 2692 10984 2744
rect 11036 2692 11066 2744
rect 11118 2692 11119 2744
rect 3223 2677 11119 2692
rect 100 2606 1939 2658
rect 1991 2606 2004 2658
rect 2056 2606 2069 2658
rect 2121 2606 2134 2658
rect 2186 2606 2199 2658
rect 2251 2606 2264 2658
rect 2316 2606 2329 2658
rect 2381 2606 2394 2658
rect 2446 2606 2459 2658
rect 2511 2606 2524 2658
rect 2576 2606 2589 2658
rect 2641 2606 2655 2658
rect 2707 2606 2721 2658
rect 2773 2606 2787 2658
rect 100 2594 2787 2606
rect 3223 2625 3938 2677
rect 3990 2625 4020 2677
rect 4072 2625 4102 2677
rect 4154 2625 4184 2677
rect 4236 2625 4762 2677
rect 4814 2625 4844 2677
rect 4896 2625 4926 2677
rect 4978 2625 5008 2677
rect 5060 2625 5586 2677
rect 5638 2625 5668 2677
rect 5720 2625 5750 2677
rect 5802 2625 5832 2677
rect 5884 2625 6410 2677
rect 6462 2625 6492 2677
rect 6544 2625 6574 2677
rect 6626 2625 6656 2677
rect 6708 2625 7524 2677
rect 7576 2625 7606 2677
rect 7658 2625 7688 2677
rect 7740 2625 7770 2677
rect 7822 2625 8348 2677
rect 8400 2625 8430 2677
rect 8482 2625 8512 2677
rect 8564 2625 8594 2677
rect 8646 2625 9172 2677
rect 9224 2625 9254 2677
rect 9306 2625 9336 2677
rect 9388 2625 9418 2677
rect 9470 2625 9996 2677
rect 10048 2625 10078 2677
rect 10130 2625 10160 2677
rect 10212 2625 10242 2677
rect 10294 2625 10820 2677
rect 10872 2625 10902 2677
rect 10954 2625 10984 2677
rect 11036 2625 11066 2677
rect 11118 2625 11119 2677
rect 3223 2610 11119 2625
rect 100 2542 1939 2594
rect 1991 2542 2004 2594
rect 2056 2542 2069 2594
rect 2121 2542 2134 2594
rect 2186 2542 2199 2594
rect 2251 2542 2264 2594
rect 2316 2542 2329 2594
rect 2381 2542 2394 2594
rect 2446 2542 2459 2594
rect 2511 2542 2525 2594
rect 2577 2542 2591 2594
rect 2643 2542 2657 2594
rect 2709 2542 2723 2594
rect 100 2530 2723 2542
rect 3223 2558 3938 2610
rect 3990 2558 4020 2610
rect 4072 2558 4102 2610
rect 4154 2558 4184 2610
rect 4236 2558 4762 2610
rect 4814 2558 4844 2610
rect 4896 2558 4926 2610
rect 4978 2558 5008 2610
rect 5060 2558 5586 2610
rect 5638 2558 5668 2610
rect 5720 2558 5750 2610
rect 5802 2558 5832 2610
rect 5884 2558 6410 2610
rect 6462 2558 6492 2610
rect 6544 2558 6574 2610
rect 6626 2558 6656 2610
rect 6708 2558 7524 2610
rect 7576 2558 7606 2610
rect 7658 2558 7688 2610
rect 7740 2558 7770 2610
rect 7822 2558 8348 2610
rect 8400 2558 8430 2610
rect 8482 2558 8512 2610
rect 8564 2558 8594 2610
rect 8646 2558 9172 2610
rect 9224 2558 9254 2610
rect 9306 2558 9336 2610
rect 9388 2558 9418 2610
rect 9470 2558 9996 2610
rect 10048 2558 10078 2610
rect 10130 2558 10160 2610
rect 10212 2558 10242 2610
rect 10294 2558 10820 2610
rect 10872 2558 10902 2610
rect 10954 2558 10984 2610
rect 11036 2558 11066 2610
rect 11118 2558 11119 2610
rect 3223 2543 11119 2558
rect 100 2478 1939 2530
rect 1991 2478 2004 2530
rect 2056 2478 2069 2530
rect 2121 2478 2134 2530
rect 2186 2478 2199 2530
rect 2251 2478 2264 2530
rect 2316 2478 2329 2530
rect 2381 2478 2395 2530
rect 2447 2478 2461 2530
rect 2513 2478 2527 2530
rect 2579 2478 2593 2530
rect 2645 2478 2659 2530
rect 100 2466 2659 2478
rect 100 2414 1939 2466
rect 1991 2414 2004 2466
rect 2056 2414 2069 2466
rect 2121 2414 2134 2466
rect 2186 2414 2199 2466
rect 2251 2414 2265 2466
rect 2317 2414 2331 2466
rect 2383 2414 2397 2466
rect 2449 2414 2463 2466
rect 2515 2414 2529 2466
rect 2581 2414 2595 2466
rect 2647 2414 2659 2466
rect 100 2402 2659 2414
rect 100 2350 1939 2402
rect 1991 2350 2004 2402
rect 2056 2350 2069 2402
rect 2121 2350 2135 2402
rect 2187 2350 2201 2402
rect 2253 2350 2267 2402
rect 2319 2350 2333 2402
rect 2385 2350 2399 2402
rect 2451 2350 2465 2402
rect 2517 2350 2531 2402
rect 2583 2401 2659 2402
rect 2583 2350 2595 2401
rect 100 2349 2595 2350
rect 2647 2350 2659 2401
rect 3223 2491 3938 2543
rect 3990 2491 4020 2543
rect 4072 2491 4102 2543
rect 4154 2491 4184 2543
rect 4236 2491 4762 2543
rect 4814 2491 4844 2543
rect 4896 2491 4926 2543
rect 4978 2491 5008 2543
rect 5060 2491 5586 2543
rect 5638 2491 5668 2543
rect 5720 2491 5750 2543
rect 5802 2491 5832 2543
rect 5884 2491 6410 2543
rect 6462 2491 6492 2543
rect 6544 2491 6574 2543
rect 6626 2491 6656 2543
rect 6708 2491 7524 2543
rect 7576 2491 7606 2543
rect 7658 2491 7688 2543
rect 7740 2491 7770 2543
rect 7822 2491 8348 2543
rect 8400 2491 8430 2543
rect 8482 2491 8512 2543
rect 8564 2491 8594 2543
rect 8646 2491 9172 2543
rect 9224 2491 9254 2543
rect 9306 2491 9336 2543
rect 9388 2491 9418 2543
rect 9470 2491 9996 2543
rect 10048 2491 10078 2543
rect 10130 2491 10160 2543
rect 10212 2491 10242 2543
rect 10294 2491 10820 2543
rect 10872 2491 10902 2543
rect 10954 2491 10984 2543
rect 11036 2491 11066 2543
rect 11118 2491 11119 2543
rect 3223 2476 11119 2491
rect 3223 2424 3938 2476
rect 3990 2424 4020 2476
rect 4072 2424 4102 2476
rect 4154 2424 4184 2476
rect 4236 2424 4762 2476
rect 4814 2424 4844 2476
rect 4896 2424 4926 2476
rect 4978 2424 5008 2476
rect 5060 2424 5586 2476
rect 5638 2424 5668 2476
rect 5720 2424 5750 2476
rect 5802 2424 5832 2476
rect 5884 2424 6410 2476
rect 6462 2424 6492 2476
rect 6544 2424 6574 2476
rect 6626 2424 6656 2476
rect 6708 2424 7524 2476
rect 7576 2424 7606 2476
rect 7658 2424 7688 2476
rect 7740 2424 7770 2476
rect 7822 2424 8348 2476
rect 8400 2424 8430 2476
rect 8482 2424 8512 2476
rect 8564 2424 8594 2476
rect 8646 2424 9172 2476
rect 9224 2424 9254 2476
rect 9306 2424 9336 2476
rect 9388 2424 9418 2476
rect 9470 2424 9996 2476
rect 10048 2424 10078 2476
rect 10130 2424 10160 2476
rect 10212 2424 10242 2476
rect 10294 2424 10820 2476
rect 10872 2424 10902 2476
rect 10954 2424 10984 2476
rect 11036 2424 11066 2476
rect 11118 2424 11119 2476
rect 3223 2409 11119 2424
rect 3223 2357 3938 2409
rect 3990 2357 4020 2409
rect 4072 2357 4102 2409
rect 4154 2357 4184 2409
rect 4236 2357 4762 2409
rect 4814 2357 4844 2409
rect 4896 2357 4926 2409
rect 4978 2357 5008 2409
rect 5060 2357 5586 2409
rect 5638 2357 5668 2409
rect 5720 2357 5750 2409
rect 5802 2357 5832 2409
rect 5884 2357 6410 2409
rect 6462 2357 6492 2409
rect 6544 2357 6574 2409
rect 6626 2357 6656 2409
rect 6708 2357 7524 2409
rect 7576 2357 7606 2409
rect 7658 2357 7688 2409
rect 7740 2357 7770 2409
rect 7822 2357 8348 2409
rect 8400 2357 8430 2409
rect 8482 2357 8512 2409
rect 8564 2357 8594 2409
rect 8646 2357 9172 2409
rect 9224 2357 9254 2409
rect 9306 2357 9336 2409
rect 9388 2357 9418 2409
rect 9470 2357 9996 2409
rect 10048 2357 10078 2409
rect 10130 2357 10160 2409
rect 10212 2357 10242 2409
rect 10294 2357 10820 2409
rect 10872 2357 10902 2409
rect 10954 2357 10984 2409
rect 11036 2357 11066 2409
rect 11118 2357 11119 2409
rect 2647 2349 2723 2350
rect 100 2338 2723 2349
rect 100 2286 1939 2338
rect 1991 2286 2005 2338
rect 2057 2286 2071 2338
rect 2123 2286 2137 2338
rect 2189 2286 2203 2338
rect 2255 2286 2269 2338
rect 2321 2286 2335 2338
rect 2387 2286 2401 2338
rect 2453 2286 2467 2338
rect 2519 2337 2723 2338
rect 2519 2286 2531 2337
rect 100 2285 2531 2286
rect 2583 2336 2659 2337
rect 2583 2285 2595 2336
rect 100 2284 2595 2285
rect 2647 2285 2659 2336
rect 2711 2286 2723 2337
rect 3223 2342 11119 2357
rect 3223 2290 3938 2342
rect 3990 2290 4020 2342
rect 4072 2290 4102 2342
rect 4154 2290 4184 2342
rect 4236 2290 4762 2342
rect 4814 2290 4844 2342
rect 4896 2290 4926 2342
rect 4978 2290 5008 2342
rect 5060 2290 5586 2342
rect 5638 2290 5668 2342
rect 5720 2290 5750 2342
rect 5802 2290 5832 2342
rect 5884 2290 6410 2342
rect 6462 2290 6492 2342
rect 6544 2290 6574 2342
rect 6626 2290 6656 2342
rect 6708 2290 7524 2342
rect 7576 2290 7606 2342
rect 7658 2290 7688 2342
rect 7740 2290 7770 2342
rect 7822 2290 8348 2342
rect 8400 2290 8430 2342
rect 8482 2290 8512 2342
rect 8564 2290 8594 2342
rect 8646 2290 9172 2342
rect 9224 2290 9254 2342
rect 9306 2290 9336 2342
rect 9388 2290 9418 2342
rect 9470 2290 9996 2342
rect 10048 2290 10078 2342
rect 10130 2290 10160 2342
rect 10212 2290 10242 2342
rect 10294 2290 10820 2342
rect 10872 2290 10902 2342
rect 10954 2290 10984 2342
rect 11036 2290 11066 2342
rect 11118 2290 11119 2342
rect 2711 2285 2787 2286
rect 2647 2284 2787 2285
rect 100 2274 2787 2284
rect 100 2222 1939 2274
rect 1991 2222 2005 2274
rect 2057 2222 2071 2274
rect 2123 2222 2137 2274
rect 2189 2222 2203 2274
rect 2255 2222 2269 2274
rect 2321 2222 2336 2274
rect 2388 2222 2403 2274
rect 2455 2273 2787 2274
rect 2455 2222 2467 2273
rect 100 2221 2467 2222
rect 2519 2272 2723 2273
rect 2519 2221 2531 2272
rect 100 2220 2531 2221
rect 2583 2271 2659 2272
rect 2583 2220 2595 2271
rect 100 2219 2595 2220
rect 2647 2220 2659 2271
rect 2711 2221 2723 2272
rect 2775 2222 2787 2273
rect 3223 2275 11119 2290
rect 3223 2223 3938 2275
rect 3990 2223 4020 2275
rect 4072 2223 4102 2275
rect 4154 2223 4184 2275
rect 4236 2223 4762 2275
rect 4814 2223 4844 2275
rect 4896 2223 4926 2275
rect 4978 2223 5008 2275
rect 5060 2223 5586 2275
rect 5638 2223 5668 2275
rect 5720 2223 5750 2275
rect 5802 2223 5832 2275
rect 5884 2223 6410 2275
rect 6462 2223 6492 2275
rect 6544 2223 6574 2275
rect 6626 2223 6656 2275
rect 6708 2223 7524 2275
rect 7576 2223 7606 2275
rect 7658 2223 7688 2275
rect 7740 2223 7770 2275
rect 7822 2223 8348 2275
rect 8400 2223 8430 2275
rect 8482 2223 8512 2275
rect 8564 2223 8594 2275
rect 8646 2223 9172 2275
rect 9224 2223 9254 2275
rect 9306 2223 9336 2275
rect 9388 2223 9418 2275
rect 9470 2223 9996 2275
rect 10048 2223 10078 2275
rect 10130 2223 10160 2275
rect 10212 2223 10242 2275
rect 10294 2223 10820 2275
rect 10872 2223 10902 2275
rect 10954 2223 10984 2275
rect 11036 2223 11066 2275
rect 11118 2223 11119 2275
rect 2775 2221 2851 2222
rect 2711 2220 2851 2221
rect 2647 2219 2851 2220
rect 100 2209 2851 2219
rect 100 2157 2403 2209
rect 2455 2208 2787 2209
rect 2455 2157 2467 2208
rect 100 2156 2467 2157
rect 2519 2207 2723 2208
rect 2519 2156 2531 2207
rect 100 2155 2531 2156
rect 2583 2206 2659 2207
rect 2583 2155 2595 2206
rect 100 2154 2595 2155
rect 2647 2155 2659 2206
rect 2711 2156 2723 2207
rect 2775 2157 2787 2208
rect 2839 2158 2851 2209
rect 3223 2208 11119 2223
rect 2839 2157 2915 2158
rect 2775 2156 2915 2157
rect 2711 2155 2915 2156
rect 2647 2154 2915 2155
rect 100 2145 2915 2154
rect 100 2144 2851 2145
rect 100 2092 2403 2144
rect 2455 2143 2787 2144
rect 2455 2092 2467 2143
rect 100 2091 2467 2092
rect 2519 2142 2723 2143
rect 2519 2091 2531 2142
rect 100 2090 2531 2091
rect 2583 2141 2659 2142
rect 2583 2090 2595 2141
rect 100 2089 2595 2090
rect 2647 2090 2659 2141
rect 2711 2091 2723 2142
rect 2775 2092 2787 2143
rect 2839 2093 2851 2144
rect 2903 2094 2915 2145
rect 3223 2156 3938 2208
rect 3990 2156 4020 2208
rect 4072 2156 4102 2208
rect 4154 2156 4184 2208
rect 4236 2156 4762 2208
rect 4814 2156 4844 2208
rect 4896 2156 4926 2208
rect 4978 2156 5008 2208
rect 5060 2156 5586 2208
rect 5638 2156 5668 2208
rect 5720 2156 5750 2208
rect 5802 2156 5832 2208
rect 5884 2156 6410 2208
rect 6462 2156 6492 2208
rect 6544 2156 6574 2208
rect 6626 2156 6656 2208
rect 6708 2156 7524 2208
rect 7576 2156 7606 2208
rect 7658 2156 7688 2208
rect 7740 2156 7770 2208
rect 7822 2156 8348 2208
rect 8400 2156 8430 2208
rect 8482 2156 8512 2208
rect 8564 2156 8594 2208
rect 8646 2156 9172 2208
rect 9224 2156 9254 2208
rect 9306 2156 9336 2208
rect 9388 2156 9418 2208
rect 9470 2156 9996 2208
rect 10048 2156 10078 2208
rect 10130 2156 10160 2208
rect 10212 2156 10242 2208
rect 10294 2156 10820 2208
rect 10872 2156 10902 2208
rect 10954 2156 10984 2208
rect 11036 2156 11066 2208
rect 11118 2156 11119 2208
rect 3223 2141 11119 2156
rect 2903 2093 2979 2094
rect 2839 2092 2979 2093
rect 2775 2091 2979 2092
rect 2711 2090 2979 2091
rect 2647 2089 2979 2090
rect 100 2081 2979 2089
rect 100 2080 2915 2081
rect 100 2079 2851 2080
rect 100 2043 2403 2079
rect 100 2027 2147 2043
tri 2147 2027 2163 2043 nw
tri 2326 2027 2342 2043 ne
rect 2342 2027 2403 2043
rect 2455 2078 2787 2079
rect 2455 2027 2467 2078
rect 100 2026 2146 2027
tri 2146 2026 2147 2027 nw
tri 2342 2026 2343 2027 ne
rect 2343 2026 2467 2027
rect 2519 2077 2723 2078
rect 2519 2026 2531 2077
rect 100 2025 2145 2026
tri 2145 2025 2146 2026 nw
tri 2343 2025 2344 2026 ne
rect 2344 2025 2531 2026
rect 2583 2076 2659 2077
rect 2583 2025 2595 2076
rect 100 2024 2144 2025
tri 2144 2024 2145 2025 nw
tri 2344 2024 2345 2025 ne
rect 2345 2024 2595 2025
rect 2647 2025 2659 2076
rect 2711 2026 2723 2077
rect 2775 2027 2787 2078
rect 2839 2028 2851 2079
rect 2903 2029 2915 2080
rect 2967 2030 2979 2081
rect 3223 2089 3938 2141
rect 3990 2089 4020 2141
rect 4072 2089 4102 2141
rect 4154 2089 4184 2141
rect 4236 2089 4762 2141
rect 4814 2089 4844 2141
rect 4896 2089 4926 2141
rect 4978 2089 5008 2141
rect 5060 2089 5586 2141
rect 5638 2089 5668 2141
rect 5720 2089 5750 2141
rect 5802 2089 5832 2141
rect 5884 2089 6410 2141
rect 6462 2089 6492 2141
rect 6544 2089 6574 2141
rect 6626 2089 6656 2141
rect 6708 2089 7524 2141
rect 7576 2089 7606 2141
rect 7658 2089 7688 2141
rect 7740 2089 7770 2141
rect 7822 2089 8348 2141
rect 8400 2089 8430 2141
rect 8482 2089 8512 2141
rect 8564 2089 8594 2141
rect 8646 2089 9172 2141
rect 9224 2089 9254 2141
rect 9306 2089 9336 2141
rect 9388 2089 9418 2141
rect 9470 2089 9996 2141
rect 10048 2089 10078 2141
rect 10130 2089 10160 2141
rect 10212 2089 10242 2141
rect 10294 2089 10820 2141
rect 10872 2089 10902 2141
rect 10954 2089 10984 2141
rect 11036 2089 11066 2141
rect 11118 2089 11119 2141
rect 3223 2074 11119 2089
rect 2967 2029 3043 2030
rect 2903 2028 3043 2029
rect 2839 2027 3043 2028
rect 2775 2026 3043 2027
rect 2711 2025 3043 2026
rect 2647 2024 3043 2025
rect 100 2017 2137 2024
tri 2137 2017 2144 2024 nw
tri 2345 2017 2352 2024 ne
rect 2352 2017 3043 2024
rect 100 2016 2136 2017
tri 2136 2016 2137 2017 nw
tri 2352 2016 2353 2017 ne
rect 2353 2016 2979 2017
rect 100 2015 2135 2016
tri 2135 2015 2136 2016 nw
tri 2353 2015 2354 2016 ne
rect 2354 2015 2915 2016
rect 100 2014 2134 2015
tri 2134 2014 2135 2015 nw
tri 2354 2014 2355 2015 ne
rect 2355 2014 2851 2015
rect 100 1994 2114 2014
tri 2114 1994 2134 2014 nw
tri 2355 1994 2375 2014 ne
rect 2375 1994 2403 2014
rect 100 1609 2084 1994
tri 2084 1964 2114 1994 nw
tri 2375 1966 2403 1994 ne
rect 2455 2013 2787 2014
rect 2455 1962 2467 2013
rect 2403 1961 2467 1962
rect 2519 2012 2723 2013
rect 2519 1961 2531 2012
rect 2403 1960 2531 1961
rect 2583 2011 2659 2012
rect 2583 1960 2595 2011
rect 2403 1959 2595 1960
rect 2647 1960 2659 2011
rect 2711 1961 2723 2012
rect 2775 1962 2787 2013
rect 2839 1963 2851 2014
rect 2903 1964 2915 2015
rect 2967 1965 2979 2016
rect 3031 1966 3043 2017
rect 3223 2022 3938 2074
rect 3990 2022 4020 2074
rect 4072 2022 4102 2074
rect 4154 2022 4184 2074
rect 4236 2022 4762 2074
rect 4814 2022 4844 2074
rect 4896 2022 4926 2074
rect 4978 2022 5008 2074
rect 5060 2022 5586 2074
rect 5638 2022 5668 2074
rect 5720 2022 5750 2074
rect 5802 2022 5832 2074
rect 5884 2022 6410 2074
rect 6462 2022 6492 2074
rect 6544 2022 6574 2074
rect 6626 2022 6656 2074
rect 6708 2022 7524 2074
rect 7576 2022 7606 2074
rect 7658 2022 7688 2074
rect 7740 2022 7770 2074
rect 7822 2022 8348 2074
rect 8400 2022 8430 2074
rect 8482 2022 8512 2074
rect 8564 2022 8594 2074
rect 8646 2022 9172 2074
rect 9224 2022 9254 2074
rect 9306 2022 9336 2074
rect 9388 2022 9418 2074
rect 9470 2022 9996 2074
rect 10048 2022 10078 2074
rect 10130 2022 10160 2074
rect 10212 2022 10242 2074
rect 10294 2022 10820 2074
rect 10872 2022 10902 2074
rect 10954 2022 10984 2074
rect 11036 2022 11066 2074
rect 11118 2022 11119 2074
rect 3223 2016 11119 2022
rect 3223 1994 3493 2016
tri 3493 1994 3515 2016 nw
rect 3223 1966 3465 1994
tri 3465 1966 3493 1994 nw
tri 11222 1966 11250 1994 se
rect 11250 1966 14940 3666
rect 3031 1965 3107 1966
rect 2967 1964 3107 1965
rect 2903 1963 3107 1964
rect 2839 1962 3107 1963
rect 2775 1961 3107 1962
rect 2711 1960 3107 1961
rect 2647 1959 3107 1960
rect 2403 1953 3107 1959
rect 2403 1952 3043 1953
rect 2403 1951 2979 1952
rect 2403 1950 2915 1951
rect 2403 1949 2851 1950
rect 2455 1948 2787 1949
rect 2455 1897 2467 1948
rect 2403 1896 2467 1897
rect 2519 1947 2723 1948
rect 2519 1896 2531 1947
rect 2403 1895 2531 1896
rect 2583 1946 2659 1947
rect 2583 1895 2595 1946
rect 2403 1894 2595 1895
rect 2647 1895 2659 1946
rect 2711 1896 2723 1947
rect 2775 1897 2787 1948
rect 2839 1898 2851 1949
rect 2903 1899 2915 1950
rect 2967 1900 2979 1951
rect 3031 1901 3043 1952
rect 3095 1902 3107 1953
rect 3223 1964 3463 1966
tri 3463 1964 3465 1966 nw
tri 11220 1964 11222 1966 se
rect 11222 1964 14940 1966
rect 3223 1908 3407 1964
tri 3407 1908 3463 1964 nw
tri 11164 1908 11220 1964 se
rect 11220 1908 14940 1964
rect 3223 1902 3401 1908
tri 3401 1902 3407 1908 nw
rect 3526 1902 10707 1908
rect 3095 1901 3372 1902
rect 3031 1900 3372 1901
rect 2967 1899 3372 1900
rect 2903 1898 3372 1899
rect 2839 1897 3372 1898
rect 2775 1896 3372 1897
rect 2711 1895 3372 1896
rect 2647 1894 3372 1895
rect 2403 1889 3372 1894
rect 2403 1888 3107 1889
rect 2403 1887 3043 1888
rect 2403 1886 2979 1887
rect 2403 1885 2915 1886
rect 2403 1884 2851 1885
rect 2455 1883 2787 1884
rect 2455 1832 2467 1883
rect 2403 1831 2467 1832
rect 2519 1882 2723 1883
rect 2519 1831 2531 1882
rect 2403 1830 2531 1831
rect 2583 1881 2659 1882
rect 2583 1830 2595 1881
rect 2403 1829 2595 1830
rect 2647 1830 2659 1881
rect 2711 1831 2723 1882
rect 2775 1832 2787 1883
rect 2839 1833 2851 1884
rect 2903 1834 2915 1885
rect 2967 1835 2979 1886
rect 3031 1836 3043 1887
rect 3095 1837 3107 1888
rect 3159 1837 3171 1889
rect 3223 1837 3372 1889
tri 3372 1873 3401 1902 nw
rect 3095 1836 3372 1837
rect 3031 1835 3372 1836
rect 2967 1834 3372 1835
rect 2903 1833 3372 1834
rect 2839 1832 3372 1833
rect 2775 1831 3372 1832
rect 2711 1830 3372 1831
rect 2647 1829 3372 1830
rect 2403 1824 3372 1829
rect 2403 1823 3107 1824
rect 2403 1822 3043 1823
rect 2403 1821 2979 1822
rect 2403 1820 2915 1821
rect 2403 1819 2851 1820
rect 2403 1818 2787 1819
rect 2455 1766 2467 1818
rect 2519 1817 2723 1818
rect 2519 1766 2531 1817
rect 2403 1765 2531 1766
rect 2583 1816 2659 1817
rect 2583 1765 2595 1816
rect 2403 1764 2595 1765
rect 2647 1765 2659 1816
rect 2711 1766 2723 1817
rect 2775 1767 2787 1818
rect 2839 1768 2851 1819
rect 2903 1769 2915 1820
rect 2967 1770 2979 1821
rect 3031 1771 3043 1822
rect 3095 1772 3107 1823
rect 3159 1772 3171 1824
rect 3223 1772 3372 1824
rect 3095 1771 3372 1772
rect 3031 1770 3372 1771
rect 2967 1769 3372 1770
rect 2903 1768 3372 1769
rect 2839 1767 3372 1768
rect 2775 1766 3372 1767
rect 2711 1765 3372 1766
rect 2647 1764 3372 1765
rect 2403 1759 3372 1764
rect 2403 1758 3107 1759
rect 2403 1757 3043 1758
rect 2403 1756 2979 1757
rect 2403 1755 2915 1756
rect 2403 1754 2851 1755
rect 2403 1753 2787 1754
rect 2403 1752 2467 1753
rect 2455 1701 2467 1752
rect 2519 1752 2723 1753
rect 2519 1701 2531 1752
rect 2455 1700 2531 1701
rect 2583 1751 2659 1752
rect 2583 1700 2595 1751
rect 2403 1699 2595 1700
rect 2647 1700 2659 1751
rect 2711 1701 2723 1752
rect 2775 1702 2787 1753
rect 2839 1703 2851 1754
rect 2903 1704 2915 1755
rect 2967 1705 2979 1756
rect 3031 1706 3043 1757
rect 3095 1707 3107 1758
rect 3159 1707 3171 1759
rect 3223 1707 3372 1759
rect 3095 1706 3372 1707
rect 3031 1705 3372 1706
rect 2967 1704 3372 1705
rect 2903 1703 3372 1704
rect 2839 1702 3372 1703
rect 2775 1701 3372 1702
rect 2711 1700 3372 1701
rect 2647 1699 3372 1700
rect 2403 1694 3372 1699
rect 2403 1693 3107 1694
rect 2403 1692 3043 1693
rect 2403 1691 2979 1692
rect 2403 1690 2915 1691
rect 2403 1689 2851 1690
rect 2403 1688 2787 1689
rect 2403 1686 2467 1688
rect 2455 1636 2467 1686
rect 2519 1687 2723 1688
rect 2519 1636 2531 1687
rect 2455 1635 2531 1636
rect 2583 1686 2659 1687
rect 2583 1635 2595 1686
rect 2455 1634 2595 1635
rect 2647 1635 2659 1686
rect 2711 1636 2723 1687
rect 2775 1637 2787 1688
rect 2839 1638 2851 1689
rect 2903 1639 2915 1690
rect 2967 1640 2979 1691
rect 3031 1641 3043 1692
rect 3095 1642 3107 1693
rect 3159 1642 3171 1694
rect 3223 1642 3372 1694
rect 3095 1641 3372 1642
rect 3031 1640 3372 1641
rect 2967 1639 3372 1640
rect 2903 1638 3372 1639
rect 2839 1637 3372 1638
rect 2775 1636 3372 1637
rect 2711 1635 3372 1636
rect 2647 1634 3372 1635
rect 2403 1629 3372 1634
rect 2403 1628 3107 1629
rect 2403 1627 3043 1628
rect 2403 1626 2979 1627
rect 2403 1625 2915 1626
rect 2403 1624 2851 1625
rect 2403 1623 2787 1624
rect 2403 1622 2723 1623
rect 2403 1620 2467 1622
tri 2084 1609 2085 1610 sw
rect 100 1568 2085 1609
tri 2085 1568 2126 1609 sw
tri 2362 1568 2403 1609 se
rect 2455 1570 2467 1620
rect 2519 1570 2531 1622
rect 2583 1621 2659 1622
rect 2583 1570 2595 1621
rect 2455 1569 2595 1570
rect 2647 1570 2659 1621
rect 2711 1571 2723 1622
rect 2775 1572 2787 1623
rect 2839 1573 2851 1624
rect 2903 1574 2915 1625
rect 2967 1575 2979 1626
rect 3031 1576 3043 1627
rect 3095 1577 3107 1628
rect 3159 1577 3171 1629
rect 3223 1577 3372 1629
rect 3095 1576 3372 1577
rect 3031 1575 3372 1576
rect 2967 1574 3372 1575
rect 2903 1573 3372 1574
rect 2839 1572 3372 1573
rect 2775 1571 3372 1572
rect 2711 1570 3372 1571
rect 2647 1569 3372 1570
rect 2455 1568 3372 1569
rect 100 1564 2126 1568
tri 2126 1564 2130 1568 sw
tri 2358 1564 2362 1568 se
rect 2362 1564 3372 1568
rect 100 1563 2130 1564
tri 2130 1563 2131 1564 sw
tri 2357 1563 2358 1564 se
rect 2358 1563 3107 1564
rect 100 1562 2131 1563
tri 2131 1562 2132 1563 sw
tri 2356 1562 2357 1563 se
rect 2357 1562 3043 1563
rect 100 1561 2132 1562
tri 2132 1561 2133 1562 sw
tri 2355 1561 2356 1562 se
rect 2356 1561 2979 1562
rect 100 1560 2133 1561
tri 2133 1560 2134 1561 sw
tri 2354 1560 2355 1561 se
rect 2355 1560 2915 1561
rect 100 1559 2134 1560
tri 2134 1559 2135 1560 sw
tri 2353 1559 2354 1560 se
rect 2354 1559 2851 1560
rect 100 1558 2135 1559
tri 2135 1558 2136 1559 sw
tri 2352 1558 2353 1559 se
rect 2353 1558 2787 1559
rect 100 1557 2136 1558
tri 2136 1557 2137 1558 sw
tri 2351 1557 2352 1558 se
rect 2352 1557 2723 1558
rect 100 1556 2137 1557
tri 2137 1556 2138 1557 sw
tri 2350 1556 2351 1557 se
rect 2351 1556 2531 1557
rect 100 1554 2138 1556
tri 2138 1554 2140 1556 sw
tri 2348 1554 2350 1556 se
rect 2350 1554 2467 1556
rect 100 1531 2140 1554
tri 2140 1531 2163 1554 sw
tri 2325 1531 2348 1554 se
rect 2348 1531 2403 1554
rect 100 1502 2403 1531
rect 2455 1504 2467 1554
rect 2519 1505 2531 1556
rect 2583 1556 2659 1557
rect 2583 1505 2595 1556
rect 2519 1504 2595 1505
rect 2647 1505 2659 1556
rect 2711 1506 2723 1557
rect 2775 1507 2787 1558
rect 2839 1508 2851 1559
rect 2903 1509 2915 1560
rect 2967 1510 2979 1561
rect 3031 1511 3043 1562
rect 3095 1512 3107 1563
rect 3159 1512 3171 1564
rect 3223 1512 3372 1564
rect 3095 1511 3372 1512
rect 3031 1510 3372 1511
rect 2967 1509 3372 1510
rect 2903 1508 3372 1509
rect 2839 1507 3372 1508
rect 2775 1506 3372 1507
rect 2711 1505 3372 1506
rect 2647 1504 3372 1505
rect 2455 1502 3372 1504
rect 100 1499 3372 1502
rect 100 1498 3107 1499
rect 100 1497 3043 1498
rect 100 1496 2979 1497
rect 100 1495 2915 1496
rect 100 1494 2851 1495
rect 100 1493 2787 1494
rect 100 1492 2723 1493
rect 100 1490 2531 1492
rect 100 1488 2467 1490
rect 100 1436 1939 1488
rect 1991 1436 2006 1488
rect 2058 1436 2073 1488
rect 2125 1436 2139 1488
rect 2191 1436 2205 1488
rect 2257 1436 2271 1488
rect 2323 1436 2337 1488
rect 2389 1436 2403 1488
rect 2455 1438 2467 1488
rect 2519 1440 2531 1490
rect 2583 1491 2659 1492
rect 2583 1440 2595 1491
rect 2519 1439 2595 1440
rect 2647 1440 2659 1491
rect 2711 1441 2723 1492
rect 2775 1442 2787 1493
rect 2839 1443 2851 1494
rect 2903 1444 2915 1495
rect 2967 1445 2979 1496
rect 3031 1446 3043 1497
rect 3095 1447 3107 1498
rect 3159 1447 3171 1499
rect 3223 1447 3372 1499
rect 3095 1446 3372 1447
rect 3031 1445 3372 1446
rect 2967 1444 3372 1445
rect 2903 1443 3372 1444
rect 2839 1442 3372 1443
rect 2775 1441 3372 1442
rect 2711 1440 3372 1441
rect 2647 1439 3372 1440
rect 2519 1438 3372 1439
rect 2455 1436 3372 1438
rect 100 1434 3372 1436
rect 100 1433 3107 1434
rect 100 1432 3043 1433
rect 100 1431 2979 1432
rect 100 1430 2915 1431
rect 100 1429 2851 1430
rect 100 1428 2787 1429
rect 100 1427 2723 1428
rect 100 1426 2659 1427
rect 100 1424 2531 1426
rect 100 1372 1939 1424
rect 1991 1372 2005 1424
rect 2057 1372 2071 1424
rect 2123 1372 2137 1424
rect 2189 1372 2203 1424
rect 2255 1372 2269 1424
rect 2321 1372 2335 1424
rect 2387 1372 2401 1424
rect 2453 1372 2467 1424
rect 2519 1374 2531 1424
rect 2583 1374 2595 1426
rect 2647 1375 2659 1426
rect 2711 1376 2723 1427
rect 2775 1377 2787 1428
rect 2839 1378 2851 1429
rect 2903 1379 2915 1430
rect 2967 1380 2979 1431
rect 3031 1381 3043 1432
rect 3095 1382 3107 1433
rect 3159 1382 3171 1434
rect 3223 1382 3372 1434
rect 3095 1381 3372 1382
rect 3031 1380 3372 1381
rect 2967 1379 3372 1380
rect 2903 1378 3372 1379
rect 2839 1377 3372 1378
rect 2775 1376 3372 1377
rect 2711 1375 3372 1376
rect 2647 1374 3372 1375
rect 2519 1372 3372 1374
rect 100 1369 3372 1372
rect 100 1368 3107 1369
rect 100 1367 3043 1368
rect 100 1366 2979 1367
rect 100 1365 2915 1366
rect 100 1364 2851 1365
rect 100 1363 2787 1364
rect 100 1362 2723 1363
rect 100 1361 2659 1362
rect 100 1360 2595 1361
rect 100 1308 1939 1360
rect 1991 1308 2005 1360
rect 2057 1308 2071 1360
rect 2123 1308 2137 1360
rect 2189 1308 2203 1360
rect 2255 1308 2269 1360
rect 2321 1308 2335 1360
rect 2387 1308 2401 1360
rect 2453 1308 2466 1360
rect 2518 1308 2531 1360
rect 2583 1309 2595 1360
rect 2647 1310 2659 1361
rect 2711 1311 2723 1362
rect 2775 1312 2787 1363
rect 2839 1313 2851 1364
rect 2903 1314 2915 1365
rect 2967 1315 2979 1366
rect 3031 1316 3043 1367
rect 3095 1317 3107 1368
rect 3159 1317 3171 1369
rect 3223 1317 3372 1369
rect 3095 1316 3372 1317
rect 3031 1315 3372 1316
rect 2967 1314 3372 1315
rect 2903 1313 3372 1314
rect 2839 1312 3372 1313
rect 2775 1311 3372 1312
rect 2711 1310 3372 1311
rect 2647 1309 3372 1310
rect 2583 1308 3372 1309
rect 100 1304 3372 1308
rect 100 1303 3107 1304
rect 100 1302 3043 1303
rect 100 1301 2979 1302
rect 100 1300 2915 1301
rect 100 1299 2851 1300
rect 100 1298 2787 1299
rect 100 1297 2723 1298
rect 100 1296 2659 1297
rect 100 1244 1939 1296
rect 1991 1244 2005 1296
rect 2057 1244 2071 1296
rect 2123 1244 2137 1296
rect 2189 1244 2203 1296
rect 2255 1244 2269 1296
rect 2321 1244 2335 1296
rect 2387 1244 2400 1296
rect 2452 1244 2465 1296
rect 2517 1244 2530 1296
rect 2582 1244 2595 1296
rect 2647 1245 2659 1296
rect 2711 1246 2723 1297
rect 2775 1247 2787 1298
rect 2839 1248 2851 1299
rect 2903 1249 2915 1300
rect 2967 1250 2979 1301
rect 3031 1251 3043 1302
rect 3095 1252 3107 1303
rect 3159 1252 3171 1304
rect 3223 1252 3372 1304
rect 3095 1251 3372 1252
rect 3031 1250 3372 1251
rect 2967 1249 3372 1250
rect 2903 1248 3372 1249
rect 2839 1247 3372 1248
rect 2775 1246 3372 1247
rect 2711 1245 3372 1246
rect 2647 1244 3372 1245
rect 100 1239 3372 1244
rect 100 1238 3107 1239
rect 100 1237 3043 1238
rect 100 1236 2979 1237
rect 100 1235 2915 1236
rect 100 1234 2851 1235
rect 100 1233 2787 1234
rect 100 1232 2723 1233
rect 100 1180 1939 1232
rect 1991 1180 2005 1232
rect 2057 1180 2071 1232
rect 2123 1180 2137 1232
rect 2189 1180 2203 1232
rect 2255 1180 2269 1232
rect 2321 1180 2334 1232
rect 2386 1180 2399 1232
rect 2451 1180 2464 1232
rect 2516 1180 2529 1232
rect 2581 1180 2594 1232
rect 2646 1180 2659 1232
rect 2711 1181 2723 1232
rect 2775 1182 2787 1233
rect 2839 1183 2851 1234
rect 2903 1184 2915 1235
rect 2967 1185 2979 1236
rect 3031 1186 3043 1237
rect 3095 1187 3107 1238
rect 3159 1187 3171 1239
rect 3223 1187 3372 1239
rect 3095 1186 3372 1187
rect 3031 1185 3372 1186
rect 2967 1184 3372 1185
rect 2903 1183 3372 1184
rect 2839 1182 3372 1183
rect 2775 1181 3372 1182
rect 2711 1180 3372 1181
rect 100 1174 3372 1180
rect 100 1173 3107 1174
rect 100 1172 3043 1173
rect 100 1171 2979 1172
rect 100 1170 2915 1171
rect 100 1169 2851 1170
rect 100 1168 2787 1169
rect 100 1116 1939 1168
rect 1991 1116 2005 1168
rect 2057 1116 2071 1168
rect 2123 1116 2137 1168
rect 2189 1116 2203 1168
rect 2255 1116 2268 1168
rect 2320 1116 2333 1168
rect 2385 1116 2398 1168
rect 2450 1116 2463 1168
rect 2515 1116 2528 1168
rect 2580 1116 2593 1168
rect 2645 1116 2658 1168
rect 2710 1116 2723 1168
rect 2775 1117 2787 1168
rect 2839 1118 2851 1169
rect 2903 1119 2915 1170
rect 2967 1120 2979 1171
rect 3031 1121 3043 1172
rect 3095 1122 3107 1173
rect 3159 1122 3171 1174
rect 3223 1122 3372 1174
rect 3095 1121 3372 1122
rect 3031 1120 3372 1121
rect 2967 1119 3372 1120
rect 2903 1118 3372 1119
rect 2839 1117 3372 1118
rect 2775 1116 3372 1117
rect 100 1109 3372 1116
rect 100 1108 3107 1109
rect 100 1107 3043 1108
rect 100 1106 2979 1107
rect 100 1105 2915 1106
rect 100 1104 2851 1105
rect 100 1052 1939 1104
rect 1991 1052 2005 1104
rect 2057 1052 2071 1104
rect 2123 1052 2137 1104
rect 2189 1052 2202 1104
rect 2254 1052 2267 1104
rect 2319 1052 2332 1104
rect 2384 1052 2397 1104
rect 2449 1052 2462 1104
rect 2514 1052 2527 1104
rect 2579 1052 2592 1104
rect 2644 1052 2657 1104
rect 2709 1052 2722 1104
rect 2774 1052 2787 1104
rect 2839 1053 2851 1104
rect 2903 1054 2915 1105
rect 2967 1055 2979 1106
rect 3031 1056 3043 1107
rect 3095 1057 3107 1108
rect 3159 1057 3171 1109
rect 3223 1057 3372 1109
rect 3095 1056 3372 1057
rect 3031 1055 3372 1056
rect 2967 1054 3372 1055
rect 2903 1053 3372 1054
rect 2839 1052 3372 1053
rect 100 1044 3372 1052
rect 100 1043 3107 1044
rect 100 1042 3043 1043
rect 100 1041 2979 1042
rect 100 1040 2915 1041
rect 100 988 1939 1040
rect 1991 988 2005 1040
rect 2057 988 2071 1040
rect 2123 988 2136 1040
rect 2188 988 2201 1040
rect 2253 988 2266 1040
rect 2318 988 2331 1040
rect 2383 988 2396 1040
rect 2448 988 2461 1040
rect 2513 988 2526 1040
rect 2578 988 2591 1040
rect 2643 988 2656 1040
rect 2708 988 2721 1040
rect 2773 988 2786 1040
rect 2838 988 2851 1040
rect 2903 989 2915 1040
rect 2967 990 2979 1041
rect 3031 991 3043 1042
rect 3095 992 3107 1043
rect 3159 992 3171 1044
rect 3223 1018 3372 1044
rect 3578 1850 3608 1902
rect 3660 1850 3690 1902
rect 3742 1850 3772 1902
rect 3824 1850 4350 1902
rect 4402 1850 4432 1902
rect 4484 1850 4514 1902
rect 4566 1850 4596 1902
rect 4648 1850 5174 1902
rect 5226 1850 5256 1902
rect 5308 1850 5338 1902
rect 5390 1850 5420 1902
rect 5472 1850 5998 1902
rect 6050 1850 6080 1902
rect 6132 1850 6162 1902
rect 6214 1850 6244 1902
rect 6296 1850 6822 1902
rect 6874 1850 6904 1902
rect 6956 1850 6986 1902
rect 7038 1850 7068 1902
rect 7120 1850 7936 1902
rect 7988 1850 8018 1902
rect 8070 1850 8100 1902
rect 8152 1850 8182 1902
rect 8234 1850 8760 1902
rect 8812 1850 8842 1902
rect 8894 1850 8924 1902
rect 8976 1850 9006 1902
rect 9058 1850 9584 1902
rect 9636 1850 9666 1902
rect 9718 1850 9748 1902
rect 9800 1850 9830 1902
rect 9882 1850 10408 1902
rect 10460 1850 10490 1902
rect 10542 1850 10572 1902
rect 10624 1850 10654 1902
rect 10706 1850 10707 1902
rect 3526 1838 10707 1850
rect 3526 1834 4350 1838
rect 3578 1782 3608 1834
rect 3660 1782 3690 1834
rect 3742 1782 3772 1834
rect 3824 1786 4350 1834
rect 4402 1786 4432 1838
rect 4484 1786 4514 1838
rect 4566 1786 4596 1838
rect 4648 1786 5174 1838
rect 5226 1786 5256 1838
rect 5308 1786 5338 1838
rect 5390 1786 5420 1838
rect 5472 1786 5998 1838
rect 6050 1786 6080 1838
rect 6132 1786 6162 1838
rect 6214 1786 6244 1838
rect 6296 1786 6822 1838
rect 6874 1786 6904 1838
rect 6956 1786 6986 1838
rect 7038 1786 7068 1838
rect 7120 1786 7936 1838
rect 7988 1786 8018 1838
rect 8070 1786 8100 1838
rect 8152 1786 8182 1838
rect 8234 1786 8760 1838
rect 8812 1786 8842 1838
rect 8894 1786 8924 1838
rect 8976 1786 9006 1838
rect 9058 1786 9584 1838
rect 9636 1786 9666 1838
rect 9718 1786 9748 1838
rect 9800 1786 9830 1838
rect 9882 1786 10408 1838
rect 10460 1786 10490 1838
rect 10542 1786 10572 1838
rect 10624 1786 10654 1838
rect 10706 1786 10707 1838
rect 3824 1782 10707 1786
rect 3526 1774 10707 1782
rect 3526 1766 4350 1774
rect 3578 1714 3608 1766
rect 3660 1714 3690 1766
rect 3742 1714 3772 1766
rect 3824 1722 4350 1766
rect 4402 1722 4432 1774
rect 4484 1722 4514 1774
rect 4566 1722 4596 1774
rect 4648 1722 5174 1774
rect 5226 1722 5256 1774
rect 5308 1722 5338 1774
rect 5390 1722 5420 1774
rect 5472 1722 5998 1774
rect 6050 1722 6080 1774
rect 6132 1722 6162 1774
rect 6214 1722 6244 1774
rect 6296 1722 6822 1774
rect 6874 1722 6904 1774
rect 6956 1722 6986 1774
rect 7038 1722 7068 1774
rect 7120 1722 7936 1774
rect 7988 1722 8018 1774
rect 8070 1722 8100 1774
rect 8152 1722 8182 1774
rect 8234 1722 8760 1774
rect 8812 1722 8842 1774
rect 8894 1722 8924 1774
rect 8976 1722 9006 1774
rect 9058 1722 9584 1774
rect 9636 1722 9666 1774
rect 9718 1722 9748 1774
rect 9800 1722 9830 1774
rect 9882 1722 10408 1774
rect 10460 1722 10490 1774
rect 10542 1722 10572 1774
rect 10624 1722 10654 1774
rect 10706 1722 10707 1774
rect 3824 1714 10707 1722
rect 3526 1710 10707 1714
rect 3526 1698 4350 1710
rect 3578 1646 3608 1698
rect 3660 1646 3690 1698
rect 3742 1646 3772 1698
rect 3824 1658 4350 1698
rect 4402 1658 4432 1710
rect 4484 1658 4514 1710
rect 4566 1658 4596 1710
rect 4648 1658 5174 1710
rect 5226 1658 5256 1710
rect 5308 1658 5338 1710
rect 5390 1658 5420 1710
rect 5472 1658 5998 1710
rect 6050 1658 6080 1710
rect 6132 1658 6162 1710
rect 6214 1658 6244 1710
rect 6296 1658 6822 1710
rect 6874 1658 6904 1710
rect 6956 1658 6986 1710
rect 7038 1658 7068 1710
rect 7120 1658 7936 1710
rect 7988 1658 8018 1710
rect 8070 1658 8100 1710
rect 8152 1658 8182 1710
rect 8234 1658 8760 1710
rect 8812 1658 8842 1710
rect 8894 1658 8924 1710
rect 8976 1658 9006 1710
rect 9058 1658 9584 1710
rect 9636 1658 9666 1710
rect 9718 1658 9748 1710
rect 9800 1658 9830 1710
rect 9882 1658 10408 1710
rect 10460 1658 10490 1710
rect 10542 1658 10572 1710
rect 10624 1658 10654 1710
rect 10706 1658 10707 1710
rect 3824 1646 10707 1658
rect 3526 1630 4350 1646
rect 3578 1578 3608 1630
rect 3660 1578 3690 1630
rect 3742 1578 3772 1630
rect 3824 1594 4350 1630
rect 4402 1594 4432 1646
rect 4484 1594 4514 1646
rect 4566 1594 4596 1646
rect 4648 1594 5174 1646
rect 5226 1594 5256 1646
rect 5308 1594 5338 1646
rect 5390 1594 5420 1646
rect 5472 1594 5998 1646
rect 6050 1594 6080 1646
rect 6132 1594 6162 1646
rect 6214 1594 6244 1646
rect 6296 1594 6822 1646
rect 6874 1594 6904 1646
rect 6956 1594 6986 1646
rect 7038 1594 7068 1646
rect 7120 1594 7936 1646
rect 7988 1594 8018 1646
rect 8070 1594 8100 1646
rect 8152 1594 8182 1646
rect 8234 1594 8760 1646
rect 8812 1594 8842 1646
rect 8894 1594 8924 1646
rect 8976 1594 9006 1646
rect 9058 1594 9584 1646
rect 9636 1594 9666 1646
rect 9718 1594 9748 1646
rect 9800 1594 9830 1646
rect 9882 1594 10408 1646
rect 10460 1594 10490 1646
rect 10542 1594 10572 1646
rect 10624 1594 10654 1646
rect 10706 1594 10707 1646
rect 3824 1582 10707 1594
rect 3824 1578 4350 1582
rect 3526 1562 4350 1578
rect 3578 1510 3608 1562
rect 3660 1510 3690 1562
rect 3742 1510 3772 1562
rect 3824 1530 4350 1562
rect 4402 1530 4432 1582
rect 4484 1530 4514 1582
rect 4566 1530 4596 1582
rect 4648 1530 5174 1582
rect 5226 1530 5256 1582
rect 5308 1530 5338 1582
rect 5390 1530 5420 1582
rect 5472 1530 5998 1582
rect 6050 1530 6080 1582
rect 6132 1530 6162 1582
rect 6214 1530 6244 1582
rect 6296 1530 6822 1582
rect 6874 1530 6904 1582
rect 6956 1530 6986 1582
rect 7038 1530 7068 1582
rect 7120 1530 7936 1582
rect 7988 1530 8018 1582
rect 8070 1530 8100 1582
rect 8152 1530 8182 1582
rect 8234 1530 8760 1582
rect 8812 1530 8842 1582
rect 8894 1530 8924 1582
rect 8976 1530 9006 1582
rect 9058 1530 9584 1582
rect 9636 1530 9666 1582
rect 9718 1530 9748 1582
rect 9800 1530 9830 1582
rect 9882 1530 10408 1582
rect 10460 1530 10490 1582
rect 10542 1530 10572 1582
rect 10624 1530 10654 1582
rect 10706 1530 10707 1582
rect 3824 1518 10707 1530
rect 3824 1510 4350 1518
rect 3526 1494 4350 1510
rect 3578 1442 3608 1494
rect 3660 1442 3690 1494
rect 3742 1442 3772 1494
rect 3824 1466 4350 1494
rect 4402 1466 4432 1518
rect 4484 1466 4514 1518
rect 4566 1466 4596 1518
rect 4648 1466 5174 1518
rect 5226 1466 5256 1518
rect 5308 1466 5338 1518
rect 5390 1466 5420 1518
rect 5472 1466 5998 1518
rect 6050 1466 6080 1518
rect 6132 1466 6162 1518
rect 6214 1466 6244 1518
rect 6296 1466 6822 1518
rect 6874 1466 6904 1518
rect 6956 1466 6986 1518
rect 7038 1466 7068 1518
rect 7120 1466 7936 1518
rect 7988 1466 8018 1518
rect 8070 1466 8100 1518
rect 8152 1466 8182 1518
rect 8234 1466 8760 1518
rect 8812 1466 8842 1518
rect 8894 1466 8924 1518
rect 8976 1466 9006 1518
rect 9058 1466 9584 1518
rect 9636 1466 9666 1518
rect 9718 1466 9748 1518
rect 9800 1466 9830 1518
rect 9882 1466 10408 1518
rect 10460 1466 10490 1518
rect 10542 1466 10572 1518
rect 10624 1466 10654 1518
rect 10706 1466 10707 1518
rect 3824 1454 10707 1466
rect 3824 1442 4350 1454
rect 3526 1426 4350 1442
rect 3578 1374 3608 1426
rect 3660 1374 3690 1426
rect 3742 1374 3772 1426
rect 3824 1402 4350 1426
rect 4402 1402 4432 1454
rect 4484 1402 4514 1454
rect 4566 1402 4596 1454
rect 4648 1402 5174 1454
rect 5226 1402 5256 1454
rect 5308 1402 5338 1454
rect 5390 1402 5420 1454
rect 5472 1402 5998 1454
rect 6050 1402 6080 1454
rect 6132 1402 6162 1454
rect 6214 1402 6244 1454
rect 6296 1402 6822 1454
rect 6874 1402 6904 1454
rect 6956 1402 6986 1454
rect 7038 1402 7068 1454
rect 7120 1402 7936 1454
rect 7988 1402 8018 1454
rect 8070 1402 8100 1454
rect 8152 1402 8182 1454
rect 8234 1402 8760 1454
rect 8812 1402 8842 1454
rect 8894 1402 8924 1454
rect 8976 1402 9006 1454
rect 9058 1402 9584 1454
rect 9636 1402 9666 1454
rect 9718 1402 9748 1454
rect 9800 1402 9830 1454
rect 9882 1402 10408 1454
rect 10460 1402 10490 1454
rect 10542 1402 10572 1454
rect 10624 1402 10654 1454
rect 10706 1402 10707 1454
rect 3824 1390 10707 1402
rect 3824 1374 4350 1390
rect 3526 1358 4350 1374
rect 3578 1306 3608 1358
rect 3660 1306 3690 1358
rect 3742 1306 3772 1358
rect 3824 1338 4350 1358
rect 4402 1338 4432 1390
rect 4484 1338 4514 1390
rect 4566 1338 4596 1390
rect 4648 1338 5174 1390
rect 5226 1338 5256 1390
rect 5308 1338 5338 1390
rect 5390 1338 5420 1390
rect 5472 1338 5998 1390
rect 6050 1338 6080 1390
rect 6132 1338 6162 1390
rect 6214 1338 6244 1390
rect 6296 1338 6822 1390
rect 6874 1338 6904 1390
rect 6956 1338 6986 1390
rect 7038 1338 7068 1390
rect 7120 1338 7936 1390
rect 7988 1338 8018 1390
rect 8070 1338 8100 1390
rect 8152 1338 8182 1390
rect 8234 1338 8760 1390
rect 8812 1338 8842 1390
rect 8894 1338 8924 1390
rect 8976 1338 9006 1390
rect 9058 1338 9584 1390
rect 9636 1338 9666 1390
rect 9718 1338 9748 1390
rect 9800 1338 9830 1390
rect 9882 1338 10408 1390
rect 10460 1338 10490 1390
rect 10542 1338 10572 1390
rect 10624 1338 10654 1390
rect 10706 1338 10707 1390
rect 3824 1326 10707 1338
rect 3824 1306 4350 1326
rect 3526 1289 4350 1306
rect 3578 1237 3608 1289
rect 3660 1237 3690 1289
rect 3742 1237 3772 1289
rect 3824 1274 4350 1289
rect 4402 1274 4432 1326
rect 4484 1274 4514 1326
rect 4566 1274 4596 1326
rect 4648 1274 5174 1326
rect 5226 1274 5256 1326
rect 5308 1274 5338 1326
rect 5390 1274 5420 1326
rect 5472 1274 5998 1326
rect 6050 1274 6080 1326
rect 6132 1274 6162 1326
rect 6214 1274 6244 1326
rect 6296 1274 6822 1326
rect 6874 1274 6904 1326
rect 6956 1274 6986 1326
rect 7038 1274 7068 1326
rect 7120 1274 7936 1326
rect 7988 1274 8018 1326
rect 8070 1274 8100 1326
rect 8152 1274 8182 1326
rect 8234 1274 8760 1326
rect 8812 1274 8842 1326
rect 8894 1274 8924 1326
rect 8976 1274 9006 1326
rect 9058 1274 9584 1326
rect 9636 1274 9666 1326
rect 9718 1274 9748 1326
rect 9800 1274 9830 1326
rect 9882 1274 10408 1326
rect 10460 1274 10490 1326
rect 10542 1274 10572 1326
rect 10624 1274 10654 1326
rect 10706 1274 10707 1326
rect 3824 1262 10707 1274
rect 3824 1237 4350 1262
rect 3526 1220 4350 1237
rect 3578 1168 3608 1220
rect 3660 1168 3690 1220
rect 3742 1168 3772 1220
rect 3824 1210 4350 1220
rect 4402 1210 4432 1262
rect 4484 1210 4514 1262
rect 4566 1210 4596 1262
rect 4648 1210 5174 1262
rect 5226 1210 5256 1262
rect 5308 1210 5338 1262
rect 5390 1210 5420 1262
rect 5472 1210 5998 1262
rect 6050 1210 6080 1262
rect 6132 1210 6162 1262
rect 6214 1210 6244 1262
rect 6296 1210 6822 1262
rect 6874 1210 6904 1262
rect 6956 1210 6986 1262
rect 7038 1210 7068 1262
rect 7120 1210 7936 1262
rect 7988 1210 8018 1262
rect 8070 1210 8100 1262
rect 8152 1210 8182 1262
rect 8234 1210 8760 1262
rect 8812 1210 8842 1262
rect 8894 1210 8924 1262
rect 8976 1210 9006 1262
rect 9058 1210 9584 1262
rect 9636 1210 9666 1262
rect 9718 1210 9748 1262
rect 9800 1210 9830 1262
rect 9882 1210 10408 1262
rect 10460 1210 10490 1262
rect 10542 1210 10572 1262
rect 10624 1210 10654 1262
rect 10706 1210 10707 1262
rect 3824 1198 10707 1210
rect 3824 1168 4350 1198
rect 3526 1151 4350 1168
rect 3578 1099 3608 1151
rect 3660 1099 3690 1151
rect 3742 1099 3772 1151
rect 3824 1146 4350 1151
rect 4402 1146 4432 1198
rect 4484 1146 4514 1198
rect 4566 1146 4596 1198
rect 4648 1146 5174 1198
rect 5226 1146 5256 1198
rect 5308 1146 5338 1198
rect 5390 1146 5420 1198
rect 5472 1146 5998 1198
rect 6050 1146 6080 1198
rect 6132 1146 6162 1198
rect 6214 1146 6244 1198
rect 6296 1146 6822 1198
rect 6874 1146 6904 1198
rect 6956 1146 6986 1198
rect 7038 1146 7068 1198
rect 7120 1146 7936 1198
rect 7988 1146 8018 1198
rect 8070 1146 8100 1198
rect 8152 1146 8182 1198
rect 8234 1146 8760 1198
rect 8812 1146 8842 1198
rect 8894 1146 8924 1198
rect 8976 1146 9006 1198
rect 9058 1146 9584 1198
rect 9636 1146 9666 1198
rect 9718 1146 9748 1198
rect 9800 1146 9830 1198
rect 9882 1146 10408 1198
rect 10460 1146 10490 1198
rect 10542 1146 10572 1198
rect 10624 1146 10654 1198
rect 10706 1146 10707 1198
rect 3824 1134 10707 1146
rect 3824 1099 4350 1134
rect 3526 1082 4350 1099
rect 4402 1082 4432 1134
rect 4484 1082 4514 1134
rect 4566 1082 4596 1134
rect 4648 1082 5174 1134
rect 5226 1082 5256 1134
rect 5308 1082 5338 1134
rect 5390 1082 5420 1134
rect 5472 1082 5998 1134
rect 6050 1082 6080 1134
rect 6132 1082 6162 1134
rect 6214 1082 6244 1134
rect 6296 1082 6822 1134
rect 6874 1082 6904 1134
rect 6956 1082 6986 1134
rect 7038 1082 7068 1134
rect 7120 1082 7936 1134
rect 7988 1082 8018 1134
rect 8070 1082 8100 1134
rect 8152 1082 8182 1134
rect 8234 1082 8760 1134
rect 8812 1082 8842 1134
rect 8894 1082 8924 1134
rect 8976 1082 9006 1134
rect 9058 1082 9584 1134
rect 9636 1082 9666 1134
rect 9718 1082 9748 1134
rect 9800 1082 9830 1134
rect 9882 1082 10408 1134
rect 10460 1082 10490 1134
rect 10542 1082 10572 1134
rect 10624 1082 10654 1134
rect 10706 1082 10707 1134
rect 3578 1030 3608 1082
rect 3660 1030 3690 1082
rect 3742 1030 3772 1082
rect 3824 1070 10707 1082
rect 3824 1030 4350 1070
tri 3372 1018 3378 1024 sw
rect 3526 1023 4350 1030
tri 3526 1018 3531 1023 ne
rect 3531 1018 4350 1023
rect 4402 1018 4432 1070
rect 4484 1018 4514 1070
rect 4566 1018 4596 1070
rect 4648 1018 5174 1070
rect 5226 1018 5256 1070
rect 5308 1018 5338 1070
rect 5390 1018 5420 1070
rect 5472 1018 5998 1070
rect 6050 1018 6080 1070
rect 6132 1018 6162 1070
rect 6214 1018 6244 1070
rect 6296 1018 6822 1070
rect 6874 1018 6904 1070
rect 6956 1018 6986 1070
rect 7038 1018 7068 1070
rect 7120 1018 7936 1070
rect 7988 1018 8018 1070
rect 8070 1018 8100 1070
rect 8152 1018 8182 1070
rect 8234 1018 8760 1070
rect 8812 1018 8842 1070
rect 8894 1018 8924 1070
rect 8976 1018 9006 1070
rect 9058 1018 9584 1070
rect 9636 1018 9666 1070
rect 9718 1018 9748 1070
rect 9800 1018 9830 1070
rect 9882 1018 10408 1070
rect 10460 1018 10490 1070
rect 10542 1018 10572 1070
rect 10624 1018 10654 1070
rect 10706 1018 10707 1070
rect 3223 992 3378 1018
rect 3095 991 3378 992
rect 3031 990 3378 991
rect 2967 989 3378 990
rect 2903 988 3378 989
rect 100 979 3378 988
rect 100 978 3107 979
rect 100 977 3043 978
rect 100 976 2979 977
rect 100 924 1939 976
rect 1991 924 2005 976
rect 2057 924 2070 976
rect 2122 924 2135 976
rect 2187 924 2200 976
rect 2252 924 2265 976
rect 2317 924 2330 976
rect 2382 924 2395 976
rect 2447 924 2460 976
rect 2512 924 2525 976
rect 2577 924 2590 976
rect 2642 924 2655 976
rect 2707 924 2720 976
rect 2772 924 2785 976
rect 2837 924 2850 976
rect 2902 924 2915 976
rect 2967 925 2979 976
rect 3031 926 3043 977
rect 3095 927 3107 978
rect 3159 927 3171 979
rect 3223 966 3378 979
tri 3378 966 3430 1018 sw
tri 3531 966 3583 1018 ne
rect 3583 966 3590 1018
rect 3642 966 3678 1018
rect 3730 966 3766 1018
rect 3818 1006 10707 1018
rect 3818 966 4350 1006
rect 3223 954 3430 966
tri 3430 954 3442 966 sw
tri 3583 954 3595 966 ne
rect 3595 954 4350 966
rect 4402 954 4432 1006
rect 4484 954 4514 1006
rect 4566 954 4596 1006
rect 4648 954 5174 1006
rect 5226 954 5256 1006
rect 5308 954 5338 1006
rect 5390 954 5420 1006
rect 5472 954 5998 1006
rect 6050 954 6080 1006
rect 6132 954 6162 1006
rect 6214 954 6244 1006
rect 6296 954 6822 1006
rect 6874 954 6904 1006
rect 6956 954 6986 1006
rect 7038 954 7068 1006
rect 7120 954 7936 1006
rect 7988 954 8018 1006
rect 8070 954 8100 1006
rect 8152 954 8182 1006
rect 8234 954 8760 1006
rect 8812 954 8842 1006
rect 8894 954 8924 1006
rect 8976 954 9006 1006
rect 9058 954 9584 1006
rect 9636 954 9666 1006
rect 9718 954 9748 1006
rect 9800 954 9830 1006
rect 9882 954 10408 1006
rect 10460 954 10490 1006
rect 10542 954 10572 1006
rect 10624 954 10654 1006
rect 10706 954 10707 1006
rect 3223 953 3442 954
tri 3442 953 3443 954 sw
tri 3595 953 3596 954 ne
rect 3596 953 10707 954
rect 3223 927 3443 953
rect 3095 926 3443 927
rect 3031 925 3443 926
rect 2967 924 3443 925
rect 100 914 3443 924
rect 100 913 3107 914
rect 100 912 3043 913
rect 100 860 1939 912
rect 1991 860 2004 912
rect 2056 860 2069 912
rect 2121 860 2134 912
rect 2186 860 2199 912
rect 2251 860 2264 912
rect 2316 860 2329 912
rect 2381 860 2394 912
rect 2446 860 2459 912
rect 2511 860 2524 912
rect 2576 860 2589 912
rect 2641 860 2654 912
rect 2706 860 2719 912
rect 2771 860 2784 912
rect 2836 860 2849 912
rect 2901 860 2914 912
rect 2966 860 2979 912
rect 3031 861 3043 912
rect 3095 862 3107 913
rect 3159 862 3171 914
rect 3223 901 3443 914
tri 3443 901 3495 953 sw
tri 3596 901 3648 953 ne
rect 3648 901 3660 953
rect 3712 901 3766 953
rect 3818 942 10707 953
rect 3818 901 4350 942
rect 3223 890 3495 901
tri 3495 890 3506 901 sw
tri 3648 890 3659 901 ne
rect 3659 890 4350 901
rect 4402 890 4432 942
rect 4484 890 4514 942
rect 4566 890 4596 942
rect 4648 890 5174 942
rect 5226 890 5256 942
rect 5308 890 5338 942
rect 5390 890 5420 942
rect 5472 890 5998 942
rect 6050 890 6080 942
rect 6132 890 6162 942
rect 6214 890 6244 942
rect 6296 890 6822 942
rect 6874 890 6904 942
rect 6956 890 6986 942
rect 7038 890 7068 942
rect 7120 890 7936 942
rect 7988 890 8018 942
rect 8070 890 8100 942
rect 8152 890 8182 942
rect 8234 890 8760 942
rect 8812 890 8842 942
rect 8894 890 8924 942
rect 8976 890 9006 942
rect 9058 890 9584 942
rect 9636 890 9666 942
rect 9718 890 9748 942
rect 9800 890 9830 942
rect 9882 890 10408 942
rect 10460 890 10490 942
rect 10542 890 10572 942
rect 10624 890 10654 942
rect 10706 890 10707 942
rect 3223 878 3506 890
tri 3506 878 3518 890 sw
tri 3659 878 3671 890 ne
rect 3671 878 10707 890
rect 3223 870 3518 878
tri 3518 870 3526 878 sw
tri 3671 870 3679 878 ne
rect 3679 870 4350 878
rect 3223 867 3526 870
tri 3526 867 3529 870 sw
tri 3679 867 3682 870 ne
rect 3682 867 4350 870
rect 3223 862 3529 867
rect 3095 861 3529 862
rect 3031 860 3529 861
rect 100 849 3529 860
rect 100 848 3107 849
rect 100 796 1939 848
rect 1991 796 2004 848
rect 2056 796 2069 848
rect 2121 796 2134 848
rect 2186 796 2199 848
rect 2251 796 2264 848
rect 2316 796 2329 848
rect 2381 796 2394 848
rect 2446 796 2459 848
rect 2511 796 2524 848
rect 2576 796 2589 848
rect 2641 796 2654 848
rect 2706 796 2719 848
rect 2771 796 2784 848
rect 2836 796 2849 848
rect 2901 796 2914 848
rect 2966 796 2979 848
rect 100 784 2979 796
rect 3095 797 3107 848
rect 3159 797 3171 849
rect 3223 815 3529 849
tri 3529 815 3581 867 sw
tri 3682 815 3734 867 ne
rect 3734 815 3753 867
rect 3805 826 4350 867
rect 4402 826 4432 878
rect 4484 826 4514 878
rect 4566 826 4596 878
rect 4648 826 5174 878
rect 5226 826 5256 878
rect 5308 826 5338 878
rect 5390 826 5420 878
rect 5472 826 5998 878
rect 6050 826 6080 878
rect 6132 826 6162 878
rect 6214 826 6244 878
rect 6296 826 6822 878
rect 6874 826 6904 878
rect 6956 826 6986 878
rect 7038 826 7068 878
rect 7120 826 7936 878
rect 7988 826 8018 878
rect 8070 826 8100 878
rect 8152 826 8182 878
rect 8234 826 8760 878
rect 8812 826 8842 878
rect 8894 826 8924 878
rect 8976 826 9006 878
rect 9058 826 9584 878
rect 9636 826 9666 878
rect 9718 826 9748 878
rect 9800 826 9830 878
rect 9882 826 10408 878
rect 10460 826 10490 878
rect 10542 826 10572 878
rect 10624 826 10654 878
rect 10706 826 10707 878
rect 3805 815 10707 826
rect 3223 814 3581 815
tri 3581 814 3582 815 sw
tri 3734 814 3735 815 ne
rect 3735 814 10707 815
rect 3223 797 3582 814
rect 3095 784 3582 797
rect 100 732 1939 784
rect 1991 732 2004 784
rect 2056 732 2069 784
rect 2121 732 2134 784
rect 2186 732 2199 784
rect 2251 732 2264 784
rect 2316 732 2329 784
rect 2381 732 2394 784
rect 2446 732 2459 784
rect 2511 732 2524 784
rect 2576 732 2589 784
rect 2641 732 2654 784
rect 2706 732 2719 784
rect 2771 732 2784 784
rect 2836 732 2849 784
rect 2901 732 2914 784
rect 2966 732 2979 784
rect 100 720 2979 732
rect 100 668 1939 720
rect 1991 668 2004 720
rect 2056 668 2069 720
rect 2121 668 2134 720
rect 2186 668 2199 720
rect 2251 668 2264 720
rect 2316 668 2329 720
rect 2381 668 2394 720
rect 2446 668 2459 720
rect 2511 668 2524 720
rect 2576 668 2589 720
rect 2641 668 2654 720
rect 2706 668 2719 720
rect 2771 668 2784 720
rect 2836 668 2849 720
rect 2901 668 2914 720
rect 2966 668 2979 720
rect 3159 732 3171 784
rect 3223 762 3582 784
tri 3582 762 3634 814 sw
tri 3735 762 3787 814 ne
rect 3787 762 4350 814
rect 4402 762 4432 814
rect 4484 762 4514 814
rect 4566 762 4596 814
rect 4648 762 5174 814
rect 5226 762 5256 814
rect 5308 762 5338 814
rect 5390 762 5420 814
rect 5472 762 5998 814
rect 6050 762 6080 814
rect 6132 762 6162 814
rect 6214 762 6244 814
rect 6296 762 6822 814
rect 6874 762 6904 814
rect 6956 762 6986 814
rect 7038 762 7068 814
rect 7120 762 7936 814
rect 7988 762 8018 814
rect 8070 762 8100 814
rect 8152 762 8182 814
rect 8234 762 8760 814
rect 8812 762 8842 814
rect 8894 762 8924 814
rect 8976 762 9006 814
rect 9058 762 9584 814
rect 9636 762 9666 814
rect 9718 762 9748 814
rect 9800 762 9830 814
rect 9882 762 10408 814
rect 10460 762 10490 814
rect 10542 762 10572 814
rect 10624 762 10654 814
rect 10706 762 10707 814
rect 3223 750 3634 762
tri 3634 750 3646 762 sw
tri 3787 750 3799 762 ne
rect 3799 750 10707 762
rect 3223 732 3646 750
rect 3159 717 3646 732
tri 3646 717 3679 750 sw
tri 3799 717 3832 750 ne
rect 3832 717 4350 750
rect 3159 698 3679 717
tri 3679 698 3698 717 sw
tri 3832 698 3851 717 ne
rect 3851 698 4350 717
rect 4402 698 4432 750
rect 4484 698 4514 750
rect 4566 698 4596 750
rect 4648 698 5174 750
rect 5226 698 5256 750
rect 5308 698 5338 750
rect 5390 698 5420 750
rect 5472 698 5998 750
rect 6050 698 6080 750
rect 6132 698 6162 750
rect 6214 698 6244 750
rect 6296 698 6822 750
rect 6874 698 6904 750
rect 6956 698 6986 750
rect 7038 698 7068 750
rect 7120 698 7936 750
rect 7988 698 8018 750
rect 8070 698 8100 750
rect 8152 698 8182 750
rect 8234 698 8760 750
rect 8812 698 8842 750
rect 8894 698 8924 750
rect 8976 698 9006 750
rect 9058 698 9584 750
rect 9636 698 9666 750
rect 9718 698 9748 750
rect 9800 698 9830 750
rect 9882 698 10408 750
rect 10460 698 10490 750
rect 10542 698 10572 750
rect 10624 698 10654 750
rect 10706 698 10707 750
rect 3159 685 3698 698
tri 3698 685 3711 698 sw
tri 3851 685 3864 698 ne
rect 3864 685 10707 698
rect 3159 668 3711 685
rect 100 633 3711 668
tri 3711 633 3763 685 sw
tri 3864 633 3916 685 ne
rect 3916 633 4350 685
rect 4402 633 4432 685
rect 4484 633 4514 685
rect 4566 633 4596 685
rect 4648 633 5174 685
rect 5226 633 5256 685
rect 5308 633 5338 685
rect 5390 633 5420 685
rect 5472 633 5998 685
rect 6050 633 6080 685
rect 6132 633 6162 685
rect 6214 633 6244 685
rect 6296 633 6822 685
rect 6874 633 6904 685
rect 6956 633 6986 685
rect 7038 633 7068 685
rect 7120 633 7936 685
rect 7988 633 8018 685
rect 8070 633 8100 685
rect 8152 633 8182 685
rect 8234 633 8760 685
rect 8812 633 8842 685
rect 8894 633 8924 685
rect 8976 633 9006 685
rect 9058 633 9584 685
rect 9636 633 9666 685
rect 9718 633 9748 685
rect 9800 633 9830 685
rect 9882 633 10408 685
rect 10460 633 10490 685
rect 10542 633 10572 685
rect 10624 633 10654 685
rect 10706 633 10707 685
rect 100 620 3763 633
tri 3763 620 3776 633 sw
tri 3916 620 3929 633 ne
rect 3929 620 10707 633
rect 100 603 3776 620
tri 3776 603 3793 620 sw
tri 3929 603 3946 620 ne
rect 3946 603 4350 620
rect 100 568 3793 603
tri 3793 568 3828 603 sw
tri 3946 568 3981 603 ne
rect 3981 568 4350 603
rect 4402 568 4432 620
rect 4484 568 4514 620
rect 4566 568 4596 620
rect 4648 568 5174 620
rect 5226 568 5256 620
rect 5308 568 5338 620
rect 5390 568 5420 620
rect 5472 568 5998 620
rect 6050 568 6080 620
rect 6132 568 6162 620
rect 6214 568 6244 620
rect 6296 568 6822 620
rect 6874 568 6904 620
rect 6956 568 6986 620
rect 7038 568 7068 620
rect 7120 568 7936 620
rect 7988 568 8018 620
rect 8070 568 8100 620
rect 8152 568 8182 620
rect 8234 568 8760 620
rect 8812 568 8842 620
rect 8894 568 8924 620
rect 8976 568 9006 620
rect 9058 568 9584 620
rect 9636 568 9666 620
rect 9718 568 9748 620
rect 9800 568 9830 620
rect 9882 568 10408 620
rect 10460 568 10490 620
rect 10542 568 10572 620
rect 10624 568 10654 620
rect 10706 568 10707 620
rect 100 555 3828 568
tri 3828 555 3841 568 sw
tri 3981 555 3994 568 ne
rect 3994 555 10707 568
rect 100 503 3841 555
tri 3841 503 3893 555 sw
tri 3994 503 4046 555 ne
rect 4046 503 4350 555
rect 4402 503 4432 555
rect 4484 503 4514 555
rect 4566 503 4596 555
rect 4648 503 5174 555
rect 5226 503 5256 555
rect 5308 503 5338 555
rect 5390 503 5420 555
rect 5472 503 5998 555
rect 6050 503 6080 555
rect 6132 503 6162 555
rect 6214 503 6244 555
rect 6296 503 6822 555
rect 6874 503 6904 555
rect 6956 503 6986 555
rect 7038 503 7068 555
rect 7120 503 7936 555
rect 7988 503 8018 555
rect 8070 503 8100 555
rect 8152 503 8182 555
rect 8234 503 8760 555
rect 8812 503 8842 555
rect 8894 503 8924 555
rect 8976 503 9006 555
rect 9058 503 9584 555
rect 9636 503 9666 555
rect 9718 503 9748 555
rect 9800 503 9830 555
rect 9882 503 10408 555
rect 10460 503 10490 555
rect 10542 503 10572 555
rect 10624 503 10654 555
rect 10706 503 10707 555
rect 100 490 3893 503
tri 3893 490 3906 503 sw
tri 4046 490 4059 503 ne
rect 4059 490 10707 503
rect 100 450 3906 490
tri 3906 450 3946 490 sw
tri 4059 450 4099 490 ne
rect 4099 450 4350 490
rect 100 438 3946 450
tri 3946 438 3958 450 sw
tri 4099 438 4111 450 ne
rect 4111 438 4350 450
rect 4402 438 4432 490
rect 4484 438 4514 490
rect 4566 438 4596 490
rect 4648 438 5174 490
rect 5226 438 5256 490
rect 5308 438 5338 490
rect 5390 438 5420 490
rect 5472 438 5998 490
rect 6050 438 6080 490
rect 6132 438 6162 490
rect 6214 438 6244 490
rect 6296 438 6822 490
rect 6874 438 6904 490
rect 6956 438 6986 490
rect 7038 438 7068 490
rect 7120 438 7936 490
rect 7988 438 8018 490
rect 8070 438 8100 490
rect 8152 438 8182 490
rect 8234 438 8760 490
rect 8812 438 8842 490
rect 8894 438 8924 490
rect 8976 438 9006 490
rect 9058 438 9584 490
rect 9636 438 9666 490
rect 9718 438 9748 490
rect 9800 438 9830 490
rect 9882 438 10408 490
rect 10460 438 10490 490
rect 10542 438 10572 490
rect 10624 438 10654 490
rect 10706 438 10707 490
rect 100 425 3958 438
tri 3958 425 3971 438 sw
tri 4111 425 4124 438 ne
rect 4124 425 10707 438
rect 100 373 3971 425
tri 3971 373 4023 425 sw
tri 4124 373 4176 425 ne
rect 4176 373 4350 425
rect 4402 373 4432 425
rect 4484 373 4514 425
rect 4566 373 4596 425
rect 4648 373 5174 425
rect 5226 373 5256 425
rect 5308 373 5338 425
rect 5390 373 5420 425
rect 5472 373 5998 425
rect 6050 373 6080 425
rect 6132 373 6162 425
rect 6214 373 6244 425
rect 6296 373 6822 425
rect 6874 373 6904 425
rect 6956 373 6986 425
rect 7038 373 7068 425
rect 7120 373 7936 425
rect 7988 373 8018 425
rect 8070 373 8100 425
rect 8152 373 8182 425
rect 8234 373 8760 425
rect 8812 373 8842 425
rect 8894 373 8924 425
rect 8976 373 9006 425
rect 9058 373 9584 425
rect 9636 373 9666 425
rect 9718 373 9748 425
rect 9800 373 9830 425
rect 9882 373 10408 425
rect 10460 373 10490 425
rect 10542 373 10572 425
rect 10624 373 10654 425
rect 10706 373 10707 425
rect 100 364 4023 373
tri 4023 364 4032 373 sw
tri 4176 364 4185 373 ne
rect 100 357 4032 364
tri 4032 357 4039 364 sw
rect 4185 357 10707 373
rect 100 356 4039 357
tri 4039 356 4040 357 sw
rect 4185 356 5149 357
rect 100 304 4040 356
tri 4040 304 4092 356 sw
rect 4185 304 4191 356
rect 4243 304 4259 356
rect 4311 304 4327 356
rect 4379 304 4395 356
rect 4447 304 4463 356
rect 4515 304 4531 356
rect 4583 304 4599 356
rect 4651 304 4666 356
rect 4718 304 4733 356
rect 4785 304 4800 356
rect 4852 304 4867 356
rect 4919 304 4934 356
rect 4986 304 5001 356
rect 5053 304 5068 356
rect 5120 305 5149 356
rect 5201 305 5221 357
rect 5273 305 5293 357
rect 5345 305 5365 357
rect 5417 305 5436 357
rect 5488 305 5507 357
rect 5559 305 5578 357
rect 5630 356 10707 357
rect 5630 305 5659 356
rect 5120 304 5659 305
rect 5711 304 5724 356
rect 5776 304 5789 356
rect 5841 304 5854 356
rect 5906 304 5919 356
rect 5971 304 5984 356
rect 6036 304 6049 356
rect 6101 304 6114 356
rect 6166 304 6179 356
rect 6231 304 6244 356
rect 6296 304 6309 356
rect 6361 304 6374 356
rect 6426 304 6439 356
rect 6491 304 6504 356
rect 6556 304 6569 356
rect 6621 304 6634 356
rect 6686 304 6699 356
rect 6751 304 6764 356
rect 6816 304 6829 356
rect 6881 304 6894 356
rect 6946 304 6959 356
rect 7011 304 7024 356
rect 7076 304 7089 356
rect 7141 304 7154 356
rect 7206 304 7219 356
rect 7271 304 7284 356
rect 7336 304 7349 356
rect 7401 304 7414 356
rect 7466 304 7479 356
rect 7531 304 7544 356
rect 7596 304 7609 356
rect 7661 304 7674 356
rect 7726 304 7739 356
rect 7791 304 7804 356
rect 7856 304 7869 356
rect 7921 304 7934 356
rect 7986 304 7999 356
rect 8051 304 8064 356
rect 8116 304 8129 356
rect 8181 304 8194 356
rect 8246 304 8259 356
rect 8311 304 8324 356
rect 8376 304 8389 356
rect 8441 304 8454 356
rect 8506 304 8519 356
rect 8571 304 8584 356
rect 8636 304 8649 356
rect 8701 304 8714 356
rect 8766 304 8779 356
rect 8831 304 8844 356
rect 8896 304 8909 356
rect 8961 304 8974 356
rect 9026 304 9039 356
rect 9091 304 9104 356
rect 9156 304 9169 356
rect 9221 304 9234 356
rect 9286 304 9299 356
rect 9351 304 9364 356
rect 9416 304 9429 356
rect 9481 304 9494 356
rect 9546 304 9559 356
rect 9611 304 9624 356
rect 9676 304 9689 356
rect 9741 304 9753 356
rect 9805 304 9817 356
rect 9869 304 9881 356
rect 9933 304 9945 356
rect 9997 304 10009 356
rect 10061 304 10073 356
rect 10125 304 10137 356
rect 10189 304 10201 356
rect 10253 304 10265 356
rect 10317 304 10329 356
rect 10381 304 10393 356
rect 10445 304 10457 356
rect 10509 304 10521 356
rect 10573 304 10585 356
rect 10637 304 10649 356
rect 10701 304 10707 356
rect 100 297 4092 304
tri 4092 297 4099 304 sw
rect 100 0 4099 297
rect 4185 282 10707 304
rect 4185 230 4191 282
rect 4243 230 4259 282
rect 4311 230 4327 282
rect 4379 230 4395 282
rect 4447 230 4463 282
rect 4515 230 4531 282
rect 4583 230 4599 282
rect 4651 230 4666 282
rect 4718 230 4733 282
rect 4785 230 4800 282
rect 4852 230 4867 282
rect 4919 230 4934 282
rect 4986 230 5001 282
rect 5053 230 5068 282
rect 5120 277 5659 282
rect 5120 230 5149 277
rect 4185 225 5149 230
rect 5201 225 5221 277
rect 5273 225 5293 277
rect 5345 225 5365 277
rect 5417 225 5436 277
rect 5488 225 5507 277
rect 5559 225 5578 277
rect 5630 230 5659 277
rect 5711 230 5724 282
rect 5776 230 5789 282
rect 5841 230 5854 282
rect 5906 230 5919 282
rect 5971 230 5984 282
rect 6036 230 6049 282
rect 6101 230 6114 282
rect 6166 230 6179 282
rect 6231 230 6244 282
rect 6296 230 6309 282
rect 6361 230 6374 282
rect 6426 230 6439 282
rect 6491 230 6504 282
rect 6556 230 6569 282
rect 6621 230 6634 282
rect 6686 230 6699 282
rect 6751 230 6764 282
rect 6816 230 6829 282
rect 6881 230 6894 282
rect 6946 230 6959 282
rect 7011 230 7024 282
rect 7076 230 7089 282
rect 7141 230 7154 282
rect 7206 230 7219 282
rect 7271 230 7284 282
rect 7336 230 7349 282
rect 7401 230 7414 282
rect 7466 230 7479 282
rect 7531 230 7544 282
rect 7596 230 7609 282
rect 7661 230 7674 282
rect 7726 230 7739 282
rect 7791 230 7804 282
rect 7856 230 7869 282
rect 7921 230 7934 282
rect 7986 230 7999 282
rect 8051 230 8064 282
rect 8116 230 8129 282
rect 8181 230 8194 282
rect 8246 230 8259 282
rect 8311 230 8324 282
rect 8376 230 8389 282
rect 8441 230 8454 282
rect 8506 230 8519 282
rect 8571 230 8584 282
rect 8636 230 8649 282
rect 8701 230 8714 282
rect 8766 230 8779 282
rect 8831 230 8844 282
rect 8896 230 8909 282
rect 8961 230 8974 282
rect 9026 230 9039 282
rect 9091 230 9104 282
rect 9156 230 9169 282
rect 9221 230 9234 282
rect 9286 230 9299 282
rect 9351 230 9364 282
rect 9416 230 9429 282
rect 9481 230 9494 282
rect 9546 230 9559 282
rect 9611 230 9624 282
rect 9676 230 9689 282
rect 9741 230 9753 282
rect 9805 230 9817 282
rect 9869 230 9881 282
rect 9933 230 9945 282
rect 9997 230 10009 282
rect 10061 230 10073 282
rect 10125 230 10137 282
rect 10189 230 10201 282
rect 10253 230 10265 282
rect 10317 230 10329 282
rect 10381 230 10393 282
rect 10445 230 10457 282
rect 10509 230 10521 282
rect 10573 230 10585 282
rect 10637 230 10649 282
rect 10701 230 10707 282
rect 5630 225 10707 230
rect 4185 208 10707 225
rect 4185 156 4191 208
rect 4243 156 4259 208
rect 4311 156 4327 208
rect 4379 156 4395 208
rect 4447 156 4463 208
rect 4515 156 4531 208
rect 4583 156 4599 208
rect 4651 156 4666 208
rect 4718 156 4733 208
rect 4785 156 4800 208
rect 4852 156 4867 208
rect 4919 156 4934 208
rect 4986 156 5001 208
rect 5053 156 5068 208
rect 5120 197 5659 208
rect 5120 156 5149 197
rect 4185 145 5149 156
rect 5201 145 5221 197
rect 5273 145 5293 197
rect 5345 145 5365 197
rect 5417 145 5436 197
rect 5488 145 5507 197
rect 5559 145 5578 197
rect 5630 156 5659 197
rect 5711 156 5724 208
rect 5776 156 5789 208
rect 5841 156 5854 208
rect 5906 156 5919 208
rect 5971 156 5984 208
rect 6036 156 6049 208
rect 6101 156 6114 208
rect 6166 156 6179 208
rect 6231 156 6244 208
rect 6296 156 6309 208
rect 6361 156 6374 208
rect 6426 156 6439 208
rect 6491 156 6504 208
rect 6556 156 6569 208
rect 6621 156 6634 208
rect 6686 156 6699 208
rect 6751 156 6764 208
rect 6816 156 6829 208
rect 6881 156 6894 208
rect 6946 156 6959 208
rect 7011 156 7024 208
rect 7076 156 7089 208
rect 7141 156 7154 208
rect 7206 156 7219 208
rect 7271 156 7284 208
rect 7336 156 7349 208
rect 7401 156 7414 208
rect 7466 156 7479 208
rect 7531 156 7544 208
rect 7596 156 7609 208
rect 7661 156 7674 208
rect 7726 156 7739 208
rect 7791 156 7804 208
rect 7856 156 7869 208
rect 7921 156 7934 208
rect 7986 156 7999 208
rect 8051 156 8064 208
rect 8116 156 8129 208
rect 8181 156 8194 208
rect 8246 156 8259 208
rect 8311 156 8324 208
rect 8376 156 8389 208
rect 8441 156 8454 208
rect 8506 156 8519 208
rect 8571 156 8584 208
rect 8636 156 8649 208
rect 8701 156 8714 208
rect 8766 156 8779 208
rect 8831 156 8844 208
rect 8896 156 8909 208
rect 8961 156 8974 208
rect 9026 156 9039 208
rect 9091 156 9104 208
rect 9156 156 9169 208
rect 9221 156 9234 208
rect 9286 156 9299 208
rect 9351 156 9364 208
rect 9416 156 9429 208
rect 9481 156 9494 208
rect 9546 156 9559 208
rect 9611 156 9624 208
rect 9676 156 9689 208
rect 9741 156 9753 208
rect 9805 156 9817 208
rect 9869 156 9881 208
rect 9933 156 9945 208
rect 9997 156 10009 208
rect 10061 156 10073 208
rect 10125 156 10137 208
rect 10189 156 10201 208
rect 10253 156 10265 208
rect 10317 156 10329 208
rect 10381 156 10393 208
rect 10445 156 10457 208
rect 10509 156 10521 208
rect 10573 156 10585 208
rect 10637 156 10649 208
rect 10701 156 10707 208
rect 5630 145 10707 156
rect 4185 134 10707 145
rect 4185 82 4191 134
rect 4243 82 4259 134
rect 4311 82 4327 134
rect 4379 82 4395 134
rect 4447 82 4463 134
rect 4515 82 4531 134
rect 4583 82 4599 134
rect 4651 82 4666 134
rect 4718 82 4733 134
rect 4785 82 4800 134
rect 4852 82 4867 134
rect 4919 82 4934 134
rect 4986 82 5001 134
rect 5053 82 5068 134
rect 5120 117 5659 134
rect 5120 82 5149 117
rect 4185 65 5149 82
rect 5201 65 5221 117
rect 5273 65 5293 117
rect 5345 65 5365 117
rect 5417 65 5436 117
rect 5488 65 5507 117
rect 5559 65 5578 117
rect 5630 82 5659 117
rect 5711 82 5724 134
rect 5776 82 5789 134
rect 5841 82 5854 134
rect 5906 82 5919 134
rect 5971 82 5984 134
rect 6036 82 6049 134
rect 6101 82 6114 134
rect 6166 82 6179 134
rect 6231 82 6244 134
rect 6296 82 6309 134
rect 6361 82 6374 134
rect 6426 82 6439 134
rect 6491 82 6504 134
rect 6556 82 6569 134
rect 6621 82 6634 134
rect 6686 82 6699 134
rect 6751 82 6764 134
rect 6816 82 6829 134
rect 6881 82 6894 134
rect 6946 82 6959 134
rect 7011 82 7024 134
rect 7076 82 7089 134
rect 7141 82 7154 134
rect 7206 82 7219 134
rect 7271 82 7284 134
rect 7336 82 7349 134
rect 7401 82 7414 134
rect 7466 82 7479 134
rect 7531 82 7544 134
rect 7596 82 7609 134
rect 7661 82 7674 134
rect 7726 82 7739 134
rect 7791 82 7804 134
rect 7856 82 7869 134
rect 7921 82 7934 134
rect 7986 82 7999 134
rect 8051 82 8064 134
rect 8116 82 8129 134
rect 8181 82 8194 134
rect 8246 82 8259 134
rect 8311 82 8324 134
rect 8376 82 8389 134
rect 8441 82 8454 134
rect 8506 82 8519 134
rect 8571 82 8584 134
rect 8636 82 8649 134
rect 8701 82 8714 134
rect 8766 82 8779 134
rect 8831 82 8844 134
rect 8896 82 8909 134
rect 8961 82 8974 134
rect 9026 82 9039 134
rect 9091 82 9104 134
rect 9156 82 9169 134
rect 9221 82 9234 134
rect 9286 82 9299 134
rect 9351 82 9364 134
rect 9416 82 9429 134
rect 9481 82 9494 134
rect 9546 82 9559 134
rect 9611 82 9624 134
rect 9676 82 9689 134
rect 9741 82 9753 134
rect 9805 82 9817 134
rect 9869 82 9881 134
rect 9933 82 9945 134
rect 9997 82 10009 134
rect 10061 82 10073 134
rect 10125 82 10137 134
rect 10189 82 10201 134
rect 10253 82 10265 134
rect 10317 82 10329 134
rect 10381 82 10393 134
rect 10445 82 10457 134
rect 10509 82 10521 134
rect 10573 82 10585 134
rect 10637 82 10649 134
rect 10701 82 10707 134
rect 5630 65 10707 82
rect 4185 60 10707 65
rect 4185 8 4191 60
rect 4243 8 4259 60
rect 4311 8 4327 60
rect 4379 8 4395 60
rect 4447 8 4463 60
rect 4515 8 4531 60
rect 4583 8 4599 60
rect 4651 8 4666 60
rect 4718 8 4733 60
rect 4785 8 4800 60
rect 4852 8 4867 60
rect 4919 8 4934 60
rect 4986 8 5001 60
rect 5053 8 5068 60
rect 5120 8 5659 60
rect 5711 8 5724 60
rect 5776 8 5789 60
rect 5841 8 5854 60
rect 5906 8 5919 60
rect 5971 8 5984 60
rect 6036 8 6049 60
rect 6101 8 6114 60
rect 6166 8 6179 60
rect 6231 8 6244 60
rect 6296 8 6309 60
rect 6361 8 6374 60
rect 6426 8 6439 60
rect 6491 8 6504 60
rect 6556 8 6569 60
rect 6621 8 6634 60
rect 6686 8 6699 60
rect 6751 8 6764 60
rect 6816 8 6829 60
rect 6881 8 6894 60
rect 6946 8 6959 60
rect 7011 8 7024 60
rect 7076 8 7089 60
rect 7141 8 7154 60
rect 7206 8 7219 60
rect 7271 8 7284 60
rect 7336 8 7349 60
rect 7401 8 7414 60
rect 7466 8 7479 60
rect 7531 8 7544 60
rect 7596 8 7609 60
rect 7661 8 7674 60
rect 7726 8 7739 60
rect 7791 8 7804 60
rect 7856 8 7869 60
rect 7921 8 7934 60
rect 7986 8 7999 60
rect 8051 8 8064 60
rect 8116 8 8129 60
rect 8181 8 8194 60
rect 8246 8 8259 60
rect 8311 8 8324 60
rect 8376 8 8389 60
rect 8441 8 8454 60
rect 8506 8 8519 60
rect 8571 8 8584 60
rect 8636 8 8649 60
rect 8701 8 8714 60
rect 8766 8 8779 60
rect 8831 8 8844 60
rect 8896 8 8909 60
rect 8961 8 8974 60
rect 9026 8 9039 60
rect 9091 8 9104 60
rect 9156 8 9169 60
rect 9221 8 9234 60
rect 9286 8 9299 60
rect 9351 8 9364 60
rect 9416 8 9429 60
rect 9481 8 9494 60
rect 9546 8 9559 60
rect 9611 8 9624 60
rect 9676 8 9689 60
rect 9741 8 9753 60
rect 9805 8 9817 60
rect 9869 8 9881 60
rect 9933 8 9945 60
rect 9997 8 10009 60
rect 10061 8 10073 60
rect 10125 8 10137 60
rect 10189 8 10201 60
rect 10253 8 10265 60
rect 10317 8 10329 60
rect 10381 8 10393 60
rect 10445 8 10457 60
rect 10509 8 10521 60
rect 10573 8 10585 60
rect 10637 8 10649 60
rect 10701 8 10707 60
rect 4185 0 10707 8
tri 10819 1563 11164 1908 se
rect 11164 1563 14940 1908
rect 10819 0 14940 1563
<< via2 >>
rect 3513 37840 3556 37892
rect 3556 37840 3569 37892
rect 3594 37840 3622 37892
rect 3622 37840 3650 37892
rect 3513 37836 3569 37840
rect 3594 37836 3650 37840
rect 3675 37836 3731 37892
rect 3756 37836 3812 37892
rect 3837 37836 3893 37892
rect 3918 37840 4058 37892
rect 4058 37840 4110 37892
rect 4110 37840 4124 37892
rect 4124 37840 4176 37892
rect 4176 37840 4612 37892
rect 4612 37840 4664 37892
rect 4664 37840 4678 37892
rect 4678 37840 4730 37892
rect 4730 37840 5014 37892
rect 5216 37840 5218 37892
rect 5218 37840 5232 37892
rect 5232 37840 5272 37892
rect 3918 37825 5014 37840
rect 5216 37836 5272 37840
rect 5297 37836 5353 37892
rect 5378 37836 5434 37892
rect 5459 37836 5515 37892
rect 5540 37836 5596 37892
rect 5621 37836 5677 37892
rect 5702 37840 5720 37892
rect 5720 37840 5758 37892
rect 5783 37840 5786 37892
rect 5786 37840 5838 37892
rect 5838 37840 5839 37892
rect 5702 37836 5758 37840
rect 5783 37836 5839 37840
rect 5864 37836 5920 37892
rect 5945 37836 6001 37892
rect 6026 37836 6082 37892
rect 6107 37836 6163 37892
rect 6188 37836 6244 37892
rect 6269 37840 6274 37892
rect 6274 37840 6325 37892
rect 6350 37840 6392 37892
rect 6392 37840 6406 37892
rect 6269 37836 6325 37840
rect 6350 37836 6406 37840
rect 6431 37836 6487 37892
rect 6512 37836 6568 37892
rect 6593 37836 6649 37892
rect 6674 37836 6730 37892
rect 6755 37836 6811 37892
rect 6836 37840 6880 37892
rect 6880 37840 6892 37892
rect 6917 37840 6946 37892
rect 6946 37840 6973 37892
rect 6836 37836 6892 37840
rect 6917 37836 6973 37840
rect 6998 37836 7054 37892
rect 7079 37836 7135 37892
rect 3513 37773 3556 37812
rect 3556 37773 3569 37812
rect 3594 37773 3622 37812
rect 3622 37773 3650 37812
rect 3513 37758 3569 37773
rect 3594 37758 3650 37773
rect 3513 37756 3556 37758
rect 3556 37756 3569 37758
rect 3594 37756 3622 37758
rect 3622 37756 3650 37758
rect 3675 37756 3731 37812
rect 3756 37756 3812 37812
rect 3837 37756 3893 37812
rect 3918 37773 4058 37825
rect 4058 37773 4110 37825
rect 4110 37773 4124 37825
rect 4124 37773 4176 37825
rect 4176 37773 4612 37825
rect 4612 37773 4664 37825
rect 4664 37773 4678 37825
rect 4678 37773 4730 37825
rect 4730 37773 5014 37825
rect 5216 37773 5218 37812
rect 5218 37773 5232 37812
rect 5232 37773 5272 37812
rect 3918 37758 5014 37773
rect 5216 37758 5272 37773
rect 3513 37706 3556 37732
rect 3556 37706 3569 37732
rect 3594 37706 3622 37732
rect 3622 37706 3650 37732
rect 3513 37691 3569 37706
rect 3594 37691 3650 37706
rect 3513 37676 3556 37691
rect 3556 37676 3569 37691
rect 3594 37676 3622 37691
rect 3622 37676 3650 37691
rect 3675 37676 3731 37732
rect 3756 37676 3812 37732
rect 3837 37676 3893 37732
rect 3918 37706 4058 37758
rect 4058 37706 4110 37758
rect 4110 37706 4124 37758
rect 4124 37706 4176 37758
rect 4176 37706 4612 37758
rect 4612 37706 4664 37758
rect 4664 37706 4678 37758
rect 4678 37706 4730 37758
rect 4730 37706 5014 37758
rect 5216 37756 5218 37758
rect 5218 37756 5232 37758
rect 5232 37756 5272 37758
rect 5297 37756 5353 37812
rect 5378 37756 5434 37812
rect 5459 37756 5515 37812
rect 5540 37756 5596 37812
rect 5621 37756 5677 37812
rect 5702 37773 5720 37812
rect 5720 37773 5758 37812
rect 5783 37773 5786 37812
rect 5786 37773 5838 37812
rect 5838 37773 5839 37812
rect 5702 37758 5758 37773
rect 5783 37758 5839 37773
rect 5702 37756 5720 37758
rect 5720 37756 5758 37758
rect 5783 37756 5786 37758
rect 5786 37756 5838 37758
rect 5838 37756 5839 37758
rect 5864 37756 5920 37812
rect 5945 37756 6001 37812
rect 6026 37756 6082 37812
rect 6107 37756 6163 37812
rect 6188 37756 6244 37812
rect 6269 37773 6274 37812
rect 6274 37773 6325 37812
rect 6350 37773 6392 37812
rect 6392 37773 6406 37812
rect 6269 37758 6325 37773
rect 6350 37758 6406 37773
rect 6269 37756 6274 37758
rect 6274 37756 6325 37758
rect 5216 37706 5218 37732
rect 5218 37706 5232 37732
rect 5232 37706 5272 37732
rect 3918 37691 5014 37706
rect 5216 37691 5272 37706
rect 3513 37639 3556 37652
rect 3556 37639 3569 37652
rect 3594 37639 3622 37652
rect 3622 37639 3650 37652
rect 3513 37624 3569 37639
rect 3594 37624 3650 37639
rect 3513 37596 3556 37624
rect 3556 37596 3569 37624
rect 3594 37596 3622 37624
rect 3622 37596 3650 37624
rect 3675 37596 3731 37652
rect 3756 37596 3812 37652
rect 3837 37596 3893 37652
rect 3918 37639 4058 37691
rect 4058 37639 4110 37691
rect 4110 37639 4124 37691
rect 4124 37639 4176 37691
rect 4176 37639 4612 37691
rect 4612 37639 4664 37691
rect 4664 37639 4678 37691
rect 4678 37639 4730 37691
rect 4730 37639 5014 37691
rect 5216 37676 5218 37691
rect 5218 37676 5232 37691
rect 5232 37676 5272 37691
rect 5297 37676 5353 37732
rect 5378 37676 5434 37732
rect 5459 37676 5515 37732
rect 5540 37676 5596 37732
rect 5621 37676 5677 37732
rect 5702 37706 5720 37732
rect 5720 37706 5758 37732
rect 5783 37706 5786 37732
rect 5786 37706 5838 37732
rect 5838 37706 5839 37732
rect 5702 37691 5758 37706
rect 5783 37691 5839 37706
rect 5702 37676 5720 37691
rect 5720 37676 5758 37691
rect 5783 37676 5786 37691
rect 5786 37676 5838 37691
rect 5838 37676 5839 37691
rect 5864 37676 5920 37732
rect 5945 37676 6001 37732
rect 6026 37676 6082 37732
rect 6107 37676 6163 37732
rect 6188 37676 6244 37732
rect 6269 37706 6274 37732
rect 6274 37706 6325 37732
rect 6350 37756 6392 37758
rect 6392 37756 6406 37758
rect 6431 37756 6487 37812
rect 6512 37756 6568 37812
rect 6593 37756 6649 37812
rect 6674 37756 6730 37812
rect 6755 37756 6811 37812
rect 6836 37773 6880 37812
rect 6880 37773 6892 37812
rect 6917 37773 6946 37812
rect 6946 37773 6973 37812
rect 6836 37758 6892 37773
rect 6917 37758 6973 37773
rect 6836 37756 6880 37758
rect 6880 37756 6892 37758
rect 6917 37756 6946 37758
rect 6946 37756 6973 37758
rect 6998 37756 7054 37812
rect 7079 37756 7135 37812
rect 6350 37706 6392 37732
rect 6392 37706 6406 37732
rect 6269 37691 6325 37706
rect 6350 37691 6406 37706
rect 6269 37676 6274 37691
rect 6274 37676 6325 37691
rect 5216 37639 5218 37652
rect 5218 37639 5232 37652
rect 5232 37639 5272 37652
rect 3918 37624 5014 37639
rect 5216 37624 5272 37639
rect 3918 37572 4058 37624
rect 4058 37572 4110 37624
rect 4110 37572 4124 37624
rect 4124 37572 4176 37624
rect 4176 37572 4612 37624
rect 4612 37572 4664 37624
rect 4664 37572 4678 37624
rect 4678 37572 4730 37624
rect 4730 37572 5014 37624
rect 5216 37596 5218 37624
rect 5218 37596 5232 37624
rect 5232 37596 5272 37624
rect 5297 37596 5353 37652
rect 5378 37596 5434 37652
rect 5459 37596 5515 37652
rect 5540 37596 5596 37652
rect 5621 37596 5677 37652
rect 5702 37639 5720 37652
rect 5720 37639 5758 37652
rect 5783 37639 5786 37652
rect 5786 37639 5838 37652
rect 5838 37639 5839 37652
rect 5702 37624 5758 37639
rect 5783 37624 5839 37639
rect 5702 37596 5720 37624
rect 5720 37596 5758 37624
rect 5783 37596 5786 37624
rect 5786 37596 5838 37624
rect 5838 37596 5839 37624
rect 5864 37596 5920 37652
rect 5945 37596 6001 37652
rect 6026 37596 6082 37652
rect 6107 37596 6163 37652
rect 6188 37596 6244 37652
rect 6269 37639 6274 37652
rect 6274 37639 6325 37652
rect 6350 37676 6392 37691
rect 6392 37676 6406 37691
rect 6431 37676 6487 37732
rect 6512 37676 6568 37732
rect 6593 37676 6649 37732
rect 6674 37676 6730 37732
rect 6755 37676 6811 37732
rect 6836 37706 6880 37732
rect 6880 37706 6892 37732
rect 6917 37706 6946 37732
rect 6946 37706 6973 37732
rect 6836 37691 6892 37706
rect 6917 37691 6973 37706
rect 6836 37676 6880 37691
rect 6880 37676 6892 37691
rect 6917 37676 6946 37691
rect 6946 37676 6973 37691
rect 6998 37676 7054 37732
rect 7079 37676 7135 37732
rect 6350 37639 6392 37652
rect 6392 37639 6406 37652
rect 6269 37624 6325 37639
rect 6350 37624 6406 37639
rect 6269 37596 6274 37624
rect 6274 37596 6325 37624
rect 6350 37596 6392 37624
rect 6392 37596 6406 37624
rect 6431 37596 6487 37652
rect 6512 37596 6568 37652
rect 6593 37596 6649 37652
rect 6674 37596 6730 37652
rect 6755 37596 6811 37652
rect 6836 37639 6880 37652
rect 6880 37639 6892 37652
rect 6917 37639 6946 37652
rect 6946 37639 6973 37652
rect 6836 37624 6892 37639
rect 6917 37624 6973 37639
rect 6836 37596 6880 37624
rect 6880 37596 6892 37624
rect 6917 37596 6946 37624
rect 6946 37596 6973 37624
rect 6998 37596 7054 37652
rect 7079 37596 7135 37652
rect 3513 37557 3569 37572
rect 3594 37557 3650 37572
rect 3513 37516 3556 37557
rect 3556 37516 3569 37557
rect 3594 37516 3622 37557
rect 3622 37516 3650 37557
rect 3675 37516 3731 37572
rect 3756 37516 3812 37572
rect 3837 37516 3893 37572
rect 3918 37557 5014 37572
rect 5216 37557 5272 37572
rect 3918 37505 4058 37557
rect 4058 37505 4110 37557
rect 4110 37505 4124 37557
rect 4124 37505 4176 37557
rect 4176 37505 4612 37557
rect 4612 37505 4664 37557
rect 4664 37505 4678 37557
rect 4678 37505 4730 37557
rect 4730 37505 5014 37557
rect 5216 37516 5218 37557
rect 5218 37516 5232 37557
rect 5232 37516 5272 37557
rect 5297 37516 5353 37572
rect 5378 37516 5434 37572
rect 5459 37516 5515 37572
rect 5540 37516 5596 37572
rect 5621 37516 5677 37572
rect 5702 37557 5758 37572
rect 5783 37557 5839 37572
rect 5702 37516 5720 37557
rect 5720 37516 5758 37557
rect 5783 37516 5786 37557
rect 5786 37516 5838 37557
rect 5838 37516 5839 37557
rect 5864 37516 5920 37572
rect 5945 37516 6001 37572
rect 6026 37516 6082 37572
rect 6107 37516 6163 37572
rect 6188 37516 6244 37572
rect 6269 37557 6325 37572
rect 6350 37557 6406 37572
rect 6269 37516 6274 37557
rect 6274 37516 6325 37557
rect 6350 37516 6392 37557
rect 6392 37516 6406 37557
rect 6431 37516 6487 37572
rect 6512 37516 6568 37572
rect 6593 37516 6649 37572
rect 6674 37516 6730 37572
rect 6755 37516 6811 37572
rect 6836 37557 6892 37572
rect 6917 37557 6973 37572
rect 6836 37516 6880 37557
rect 6880 37516 6892 37557
rect 6917 37516 6946 37557
rect 6946 37516 6973 37557
rect 6998 37516 7054 37572
rect 7079 37516 7135 37572
rect 3513 37490 3569 37492
rect 3594 37490 3650 37492
rect 3513 37438 3556 37490
rect 3556 37438 3569 37490
rect 3594 37438 3622 37490
rect 3622 37438 3650 37490
rect 3513 37436 3569 37438
rect 3594 37436 3650 37438
rect 3675 37436 3731 37492
rect 3756 37436 3812 37492
rect 3837 37436 3893 37492
rect 3918 37490 5014 37505
rect 5216 37490 5272 37492
rect 3918 37438 4058 37490
rect 4058 37438 4110 37490
rect 4110 37438 4124 37490
rect 4124 37438 4176 37490
rect 4176 37438 4612 37490
rect 4612 37438 4664 37490
rect 4664 37438 4678 37490
rect 4678 37438 4730 37490
rect 4730 37438 5014 37490
rect 5216 37438 5218 37490
rect 5218 37438 5232 37490
rect 5232 37438 5272 37490
rect 3918 37423 5014 37438
rect 5216 37436 5272 37438
rect 5297 37436 5353 37492
rect 5378 37436 5434 37492
rect 5459 37436 5515 37492
rect 5540 37436 5596 37492
rect 5621 37436 5677 37492
rect 5702 37490 5758 37492
rect 5783 37490 5839 37492
rect 5702 37438 5720 37490
rect 5720 37438 5758 37490
rect 5783 37438 5786 37490
rect 5786 37438 5838 37490
rect 5838 37438 5839 37490
rect 5702 37436 5758 37438
rect 5783 37436 5839 37438
rect 5864 37436 5920 37492
rect 5945 37436 6001 37492
rect 6026 37436 6082 37492
rect 6107 37436 6163 37492
rect 6188 37436 6244 37492
rect 6269 37490 6325 37492
rect 6350 37490 6406 37492
rect 6269 37438 6274 37490
rect 6274 37438 6325 37490
rect 6350 37438 6392 37490
rect 6392 37438 6406 37490
rect 6269 37436 6325 37438
rect 6350 37436 6406 37438
rect 6431 37436 6487 37492
rect 6512 37436 6568 37492
rect 6593 37436 6649 37492
rect 6674 37436 6730 37492
rect 6755 37436 6811 37492
rect 6836 37490 6892 37492
rect 6917 37490 6973 37492
rect 6836 37438 6880 37490
rect 6880 37438 6892 37490
rect 6917 37438 6946 37490
rect 6946 37438 6973 37490
rect 6836 37436 6892 37438
rect 6917 37436 6973 37438
rect 6998 37436 7054 37492
rect 7079 37436 7135 37492
rect 3513 37371 3556 37412
rect 3556 37371 3569 37412
rect 3594 37371 3622 37412
rect 3622 37371 3650 37412
rect 3513 37356 3569 37371
rect 3594 37356 3650 37371
rect 3675 37356 3731 37412
rect 3756 37356 3812 37412
rect 3837 37356 3893 37412
rect 3918 37371 4058 37423
rect 4058 37371 4110 37423
rect 4110 37371 4124 37423
rect 4124 37371 4176 37423
rect 4176 37371 4612 37423
rect 4612 37371 4664 37423
rect 4664 37371 4678 37423
rect 4678 37371 4730 37423
rect 4730 37371 5014 37423
rect 5216 37371 5218 37412
rect 5218 37371 5232 37412
rect 5232 37371 5272 37412
rect 3918 37356 5014 37371
rect 5216 37356 5272 37371
rect 5297 37356 5353 37412
rect 5378 37356 5434 37412
rect 5459 37356 5515 37412
rect 5540 37356 5596 37412
rect 5621 37356 5677 37412
rect 5702 37371 5720 37412
rect 5720 37371 5758 37412
rect 5783 37371 5786 37412
rect 5786 37371 5838 37412
rect 5838 37371 5839 37412
rect 5702 37356 5758 37371
rect 5783 37356 5839 37371
rect 5864 37356 5920 37412
rect 5945 37356 6001 37412
rect 6026 37356 6082 37412
rect 6107 37356 6163 37412
rect 6188 37356 6244 37412
rect 6269 37371 6274 37412
rect 6274 37371 6325 37412
rect 6350 37371 6392 37412
rect 6392 37371 6406 37412
rect 6269 37356 6325 37371
rect 6350 37356 6406 37371
rect 6431 37356 6487 37412
rect 6512 37356 6568 37412
rect 6593 37356 6649 37412
rect 6674 37356 6730 37412
rect 6755 37356 6811 37412
rect 6836 37371 6880 37412
rect 6880 37371 6892 37412
rect 6917 37371 6946 37412
rect 6946 37371 6973 37412
rect 6836 37356 6892 37371
rect 6917 37356 6973 37371
rect 6998 37356 7054 37412
rect 7079 37356 7135 37412
rect 3513 37304 3556 37332
rect 3556 37304 3569 37332
rect 3594 37304 3622 37332
rect 3622 37304 3650 37332
rect 3513 37289 3569 37304
rect 3594 37289 3650 37304
rect 3513 37276 3556 37289
rect 3556 37276 3569 37289
rect 3594 37276 3622 37289
rect 3622 37276 3650 37289
rect 3675 37276 3731 37332
rect 3756 37276 3812 37332
rect 3837 37276 3893 37332
rect 3918 37304 4058 37356
rect 4058 37304 4110 37356
rect 4110 37304 4124 37356
rect 4124 37304 4176 37356
rect 4176 37304 4612 37356
rect 4612 37304 4664 37356
rect 4664 37304 4678 37356
rect 4678 37304 4730 37356
rect 4730 37304 5014 37356
rect 5216 37304 5218 37332
rect 5218 37304 5232 37332
rect 5232 37304 5272 37332
rect 3918 37289 5014 37304
rect 5216 37289 5272 37304
rect 3513 37237 3556 37252
rect 3556 37237 3569 37252
rect 3594 37237 3622 37252
rect 3622 37237 3650 37252
rect 3513 37222 3569 37237
rect 3594 37222 3650 37237
rect 3513 37196 3556 37222
rect 3556 37196 3569 37222
rect 3594 37196 3622 37222
rect 3622 37196 3650 37222
rect 3675 37196 3731 37252
rect 3756 37196 3812 37252
rect 3837 37196 3893 37252
rect 3918 37237 4058 37289
rect 4058 37237 4110 37289
rect 4110 37237 4124 37289
rect 4124 37237 4176 37289
rect 4176 37237 4612 37289
rect 4612 37237 4664 37289
rect 4664 37237 4678 37289
rect 4678 37237 4730 37289
rect 4730 37237 5014 37289
rect 5216 37276 5218 37289
rect 5218 37276 5232 37289
rect 5232 37276 5272 37289
rect 5297 37276 5353 37332
rect 5378 37276 5434 37332
rect 5459 37276 5515 37332
rect 5540 37276 5596 37332
rect 5621 37276 5677 37332
rect 5702 37304 5720 37332
rect 5720 37304 5758 37332
rect 5783 37304 5786 37332
rect 5786 37304 5838 37332
rect 5838 37304 5839 37332
rect 5702 37289 5758 37304
rect 5783 37289 5839 37304
rect 5702 37276 5720 37289
rect 5720 37276 5758 37289
rect 5783 37276 5786 37289
rect 5786 37276 5838 37289
rect 5838 37276 5839 37289
rect 5864 37276 5920 37332
rect 5945 37276 6001 37332
rect 6026 37276 6082 37332
rect 6107 37276 6163 37332
rect 6188 37276 6244 37332
rect 6269 37304 6274 37332
rect 6274 37304 6325 37332
rect 6350 37304 6392 37332
rect 6392 37304 6406 37332
rect 6269 37289 6325 37304
rect 6350 37289 6406 37304
rect 6269 37276 6274 37289
rect 6274 37276 6325 37289
rect 5216 37237 5218 37252
rect 5218 37237 5232 37252
rect 5232 37237 5272 37252
rect 3918 37222 5014 37237
rect 5216 37222 5272 37237
rect 3513 37170 3556 37172
rect 3556 37170 3569 37172
rect 3594 37170 3622 37172
rect 3622 37170 3650 37172
rect 3513 37155 3569 37170
rect 3594 37155 3650 37170
rect 3513 37116 3556 37155
rect 3556 37116 3569 37155
rect 3594 37116 3622 37155
rect 3622 37116 3650 37155
rect 3675 37116 3731 37172
rect 3756 37116 3812 37172
rect 3837 37116 3893 37172
rect 3918 37170 4058 37222
rect 4058 37170 4110 37222
rect 4110 37170 4124 37222
rect 4124 37170 4176 37222
rect 4176 37170 4612 37222
rect 4612 37170 4664 37222
rect 4664 37170 4678 37222
rect 4678 37170 4730 37222
rect 4730 37170 5014 37222
rect 5216 37196 5218 37222
rect 5218 37196 5232 37222
rect 5232 37196 5272 37222
rect 5297 37196 5353 37252
rect 5378 37196 5434 37252
rect 5459 37196 5515 37252
rect 5540 37196 5596 37252
rect 5621 37196 5677 37252
rect 5702 37237 5720 37252
rect 5720 37237 5758 37252
rect 5783 37237 5786 37252
rect 5786 37237 5838 37252
rect 5838 37237 5839 37252
rect 5702 37222 5758 37237
rect 5783 37222 5839 37237
rect 5702 37196 5720 37222
rect 5720 37196 5758 37222
rect 5783 37196 5786 37222
rect 5786 37196 5838 37222
rect 5838 37196 5839 37222
rect 5864 37196 5920 37252
rect 5945 37196 6001 37252
rect 6026 37196 6082 37252
rect 6107 37196 6163 37252
rect 6188 37196 6244 37252
rect 6269 37237 6274 37252
rect 6274 37237 6325 37252
rect 6350 37276 6392 37289
rect 6392 37276 6406 37289
rect 6431 37276 6487 37332
rect 6512 37276 6568 37332
rect 6593 37276 6649 37332
rect 6674 37276 6730 37332
rect 6755 37276 6811 37332
rect 6836 37304 6880 37332
rect 6880 37304 6892 37332
rect 6917 37304 6946 37332
rect 6946 37304 6973 37332
rect 6836 37289 6892 37304
rect 6917 37289 6973 37304
rect 6836 37276 6880 37289
rect 6880 37276 6892 37289
rect 6917 37276 6946 37289
rect 6946 37276 6973 37289
rect 6998 37276 7054 37332
rect 7079 37276 7135 37332
rect 6350 37237 6392 37252
rect 6392 37237 6406 37252
rect 6269 37222 6325 37237
rect 6350 37222 6406 37237
rect 6269 37196 6274 37222
rect 6274 37196 6325 37222
rect 5216 37170 5218 37172
rect 5218 37170 5232 37172
rect 5232 37170 5272 37172
rect 3918 37155 5014 37170
rect 5216 37155 5272 37170
rect 3918 37103 4058 37155
rect 4058 37103 4110 37155
rect 4110 37103 4124 37155
rect 4124 37103 4176 37155
rect 4176 37103 4612 37155
rect 4612 37103 4664 37155
rect 4664 37103 4678 37155
rect 4678 37103 4730 37155
rect 4730 37103 5014 37155
rect 5216 37116 5218 37155
rect 5218 37116 5232 37155
rect 5232 37116 5272 37155
rect 5297 37116 5353 37172
rect 5378 37116 5434 37172
rect 5459 37116 5515 37172
rect 5540 37116 5596 37172
rect 5621 37116 5677 37172
rect 5702 37170 5720 37172
rect 5720 37170 5758 37172
rect 5783 37170 5786 37172
rect 5786 37170 5838 37172
rect 5838 37170 5839 37172
rect 5702 37155 5758 37170
rect 5783 37155 5839 37170
rect 5702 37116 5720 37155
rect 5720 37116 5758 37155
rect 5783 37116 5786 37155
rect 5786 37116 5838 37155
rect 5838 37116 5839 37155
rect 5864 37116 5920 37172
rect 5945 37116 6001 37172
rect 6026 37116 6082 37172
rect 6107 37116 6163 37172
rect 6188 37116 6244 37172
rect 6269 37170 6274 37172
rect 6274 37170 6325 37172
rect 6350 37196 6392 37222
rect 6392 37196 6406 37222
rect 6431 37196 6487 37252
rect 6512 37196 6568 37252
rect 6593 37196 6649 37252
rect 6674 37196 6730 37252
rect 6755 37196 6811 37252
rect 6836 37237 6880 37252
rect 6880 37237 6892 37252
rect 6917 37237 6946 37252
rect 6946 37237 6973 37252
rect 6836 37222 6892 37237
rect 6917 37222 6973 37237
rect 6836 37196 6880 37222
rect 6880 37196 6892 37222
rect 6917 37196 6946 37222
rect 6946 37196 6973 37222
rect 6998 37196 7054 37252
rect 7079 37196 7135 37252
rect 6350 37170 6392 37172
rect 6392 37170 6406 37172
rect 6269 37155 6325 37170
rect 6350 37155 6406 37170
rect 6269 37116 6274 37155
rect 6274 37116 6325 37155
rect 6350 37116 6392 37155
rect 6392 37116 6406 37155
rect 6431 37116 6487 37172
rect 6512 37116 6568 37172
rect 6593 37116 6649 37172
rect 6674 37116 6730 37172
rect 6755 37116 6811 37172
rect 6836 37170 6880 37172
rect 6880 37170 6892 37172
rect 6917 37170 6946 37172
rect 6946 37170 6973 37172
rect 6836 37155 6892 37170
rect 6917 37155 6973 37170
rect 6836 37116 6880 37155
rect 6880 37116 6892 37155
rect 6917 37116 6946 37155
rect 6946 37116 6973 37155
rect 6998 37116 7054 37172
rect 7079 37116 7135 37172
rect 3513 37088 3569 37092
rect 3594 37088 3650 37092
rect 3513 37036 3556 37088
rect 3556 37036 3569 37088
rect 3594 37036 3622 37088
rect 3622 37036 3650 37088
rect 3675 37036 3731 37092
rect 3756 37036 3812 37092
rect 3837 37036 3893 37092
rect 3918 37088 5014 37103
rect 5216 37088 5272 37092
rect 3918 37036 4058 37088
rect 4058 37036 4110 37088
rect 4110 37036 4124 37088
rect 4124 37036 4176 37088
rect 4176 37036 4612 37088
rect 4612 37036 4664 37088
rect 4664 37036 4678 37088
rect 4678 37036 4730 37088
rect 4730 37036 5014 37088
rect 5216 37036 5218 37088
rect 5218 37036 5232 37088
rect 5232 37036 5272 37088
rect 5297 37036 5353 37092
rect 5378 37036 5434 37092
rect 5459 37036 5515 37092
rect 5540 37036 5596 37092
rect 5621 37036 5677 37092
rect 5702 37088 5758 37092
rect 5783 37088 5839 37092
rect 5702 37036 5720 37088
rect 5720 37036 5758 37088
rect 5783 37036 5786 37088
rect 5786 37036 5838 37088
rect 5838 37036 5839 37088
rect 5864 37036 5920 37092
rect 5945 37036 6001 37092
rect 6026 37036 6082 37092
rect 6107 37036 6163 37092
rect 6188 37036 6244 37092
rect 6269 37088 6325 37092
rect 6350 37088 6406 37092
rect 6269 37036 6274 37088
rect 6274 37036 6325 37088
rect 6350 37036 6392 37088
rect 6392 37036 6406 37088
rect 6431 37036 6487 37092
rect 6512 37036 6568 37092
rect 6593 37036 6649 37092
rect 6674 37036 6730 37092
rect 6755 37036 6811 37092
rect 6836 37088 6892 37092
rect 6917 37088 6973 37092
rect 6836 37036 6880 37088
rect 6880 37036 6892 37088
rect 6917 37036 6946 37088
rect 6946 37036 6973 37088
rect 6998 37036 7054 37092
rect 7079 37036 7135 37092
rect 7160 37036 7376 37892
rect 7598 37836 7654 37892
rect 7679 37836 7735 37892
rect 7760 37836 7816 37892
rect 7841 37836 7897 37892
rect 7922 37840 7936 37892
rect 7936 37840 7978 37892
rect 8003 37840 8054 37892
rect 8054 37840 8059 37892
rect 7922 37836 7978 37840
rect 8003 37836 8059 37840
rect 8084 37836 8140 37892
rect 8165 37836 8221 37892
rect 8246 37836 8302 37892
rect 8327 37836 8383 37892
rect 8408 37836 8464 37892
rect 8489 37840 8490 37892
rect 8490 37840 8542 37892
rect 8542 37840 8545 37892
rect 8570 37840 8608 37892
rect 8608 37840 8626 37892
rect 8489 37836 8545 37840
rect 8570 37836 8626 37840
rect 8651 37836 8707 37892
rect 8732 37836 8788 37892
rect 8813 37836 8869 37892
rect 8894 37836 8950 37892
rect 8975 37836 9031 37892
rect 9056 37840 9096 37892
rect 9096 37840 9110 37892
rect 9110 37840 9112 37892
rect 9137 37840 9162 37892
rect 9162 37840 9193 37892
rect 9056 37836 9112 37840
rect 9137 37836 9193 37840
rect 9218 37836 9274 37892
rect 9299 37836 9355 37892
rect 9380 37836 9436 37892
rect 9461 37836 9517 37892
rect 9542 37840 9598 37892
rect 9598 37840 9650 37892
rect 9650 37840 9664 37892
rect 9664 37840 9716 37892
rect 9716 37840 9758 37892
rect 9542 37825 9758 37840
rect 9983 37836 10039 37892
rect 10064 37836 10120 37892
rect 10145 37840 10152 37892
rect 10152 37840 10201 37892
rect 10226 37840 10270 37892
rect 10270 37840 10282 37892
rect 10145 37836 10201 37840
rect 10226 37836 10282 37840
rect 10307 37836 10363 37892
rect 10388 37836 10444 37892
rect 10469 37836 10525 37892
rect 10550 37836 10606 37892
rect 10631 37836 10687 37892
rect 10712 37840 10758 37892
rect 10758 37840 10768 37892
rect 10793 37840 10824 37892
rect 10824 37840 10849 37892
rect 10712 37836 10768 37840
rect 10793 37836 10849 37840
rect 10874 37836 10930 37892
rect 10955 37836 11011 37892
rect 11036 37836 11092 37892
rect 11117 37836 11173 37892
rect 11198 37836 11254 37892
rect 11279 37840 11312 37892
rect 11312 37840 11326 37892
rect 11326 37840 11335 37892
rect 11360 37840 11378 37892
rect 11378 37840 11416 37892
rect 11279 37836 11335 37840
rect 11360 37836 11416 37840
rect 11441 37840 11814 37892
rect 11814 37840 11866 37892
rect 11866 37840 11880 37892
rect 11880 37840 11932 37892
rect 11932 37840 12057 37892
rect 11441 37825 12057 37840
rect 7598 37756 7654 37812
rect 7679 37756 7735 37812
rect 7760 37756 7816 37812
rect 7841 37756 7897 37812
rect 7922 37773 7936 37812
rect 7936 37773 7978 37812
rect 8003 37773 8054 37812
rect 8054 37773 8059 37812
rect 7922 37758 7978 37773
rect 8003 37758 8059 37773
rect 7922 37756 7936 37758
rect 7936 37756 7978 37758
rect 7598 37676 7654 37732
rect 7679 37676 7735 37732
rect 7760 37676 7816 37732
rect 7841 37676 7897 37732
rect 7922 37706 7936 37732
rect 7936 37706 7978 37732
rect 8003 37756 8054 37758
rect 8054 37756 8059 37758
rect 8084 37756 8140 37812
rect 8165 37756 8221 37812
rect 8246 37756 8302 37812
rect 8327 37756 8383 37812
rect 8408 37756 8464 37812
rect 8489 37773 8490 37812
rect 8490 37773 8542 37812
rect 8542 37773 8545 37812
rect 8570 37773 8608 37812
rect 8608 37773 8626 37812
rect 8489 37758 8545 37773
rect 8570 37758 8626 37773
rect 8489 37756 8490 37758
rect 8490 37756 8542 37758
rect 8542 37756 8545 37758
rect 8570 37756 8608 37758
rect 8608 37756 8626 37758
rect 8651 37756 8707 37812
rect 8732 37756 8788 37812
rect 8813 37756 8869 37812
rect 8894 37756 8950 37812
rect 8975 37756 9031 37812
rect 9056 37773 9096 37812
rect 9096 37773 9110 37812
rect 9110 37773 9112 37812
rect 9137 37773 9162 37812
rect 9162 37773 9193 37812
rect 9056 37758 9112 37773
rect 9137 37758 9193 37773
rect 9056 37756 9096 37758
rect 9096 37756 9110 37758
rect 9110 37756 9112 37758
rect 9137 37756 9162 37758
rect 9162 37756 9193 37758
rect 9218 37756 9274 37812
rect 9299 37756 9355 37812
rect 9380 37756 9436 37812
rect 9461 37756 9517 37812
rect 9542 37773 9598 37825
rect 9598 37773 9650 37825
rect 9650 37773 9664 37825
rect 9664 37773 9716 37825
rect 9716 37773 9758 37825
rect 9542 37758 9758 37773
rect 8003 37706 8054 37732
rect 8054 37706 8059 37732
rect 7922 37691 7978 37706
rect 8003 37691 8059 37706
rect 7922 37676 7936 37691
rect 7936 37676 7978 37691
rect 7598 37596 7654 37652
rect 7679 37596 7735 37652
rect 7760 37596 7816 37652
rect 7841 37596 7897 37652
rect 7922 37639 7936 37652
rect 7936 37639 7978 37652
rect 8003 37676 8054 37691
rect 8054 37676 8059 37691
rect 8084 37676 8140 37732
rect 8165 37676 8221 37732
rect 8246 37676 8302 37732
rect 8327 37676 8383 37732
rect 8408 37676 8464 37732
rect 8489 37706 8490 37732
rect 8490 37706 8542 37732
rect 8542 37706 8545 37732
rect 8570 37706 8608 37732
rect 8608 37706 8626 37732
rect 8489 37691 8545 37706
rect 8570 37691 8626 37706
rect 8489 37676 8490 37691
rect 8490 37676 8542 37691
rect 8542 37676 8545 37691
rect 8570 37676 8608 37691
rect 8608 37676 8626 37691
rect 8651 37676 8707 37732
rect 8732 37676 8788 37732
rect 8813 37676 8869 37732
rect 8894 37676 8950 37732
rect 8975 37676 9031 37732
rect 9056 37706 9096 37732
rect 9096 37706 9110 37732
rect 9110 37706 9112 37732
rect 9137 37706 9162 37732
rect 9162 37706 9193 37732
rect 9056 37691 9112 37706
rect 9137 37691 9193 37706
rect 9056 37676 9096 37691
rect 9096 37676 9110 37691
rect 9110 37676 9112 37691
rect 9137 37676 9162 37691
rect 9162 37676 9193 37691
rect 9218 37676 9274 37732
rect 9299 37676 9355 37732
rect 9380 37676 9436 37732
rect 9461 37676 9517 37732
rect 9542 37706 9598 37758
rect 9598 37706 9650 37758
rect 9650 37706 9664 37758
rect 9664 37706 9716 37758
rect 9716 37706 9758 37758
rect 9983 37756 10039 37812
rect 10064 37756 10120 37812
rect 10145 37773 10152 37812
rect 10152 37773 10201 37812
rect 10226 37773 10270 37812
rect 10270 37773 10282 37812
rect 10145 37758 10201 37773
rect 10226 37758 10282 37773
rect 10145 37756 10152 37758
rect 10152 37756 10201 37758
rect 9542 37691 9758 37706
rect 8003 37639 8054 37652
rect 8054 37639 8059 37652
rect 7922 37624 7978 37639
rect 8003 37624 8059 37639
rect 7922 37596 7936 37624
rect 7936 37596 7978 37624
rect 8003 37596 8054 37624
rect 8054 37596 8059 37624
rect 8084 37596 8140 37652
rect 8165 37596 8221 37652
rect 8246 37596 8302 37652
rect 8327 37596 8383 37652
rect 8408 37596 8464 37652
rect 8489 37639 8490 37652
rect 8490 37639 8542 37652
rect 8542 37639 8545 37652
rect 8570 37639 8608 37652
rect 8608 37639 8626 37652
rect 8489 37624 8545 37639
rect 8570 37624 8626 37639
rect 8489 37596 8490 37624
rect 8490 37596 8542 37624
rect 8542 37596 8545 37624
rect 8570 37596 8608 37624
rect 8608 37596 8626 37624
rect 8651 37596 8707 37652
rect 8732 37596 8788 37652
rect 8813 37596 8869 37652
rect 8894 37596 8950 37652
rect 8975 37596 9031 37652
rect 9056 37639 9096 37652
rect 9096 37639 9110 37652
rect 9110 37639 9112 37652
rect 9137 37639 9162 37652
rect 9162 37639 9193 37652
rect 9056 37624 9112 37639
rect 9137 37624 9193 37639
rect 9056 37596 9096 37624
rect 9096 37596 9110 37624
rect 9110 37596 9112 37624
rect 9137 37596 9162 37624
rect 9162 37596 9193 37624
rect 9218 37596 9274 37652
rect 9299 37596 9355 37652
rect 9380 37596 9436 37652
rect 9461 37596 9517 37652
rect 9542 37639 9598 37691
rect 9598 37639 9650 37691
rect 9650 37639 9664 37691
rect 9664 37639 9716 37691
rect 9716 37639 9758 37691
rect 9983 37676 10039 37732
rect 10064 37676 10120 37732
rect 10145 37706 10152 37732
rect 10152 37706 10201 37732
rect 10226 37756 10270 37758
rect 10270 37756 10282 37758
rect 10307 37756 10363 37812
rect 10388 37756 10444 37812
rect 10469 37756 10525 37812
rect 10550 37756 10606 37812
rect 10631 37756 10687 37812
rect 10712 37773 10758 37812
rect 10758 37773 10768 37812
rect 10793 37773 10824 37812
rect 10824 37773 10849 37812
rect 10712 37758 10768 37773
rect 10793 37758 10849 37773
rect 10712 37756 10758 37758
rect 10758 37756 10768 37758
rect 10793 37756 10824 37758
rect 10824 37756 10849 37758
rect 10874 37756 10930 37812
rect 10955 37756 11011 37812
rect 11036 37756 11092 37812
rect 11117 37756 11173 37812
rect 11198 37756 11254 37812
rect 11279 37773 11312 37812
rect 11312 37773 11326 37812
rect 11326 37773 11335 37812
rect 11360 37773 11378 37812
rect 11378 37773 11416 37812
rect 11279 37758 11335 37773
rect 11360 37758 11416 37773
rect 11279 37756 11312 37758
rect 11312 37756 11326 37758
rect 11326 37756 11335 37758
rect 11360 37756 11378 37758
rect 11378 37756 11416 37758
rect 11441 37773 11814 37825
rect 11814 37773 11866 37825
rect 11866 37773 11880 37825
rect 11880 37773 11932 37825
rect 11932 37773 12057 37825
rect 11441 37758 12057 37773
rect 10226 37706 10270 37732
rect 10270 37706 10282 37732
rect 10145 37691 10201 37706
rect 10226 37691 10282 37706
rect 10145 37676 10152 37691
rect 10152 37676 10201 37691
rect 9542 37624 9758 37639
rect 9542 37572 9598 37624
rect 9598 37572 9650 37624
rect 9650 37572 9664 37624
rect 9664 37572 9716 37624
rect 9716 37572 9758 37624
rect 9983 37596 10039 37652
rect 10064 37596 10120 37652
rect 10145 37639 10152 37652
rect 10152 37639 10201 37652
rect 10226 37676 10270 37691
rect 10270 37676 10282 37691
rect 10307 37676 10363 37732
rect 10388 37676 10444 37732
rect 10469 37676 10525 37732
rect 10550 37676 10606 37732
rect 10631 37676 10687 37732
rect 10712 37706 10758 37732
rect 10758 37706 10768 37732
rect 10793 37706 10824 37732
rect 10824 37706 10849 37732
rect 10712 37691 10768 37706
rect 10793 37691 10849 37706
rect 10712 37676 10758 37691
rect 10758 37676 10768 37691
rect 10793 37676 10824 37691
rect 10824 37676 10849 37691
rect 10874 37676 10930 37732
rect 10955 37676 11011 37732
rect 11036 37676 11092 37732
rect 11117 37676 11173 37732
rect 11198 37676 11254 37732
rect 11279 37706 11312 37732
rect 11312 37706 11326 37732
rect 11326 37706 11335 37732
rect 11360 37706 11378 37732
rect 11378 37706 11416 37732
rect 11279 37691 11335 37706
rect 11360 37691 11416 37706
rect 11279 37676 11312 37691
rect 11312 37676 11326 37691
rect 11326 37676 11335 37691
rect 11360 37676 11378 37691
rect 11378 37676 11416 37691
rect 11441 37706 11814 37758
rect 11814 37706 11866 37758
rect 11866 37706 11880 37758
rect 11880 37706 11932 37758
rect 11932 37706 12057 37758
rect 11441 37691 12057 37706
rect 10226 37639 10270 37652
rect 10270 37639 10282 37652
rect 10145 37624 10201 37639
rect 10226 37624 10282 37639
rect 10145 37596 10152 37624
rect 10152 37596 10201 37624
rect 10226 37596 10270 37624
rect 10270 37596 10282 37624
rect 10307 37596 10363 37652
rect 10388 37596 10444 37652
rect 10469 37596 10525 37652
rect 10550 37596 10606 37652
rect 10631 37596 10687 37652
rect 10712 37639 10758 37652
rect 10758 37639 10768 37652
rect 10793 37639 10824 37652
rect 10824 37639 10849 37652
rect 10712 37624 10768 37639
rect 10793 37624 10849 37639
rect 10712 37596 10758 37624
rect 10758 37596 10768 37624
rect 10793 37596 10824 37624
rect 10824 37596 10849 37624
rect 10874 37596 10930 37652
rect 10955 37596 11011 37652
rect 11036 37596 11092 37652
rect 11117 37596 11173 37652
rect 11198 37596 11254 37652
rect 11279 37639 11312 37652
rect 11312 37639 11326 37652
rect 11326 37639 11335 37652
rect 11360 37639 11378 37652
rect 11378 37639 11416 37652
rect 11279 37624 11335 37639
rect 11360 37624 11416 37639
rect 11279 37596 11312 37624
rect 11312 37596 11326 37624
rect 11326 37596 11335 37624
rect 11360 37596 11378 37624
rect 11378 37596 11416 37624
rect 11441 37639 11814 37691
rect 11814 37639 11866 37691
rect 11866 37639 11880 37691
rect 11880 37639 11932 37691
rect 11932 37639 12057 37691
rect 11441 37624 12057 37639
rect 11441 37572 11814 37624
rect 11814 37572 11866 37624
rect 11866 37572 11880 37624
rect 11880 37572 11932 37624
rect 11932 37572 12057 37624
rect 7598 37516 7654 37572
rect 7679 37516 7735 37572
rect 7760 37516 7816 37572
rect 7841 37516 7897 37572
rect 7922 37557 7978 37572
rect 8003 37557 8059 37572
rect 7922 37516 7936 37557
rect 7936 37516 7978 37557
rect 8003 37516 8054 37557
rect 8054 37516 8059 37557
rect 8084 37516 8140 37572
rect 8165 37516 8221 37572
rect 8246 37516 8302 37572
rect 8327 37516 8383 37572
rect 8408 37516 8464 37572
rect 8489 37557 8545 37572
rect 8570 37557 8626 37572
rect 8489 37516 8490 37557
rect 8490 37516 8542 37557
rect 8542 37516 8545 37557
rect 8570 37516 8608 37557
rect 8608 37516 8626 37557
rect 8651 37516 8707 37572
rect 8732 37516 8788 37572
rect 8813 37516 8869 37572
rect 8894 37516 8950 37572
rect 8975 37516 9031 37572
rect 9056 37557 9112 37572
rect 9137 37557 9193 37572
rect 9056 37516 9096 37557
rect 9096 37516 9110 37557
rect 9110 37516 9112 37557
rect 9137 37516 9162 37557
rect 9162 37516 9193 37557
rect 9218 37516 9274 37572
rect 9299 37516 9355 37572
rect 9380 37516 9436 37572
rect 9461 37516 9517 37572
rect 9542 37557 9758 37572
rect 9542 37505 9598 37557
rect 9598 37505 9650 37557
rect 9650 37505 9664 37557
rect 9664 37505 9716 37557
rect 9716 37505 9758 37557
rect 9983 37516 10039 37572
rect 10064 37516 10120 37572
rect 10145 37557 10201 37572
rect 10226 37557 10282 37572
rect 10145 37516 10152 37557
rect 10152 37516 10201 37557
rect 10226 37516 10270 37557
rect 10270 37516 10282 37557
rect 10307 37516 10363 37572
rect 10388 37516 10444 37572
rect 10469 37516 10525 37572
rect 10550 37516 10606 37572
rect 10631 37516 10687 37572
rect 10712 37557 10768 37572
rect 10793 37557 10849 37572
rect 10712 37516 10758 37557
rect 10758 37516 10768 37557
rect 10793 37516 10824 37557
rect 10824 37516 10849 37557
rect 10874 37516 10930 37572
rect 10955 37516 11011 37572
rect 11036 37516 11092 37572
rect 11117 37516 11173 37572
rect 11198 37516 11254 37572
rect 11279 37557 11335 37572
rect 11360 37557 11416 37572
rect 11279 37516 11312 37557
rect 11312 37516 11326 37557
rect 11326 37516 11335 37557
rect 11360 37516 11378 37557
rect 11378 37516 11416 37557
rect 11441 37557 12057 37572
rect 11441 37505 11814 37557
rect 11814 37505 11866 37557
rect 11866 37505 11880 37557
rect 11880 37505 11932 37557
rect 11932 37505 12057 37557
rect 7598 37436 7654 37492
rect 7679 37436 7735 37492
rect 7760 37436 7816 37492
rect 7841 37436 7897 37492
rect 7922 37490 7978 37492
rect 8003 37490 8059 37492
rect 7922 37438 7936 37490
rect 7936 37438 7978 37490
rect 8003 37438 8054 37490
rect 8054 37438 8059 37490
rect 7922 37436 7978 37438
rect 8003 37436 8059 37438
rect 8084 37436 8140 37492
rect 8165 37436 8221 37492
rect 8246 37436 8302 37492
rect 8327 37436 8383 37492
rect 8408 37436 8464 37492
rect 8489 37490 8545 37492
rect 8570 37490 8626 37492
rect 8489 37438 8490 37490
rect 8490 37438 8542 37490
rect 8542 37438 8545 37490
rect 8570 37438 8608 37490
rect 8608 37438 8626 37490
rect 8489 37436 8545 37438
rect 8570 37436 8626 37438
rect 8651 37436 8707 37492
rect 8732 37436 8788 37492
rect 8813 37436 8869 37492
rect 8894 37436 8950 37492
rect 8975 37436 9031 37492
rect 9056 37490 9112 37492
rect 9137 37490 9193 37492
rect 9056 37438 9096 37490
rect 9096 37438 9110 37490
rect 9110 37438 9112 37490
rect 9137 37438 9162 37490
rect 9162 37438 9193 37490
rect 9056 37436 9112 37438
rect 9137 37436 9193 37438
rect 9218 37436 9274 37492
rect 9299 37436 9355 37492
rect 9380 37436 9436 37492
rect 9461 37436 9517 37492
rect 9542 37490 9758 37505
rect 9542 37438 9598 37490
rect 9598 37438 9650 37490
rect 9650 37438 9664 37490
rect 9664 37438 9716 37490
rect 9716 37438 9758 37490
rect 9542 37423 9758 37438
rect 9983 37436 10039 37492
rect 10064 37436 10120 37492
rect 10145 37490 10201 37492
rect 10226 37490 10282 37492
rect 10145 37438 10152 37490
rect 10152 37438 10201 37490
rect 10226 37438 10270 37490
rect 10270 37438 10282 37490
rect 10145 37436 10201 37438
rect 10226 37436 10282 37438
rect 10307 37436 10363 37492
rect 10388 37436 10444 37492
rect 10469 37436 10525 37492
rect 10550 37436 10606 37492
rect 10631 37436 10687 37492
rect 10712 37490 10768 37492
rect 10793 37490 10849 37492
rect 10712 37438 10758 37490
rect 10758 37438 10768 37490
rect 10793 37438 10824 37490
rect 10824 37438 10849 37490
rect 10712 37436 10768 37438
rect 10793 37436 10849 37438
rect 10874 37436 10930 37492
rect 10955 37436 11011 37492
rect 11036 37436 11092 37492
rect 11117 37436 11173 37492
rect 11198 37436 11254 37492
rect 11279 37490 11335 37492
rect 11360 37490 11416 37492
rect 11279 37438 11312 37490
rect 11312 37438 11326 37490
rect 11326 37438 11335 37490
rect 11360 37438 11378 37490
rect 11378 37438 11416 37490
rect 11279 37436 11335 37438
rect 11360 37436 11416 37438
rect 11441 37490 12057 37505
rect 11441 37438 11814 37490
rect 11814 37438 11866 37490
rect 11866 37438 11880 37490
rect 11880 37438 11932 37490
rect 11932 37438 12057 37490
rect 11441 37423 12057 37438
rect 7598 37356 7654 37412
rect 7679 37356 7735 37412
rect 7760 37356 7816 37412
rect 7841 37356 7897 37412
rect 7922 37371 7936 37412
rect 7936 37371 7978 37412
rect 8003 37371 8054 37412
rect 8054 37371 8059 37412
rect 7922 37356 7978 37371
rect 8003 37356 8059 37371
rect 8084 37356 8140 37412
rect 8165 37356 8221 37412
rect 8246 37356 8302 37412
rect 8327 37356 8383 37412
rect 8408 37356 8464 37412
rect 8489 37371 8490 37412
rect 8490 37371 8542 37412
rect 8542 37371 8545 37412
rect 8570 37371 8608 37412
rect 8608 37371 8626 37412
rect 8489 37356 8545 37371
rect 8570 37356 8626 37371
rect 8651 37356 8707 37412
rect 8732 37356 8788 37412
rect 8813 37356 8869 37412
rect 8894 37356 8950 37412
rect 8975 37356 9031 37412
rect 9056 37371 9096 37412
rect 9096 37371 9110 37412
rect 9110 37371 9112 37412
rect 9137 37371 9162 37412
rect 9162 37371 9193 37412
rect 9056 37356 9112 37371
rect 9137 37356 9193 37371
rect 9218 37356 9274 37412
rect 9299 37356 9355 37412
rect 9380 37356 9436 37412
rect 9461 37356 9517 37412
rect 9542 37371 9598 37423
rect 9598 37371 9650 37423
rect 9650 37371 9664 37423
rect 9664 37371 9716 37423
rect 9716 37371 9758 37423
rect 9542 37356 9758 37371
rect 9983 37356 10039 37412
rect 10064 37356 10120 37412
rect 10145 37371 10152 37412
rect 10152 37371 10201 37412
rect 10226 37371 10270 37412
rect 10270 37371 10282 37412
rect 10145 37356 10201 37371
rect 10226 37356 10282 37371
rect 10307 37356 10363 37412
rect 10388 37356 10444 37412
rect 10469 37356 10525 37412
rect 10550 37356 10606 37412
rect 10631 37356 10687 37412
rect 10712 37371 10758 37412
rect 10758 37371 10768 37412
rect 10793 37371 10824 37412
rect 10824 37371 10849 37412
rect 10712 37356 10768 37371
rect 10793 37356 10849 37371
rect 10874 37356 10930 37412
rect 10955 37356 11011 37412
rect 11036 37356 11092 37412
rect 11117 37356 11173 37412
rect 11198 37356 11254 37412
rect 11279 37371 11312 37412
rect 11312 37371 11326 37412
rect 11326 37371 11335 37412
rect 11360 37371 11378 37412
rect 11378 37371 11416 37412
rect 11279 37356 11335 37371
rect 11360 37356 11416 37371
rect 11441 37371 11814 37423
rect 11814 37371 11866 37423
rect 11866 37371 11880 37423
rect 11880 37371 11932 37423
rect 11932 37371 12057 37423
rect 11441 37356 12057 37371
rect 7598 37276 7654 37332
rect 7679 37276 7735 37332
rect 7760 37276 7816 37332
rect 7841 37276 7897 37332
rect 7922 37304 7936 37332
rect 7936 37304 7978 37332
rect 8003 37304 8054 37332
rect 8054 37304 8059 37332
rect 7922 37289 7978 37304
rect 8003 37289 8059 37304
rect 7922 37276 7936 37289
rect 7936 37276 7978 37289
rect 7598 37196 7654 37252
rect 7679 37196 7735 37252
rect 7760 37196 7816 37252
rect 7841 37196 7897 37252
rect 7922 37237 7936 37252
rect 7936 37237 7978 37252
rect 8003 37276 8054 37289
rect 8054 37276 8059 37289
rect 8084 37276 8140 37332
rect 8165 37276 8221 37332
rect 8246 37276 8302 37332
rect 8327 37276 8383 37332
rect 8408 37276 8464 37332
rect 8489 37304 8490 37332
rect 8490 37304 8542 37332
rect 8542 37304 8545 37332
rect 8570 37304 8608 37332
rect 8608 37304 8626 37332
rect 8489 37289 8545 37304
rect 8570 37289 8626 37304
rect 8489 37276 8490 37289
rect 8490 37276 8542 37289
rect 8542 37276 8545 37289
rect 8570 37276 8608 37289
rect 8608 37276 8626 37289
rect 8651 37276 8707 37332
rect 8732 37276 8788 37332
rect 8813 37276 8869 37332
rect 8894 37276 8950 37332
rect 8975 37276 9031 37332
rect 9056 37304 9096 37332
rect 9096 37304 9110 37332
rect 9110 37304 9112 37332
rect 9137 37304 9162 37332
rect 9162 37304 9193 37332
rect 9056 37289 9112 37304
rect 9137 37289 9193 37304
rect 9056 37276 9096 37289
rect 9096 37276 9110 37289
rect 9110 37276 9112 37289
rect 9137 37276 9162 37289
rect 9162 37276 9193 37289
rect 9218 37276 9274 37332
rect 9299 37276 9355 37332
rect 9380 37276 9436 37332
rect 9461 37276 9517 37332
rect 9542 37304 9598 37356
rect 9598 37304 9650 37356
rect 9650 37304 9664 37356
rect 9664 37304 9716 37356
rect 9716 37304 9758 37356
rect 9542 37289 9758 37304
rect 8003 37237 8054 37252
rect 8054 37237 8059 37252
rect 7922 37222 7978 37237
rect 8003 37222 8059 37237
rect 7922 37196 7936 37222
rect 7936 37196 7978 37222
rect 7598 37116 7654 37172
rect 7679 37116 7735 37172
rect 7760 37116 7816 37172
rect 7841 37116 7897 37172
rect 7922 37170 7936 37172
rect 7936 37170 7978 37172
rect 8003 37196 8054 37222
rect 8054 37196 8059 37222
rect 8084 37196 8140 37252
rect 8165 37196 8221 37252
rect 8246 37196 8302 37252
rect 8327 37196 8383 37252
rect 8408 37196 8464 37252
rect 8489 37237 8490 37252
rect 8490 37237 8542 37252
rect 8542 37237 8545 37252
rect 8570 37237 8608 37252
rect 8608 37237 8626 37252
rect 8489 37222 8545 37237
rect 8570 37222 8626 37237
rect 8489 37196 8490 37222
rect 8490 37196 8542 37222
rect 8542 37196 8545 37222
rect 8570 37196 8608 37222
rect 8608 37196 8626 37222
rect 8651 37196 8707 37252
rect 8732 37196 8788 37252
rect 8813 37196 8869 37252
rect 8894 37196 8950 37252
rect 8975 37196 9031 37252
rect 9056 37237 9096 37252
rect 9096 37237 9110 37252
rect 9110 37237 9112 37252
rect 9137 37237 9162 37252
rect 9162 37237 9193 37252
rect 9056 37222 9112 37237
rect 9137 37222 9193 37237
rect 9056 37196 9096 37222
rect 9096 37196 9110 37222
rect 9110 37196 9112 37222
rect 9137 37196 9162 37222
rect 9162 37196 9193 37222
rect 9218 37196 9274 37252
rect 9299 37196 9355 37252
rect 9380 37196 9436 37252
rect 9461 37196 9517 37252
rect 9542 37237 9598 37289
rect 9598 37237 9650 37289
rect 9650 37237 9664 37289
rect 9664 37237 9716 37289
rect 9716 37237 9758 37289
rect 9983 37276 10039 37332
rect 10064 37276 10120 37332
rect 10145 37304 10152 37332
rect 10152 37304 10201 37332
rect 10226 37304 10270 37332
rect 10270 37304 10282 37332
rect 10145 37289 10201 37304
rect 10226 37289 10282 37304
rect 10145 37276 10152 37289
rect 10152 37276 10201 37289
rect 9542 37222 9758 37237
rect 8003 37170 8054 37172
rect 8054 37170 8059 37172
rect 7922 37155 7978 37170
rect 8003 37155 8059 37170
rect 7922 37116 7936 37155
rect 7936 37116 7978 37155
rect 8003 37116 8054 37155
rect 8054 37116 8059 37155
rect 8084 37116 8140 37172
rect 8165 37116 8221 37172
rect 8246 37116 8302 37172
rect 8327 37116 8383 37172
rect 8408 37116 8464 37172
rect 8489 37170 8490 37172
rect 8490 37170 8542 37172
rect 8542 37170 8545 37172
rect 8570 37170 8608 37172
rect 8608 37170 8626 37172
rect 8489 37155 8545 37170
rect 8570 37155 8626 37170
rect 8489 37116 8490 37155
rect 8490 37116 8542 37155
rect 8542 37116 8545 37155
rect 8570 37116 8608 37155
rect 8608 37116 8626 37155
rect 8651 37116 8707 37172
rect 8732 37116 8788 37172
rect 8813 37116 8869 37172
rect 8894 37116 8950 37172
rect 8975 37116 9031 37172
rect 9056 37170 9096 37172
rect 9096 37170 9110 37172
rect 9110 37170 9112 37172
rect 9137 37170 9162 37172
rect 9162 37170 9193 37172
rect 9056 37155 9112 37170
rect 9137 37155 9193 37170
rect 9056 37116 9096 37155
rect 9096 37116 9110 37155
rect 9110 37116 9112 37155
rect 9137 37116 9162 37155
rect 9162 37116 9193 37155
rect 9218 37116 9274 37172
rect 9299 37116 9355 37172
rect 9380 37116 9436 37172
rect 9461 37116 9517 37172
rect 9542 37170 9598 37222
rect 9598 37170 9650 37222
rect 9650 37170 9664 37222
rect 9664 37170 9716 37222
rect 9716 37170 9758 37222
rect 9983 37196 10039 37252
rect 10064 37196 10120 37252
rect 10145 37237 10152 37252
rect 10152 37237 10201 37252
rect 10226 37276 10270 37289
rect 10270 37276 10282 37289
rect 10307 37276 10363 37332
rect 10388 37276 10444 37332
rect 10469 37276 10525 37332
rect 10550 37276 10606 37332
rect 10631 37276 10687 37332
rect 10712 37304 10758 37332
rect 10758 37304 10768 37332
rect 10793 37304 10824 37332
rect 10824 37304 10849 37332
rect 10712 37289 10768 37304
rect 10793 37289 10849 37304
rect 10712 37276 10758 37289
rect 10758 37276 10768 37289
rect 10793 37276 10824 37289
rect 10824 37276 10849 37289
rect 10874 37276 10930 37332
rect 10955 37276 11011 37332
rect 11036 37276 11092 37332
rect 11117 37276 11173 37332
rect 11198 37276 11254 37332
rect 11279 37304 11312 37332
rect 11312 37304 11326 37332
rect 11326 37304 11335 37332
rect 11360 37304 11378 37332
rect 11378 37304 11416 37332
rect 11279 37289 11335 37304
rect 11360 37289 11416 37304
rect 11279 37276 11312 37289
rect 11312 37276 11326 37289
rect 11326 37276 11335 37289
rect 11360 37276 11378 37289
rect 11378 37276 11416 37289
rect 11441 37304 11814 37356
rect 11814 37304 11866 37356
rect 11866 37304 11880 37356
rect 11880 37304 11932 37356
rect 11932 37304 12057 37356
rect 11441 37289 12057 37304
rect 10226 37237 10270 37252
rect 10270 37237 10282 37252
rect 10145 37222 10201 37237
rect 10226 37222 10282 37237
rect 10145 37196 10152 37222
rect 10152 37196 10201 37222
rect 9542 37155 9758 37170
rect 9542 37103 9598 37155
rect 9598 37103 9650 37155
rect 9650 37103 9664 37155
rect 9664 37103 9716 37155
rect 9716 37103 9758 37155
rect 9983 37116 10039 37172
rect 10064 37116 10120 37172
rect 10145 37170 10152 37172
rect 10152 37170 10201 37172
rect 10226 37196 10270 37222
rect 10270 37196 10282 37222
rect 10307 37196 10363 37252
rect 10388 37196 10444 37252
rect 10469 37196 10525 37252
rect 10550 37196 10606 37252
rect 10631 37196 10687 37252
rect 10712 37237 10758 37252
rect 10758 37237 10768 37252
rect 10793 37237 10824 37252
rect 10824 37237 10849 37252
rect 10712 37222 10768 37237
rect 10793 37222 10849 37237
rect 10712 37196 10758 37222
rect 10758 37196 10768 37222
rect 10793 37196 10824 37222
rect 10824 37196 10849 37222
rect 10874 37196 10930 37252
rect 10955 37196 11011 37252
rect 11036 37196 11092 37252
rect 11117 37196 11173 37252
rect 11198 37196 11254 37252
rect 11279 37237 11312 37252
rect 11312 37237 11326 37252
rect 11326 37237 11335 37252
rect 11360 37237 11378 37252
rect 11378 37237 11416 37252
rect 11279 37222 11335 37237
rect 11360 37222 11416 37237
rect 11279 37196 11312 37222
rect 11312 37196 11326 37222
rect 11326 37196 11335 37222
rect 11360 37196 11378 37222
rect 11378 37196 11416 37222
rect 11441 37237 11814 37289
rect 11814 37237 11866 37289
rect 11866 37237 11880 37289
rect 11880 37237 11932 37289
rect 11932 37237 12057 37289
rect 11441 37222 12057 37237
rect 10226 37170 10270 37172
rect 10270 37170 10282 37172
rect 10145 37155 10201 37170
rect 10226 37155 10282 37170
rect 10145 37116 10152 37155
rect 10152 37116 10201 37155
rect 10226 37116 10270 37155
rect 10270 37116 10282 37155
rect 10307 37116 10363 37172
rect 10388 37116 10444 37172
rect 10469 37116 10525 37172
rect 10550 37116 10606 37172
rect 10631 37116 10687 37172
rect 10712 37170 10758 37172
rect 10758 37170 10768 37172
rect 10793 37170 10824 37172
rect 10824 37170 10849 37172
rect 10712 37155 10768 37170
rect 10793 37155 10849 37170
rect 10712 37116 10758 37155
rect 10758 37116 10768 37155
rect 10793 37116 10824 37155
rect 10824 37116 10849 37155
rect 10874 37116 10930 37172
rect 10955 37116 11011 37172
rect 11036 37116 11092 37172
rect 11117 37116 11173 37172
rect 11198 37116 11254 37172
rect 11279 37170 11312 37172
rect 11312 37170 11326 37172
rect 11326 37170 11335 37172
rect 11360 37170 11378 37172
rect 11378 37170 11416 37172
rect 11279 37155 11335 37170
rect 11360 37155 11416 37170
rect 11279 37116 11312 37155
rect 11312 37116 11326 37155
rect 11326 37116 11335 37155
rect 11360 37116 11378 37155
rect 11378 37116 11416 37155
rect 11441 37170 11814 37222
rect 11814 37170 11866 37222
rect 11866 37170 11880 37222
rect 11880 37170 11932 37222
rect 11932 37170 12057 37222
rect 11441 37155 12057 37170
rect 11441 37103 11814 37155
rect 11814 37103 11866 37155
rect 11866 37103 11880 37155
rect 11880 37103 11932 37155
rect 11932 37103 12057 37155
rect 7598 37036 7654 37092
rect 7679 37036 7735 37092
rect 7760 37036 7816 37092
rect 7841 37036 7897 37092
rect 7922 37088 7978 37092
rect 8003 37088 8059 37092
rect 7922 37036 7936 37088
rect 7936 37036 7978 37088
rect 8003 37036 8054 37088
rect 8054 37036 8059 37088
rect 8084 37036 8140 37092
rect 8165 37036 8221 37092
rect 8246 37036 8302 37092
rect 8327 37036 8383 37092
rect 8408 37036 8464 37092
rect 8489 37088 8545 37092
rect 8570 37088 8626 37092
rect 8489 37036 8490 37088
rect 8490 37036 8542 37088
rect 8542 37036 8545 37088
rect 8570 37036 8608 37088
rect 8608 37036 8626 37088
rect 8651 37036 8707 37092
rect 8732 37036 8788 37092
rect 8813 37036 8869 37092
rect 8894 37036 8950 37092
rect 8975 37036 9031 37092
rect 9056 37088 9112 37092
rect 9137 37088 9193 37092
rect 9056 37036 9096 37088
rect 9096 37036 9110 37088
rect 9110 37036 9112 37088
rect 9137 37036 9162 37088
rect 9162 37036 9193 37088
rect 9218 37036 9274 37092
rect 9299 37036 9355 37092
rect 9380 37036 9436 37092
rect 9461 37036 9517 37092
rect 9542 37088 9758 37103
rect 9542 37036 9598 37088
rect 9598 37036 9650 37088
rect 9650 37036 9664 37088
rect 9664 37036 9716 37088
rect 9716 37036 9758 37088
rect 9983 37036 10039 37092
rect 10064 37036 10120 37092
rect 10145 37088 10201 37092
rect 10226 37088 10282 37092
rect 10145 37036 10152 37088
rect 10152 37036 10201 37088
rect 10226 37036 10270 37088
rect 10270 37036 10282 37088
rect 10307 37036 10363 37092
rect 10388 37036 10444 37092
rect 10469 37036 10525 37092
rect 10550 37036 10606 37092
rect 10631 37036 10687 37092
rect 10712 37088 10768 37092
rect 10793 37088 10849 37092
rect 10712 37036 10758 37088
rect 10758 37036 10768 37088
rect 10793 37036 10824 37088
rect 10824 37036 10849 37088
rect 10874 37036 10930 37092
rect 10955 37036 11011 37092
rect 11036 37036 11092 37092
rect 11117 37036 11173 37092
rect 11198 37036 11254 37092
rect 11279 37088 11335 37092
rect 11360 37088 11416 37092
rect 11279 37036 11312 37088
rect 11312 37036 11326 37088
rect 11326 37036 11335 37088
rect 11360 37036 11378 37088
rect 11378 37036 11416 37088
rect 11441 37088 12057 37103
rect 11441 37036 11814 37088
rect 11814 37036 11866 37088
rect 11866 37036 11880 37088
rect 11880 37036 11932 37088
rect 11932 37036 12057 37088
rect 3513 35892 3569 35896
rect 3593 35892 3649 35896
rect 3513 35840 3556 35892
rect 3556 35840 3569 35892
rect 3593 35840 3622 35892
rect 3622 35840 3649 35892
rect 3673 35840 3729 35896
rect 3753 35840 3809 35896
rect 3833 35840 3889 35896
rect 3913 35840 3969 35896
rect 3993 35840 4049 35896
rect 4073 35892 4129 35896
rect 4153 35892 4209 35896
rect 4073 35840 4110 35892
rect 4110 35840 4124 35892
rect 4124 35840 4129 35892
rect 4153 35840 4176 35892
rect 4176 35840 4209 35892
rect 4233 35840 4289 35896
rect 4314 35840 4370 35896
rect 4395 35840 4451 35896
rect 4476 35840 4532 35896
rect 4557 35892 4613 35896
rect 4638 35892 4694 35896
rect 4719 35892 4775 35896
rect 4557 35840 4612 35892
rect 4612 35840 4613 35892
rect 4638 35840 4664 35892
rect 4664 35840 4678 35892
rect 4678 35840 4694 35892
rect 4719 35840 4730 35892
rect 4730 35840 4775 35892
rect 4800 35840 4856 35896
rect 4881 35840 4937 35896
rect 4962 35840 5018 35896
rect 5215 35840 5218 35877
rect 5218 35840 5232 35877
rect 5232 35840 5271 35877
rect 5215 35826 5271 35840
rect 5215 35821 5218 35826
rect 5218 35821 5232 35826
rect 5232 35821 5271 35826
rect 5296 35821 5352 35877
rect 5377 35821 5433 35877
rect 5458 35821 5514 35877
rect 5539 35821 5595 35877
rect 5620 35821 5676 35877
rect 5701 35840 5720 35877
rect 5720 35840 5757 35877
rect 5782 35840 5786 35877
rect 5786 35840 5838 35877
rect 5701 35826 5757 35840
rect 5782 35826 5838 35840
rect 5701 35821 5720 35826
rect 5720 35821 5757 35826
rect 5782 35821 5786 35826
rect 5786 35821 5838 35826
rect 5863 35821 5919 35877
rect 5944 35821 6000 35877
rect 6025 35821 6081 35877
rect 6106 35821 6162 35877
rect 6187 35821 6243 35877
rect 6268 35840 6274 35877
rect 6274 35840 6324 35877
rect 6349 35840 6392 35877
rect 6392 35840 6405 35877
rect 6268 35826 6324 35840
rect 6349 35826 6405 35840
rect 6268 35821 6274 35826
rect 6274 35821 6324 35826
rect 3513 35774 3556 35802
rect 3556 35774 3569 35802
rect 3593 35774 3622 35802
rect 3622 35774 3649 35802
rect 3513 35760 3569 35774
rect 3593 35760 3649 35774
rect 3513 35746 3556 35760
rect 3556 35746 3569 35760
rect 3593 35746 3622 35760
rect 3622 35746 3649 35760
rect 3673 35746 3729 35802
rect 3753 35746 3809 35802
rect 3833 35746 3889 35802
rect 3913 35746 3969 35802
rect 3993 35746 4049 35802
rect 4073 35774 4110 35802
rect 4110 35774 4124 35802
rect 4124 35774 4129 35802
rect 4153 35774 4176 35802
rect 4176 35774 4209 35802
rect 4073 35760 4129 35774
rect 4153 35760 4209 35774
rect 4073 35746 4110 35760
rect 4110 35746 4124 35760
rect 4124 35746 4129 35760
rect 4153 35746 4176 35760
rect 4176 35746 4209 35760
rect 4233 35746 4289 35802
rect 4314 35746 4370 35802
rect 4395 35746 4451 35802
rect 4476 35746 4532 35802
rect 4557 35774 4612 35802
rect 4612 35774 4613 35802
rect 4638 35774 4664 35802
rect 4664 35774 4678 35802
rect 4678 35774 4694 35802
rect 4719 35774 4730 35802
rect 4730 35774 4775 35802
rect 4557 35760 4613 35774
rect 4638 35760 4694 35774
rect 4719 35760 4775 35774
rect 4557 35746 4612 35760
rect 4612 35746 4613 35760
rect 4638 35746 4664 35760
rect 4664 35746 4678 35760
rect 4678 35746 4694 35760
rect 4719 35746 4730 35760
rect 4730 35746 4775 35760
rect 4800 35746 4856 35802
rect 4881 35746 4937 35802
rect 4962 35746 5018 35802
rect 5215 35774 5218 35789
rect 5218 35774 5232 35789
rect 5232 35774 5271 35789
rect 5215 35760 5271 35774
rect 5215 35733 5218 35760
rect 5218 35733 5232 35760
rect 5232 35733 5271 35760
rect 5296 35733 5352 35789
rect 5377 35733 5433 35789
rect 5458 35733 5514 35789
rect 5539 35733 5595 35789
rect 5620 35733 5676 35789
rect 5701 35774 5720 35789
rect 5720 35774 5757 35789
rect 5782 35774 5786 35789
rect 5786 35774 5838 35789
rect 5701 35760 5757 35774
rect 5782 35760 5838 35774
rect 5701 35733 5720 35760
rect 5720 35733 5757 35760
rect 5782 35733 5786 35760
rect 5786 35733 5838 35760
rect 5863 35733 5919 35789
rect 5944 35733 6000 35789
rect 6025 35733 6081 35789
rect 6106 35733 6162 35789
rect 6187 35733 6243 35789
rect 6268 35774 6274 35789
rect 6274 35774 6324 35789
rect 6349 35821 6392 35826
rect 6392 35821 6405 35826
rect 6430 35821 6486 35877
rect 6511 35821 6567 35877
rect 6592 35821 6648 35877
rect 6673 35821 6729 35877
rect 6754 35821 6810 35877
rect 6835 35840 6880 35877
rect 6880 35840 6891 35877
rect 6916 35840 6946 35877
rect 6946 35840 6972 35877
rect 6835 35826 6891 35840
rect 6916 35826 6972 35840
rect 6835 35821 6880 35826
rect 6880 35821 6891 35826
rect 6916 35821 6946 35826
rect 6946 35821 6972 35826
rect 6997 35821 7053 35877
rect 7078 35821 7134 35877
rect 7159 35821 7215 35877
rect 7240 35821 7296 35877
rect 7320 35821 7376 35877
rect 6349 35774 6392 35789
rect 6392 35774 6405 35789
rect 6268 35760 6324 35774
rect 6349 35760 6405 35774
rect 6268 35733 6274 35760
rect 6274 35733 6324 35760
rect 6349 35733 6392 35760
rect 6392 35733 6405 35760
rect 6430 35733 6486 35789
rect 6511 35733 6567 35789
rect 6592 35733 6648 35789
rect 6673 35733 6729 35789
rect 6754 35733 6810 35789
rect 6835 35774 6880 35789
rect 6880 35774 6891 35789
rect 6916 35774 6946 35789
rect 6946 35774 6972 35789
rect 6835 35760 6891 35774
rect 6916 35760 6972 35774
rect 6835 35733 6880 35760
rect 6880 35733 6891 35760
rect 6916 35733 6946 35760
rect 6946 35733 6972 35760
rect 6997 35733 7053 35789
rect 7078 35733 7134 35789
rect 7159 35733 7215 35789
rect 7240 35733 7296 35789
rect 7320 35733 7376 35789
rect 7598 35821 7654 35877
rect 7678 35821 7734 35877
rect 7759 35821 7815 35877
rect 7840 35821 7896 35877
rect 7921 35840 7936 35877
rect 7936 35840 7977 35877
rect 8002 35840 8054 35877
rect 8054 35840 8058 35877
rect 7921 35826 7977 35840
rect 8002 35826 8058 35840
rect 7921 35821 7936 35826
rect 7936 35821 7977 35826
rect 7598 35733 7654 35789
rect 7678 35733 7734 35789
rect 7759 35733 7815 35789
rect 7840 35733 7896 35789
rect 7921 35774 7936 35789
rect 7936 35774 7977 35789
rect 8002 35821 8054 35826
rect 8054 35821 8058 35826
rect 8083 35821 8139 35877
rect 8164 35821 8220 35877
rect 8245 35821 8301 35877
rect 8326 35821 8382 35877
rect 8407 35821 8463 35877
rect 8488 35840 8490 35877
rect 8490 35840 8542 35877
rect 8542 35840 8544 35877
rect 8569 35840 8608 35877
rect 8608 35840 8625 35877
rect 8488 35826 8544 35840
rect 8569 35826 8625 35840
rect 8488 35821 8490 35826
rect 8490 35821 8542 35826
rect 8542 35821 8544 35826
rect 8569 35821 8608 35826
rect 8608 35821 8625 35826
rect 8650 35821 8706 35877
rect 8731 35821 8787 35877
rect 8812 35821 8868 35877
rect 8893 35821 8949 35877
rect 8974 35821 9030 35877
rect 9055 35840 9096 35877
rect 9096 35840 9110 35877
rect 9110 35840 9111 35877
rect 9136 35840 9162 35877
rect 9162 35840 9192 35877
rect 9055 35826 9111 35840
rect 9136 35826 9192 35840
rect 9055 35821 9096 35826
rect 9096 35821 9110 35826
rect 9110 35821 9111 35826
rect 9136 35821 9162 35826
rect 9162 35821 9192 35826
rect 9217 35821 9273 35877
rect 9298 35821 9354 35877
rect 9379 35821 9435 35877
rect 9460 35821 9516 35877
rect 9541 35821 9597 35877
rect 9622 35840 9650 35877
rect 9650 35840 9664 35877
rect 9664 35840 9678 35877
rect 9703 35840 9716 35877
rect 9716 35840 9759 35877
rect 9622 35826 9678 35840
rect 9703 35826 9759 35840
rect 9622 35821 9650 35826
rect 9650 35821 9664 35826
rect 9664 35821 9678 35826
rect 9703 35821 9716 35826
rect 9716 35821 9759 35826
rect 9983 35821 10039 35877
rect 10063 35821 10119 35877
rect 10143 35840 10152 35877
rect 10152 35840 10199 35877
rect 10223 35840 10270 35877
rect 10270 35840 10279 35877
rect 10143 35826 10199 35840
rect 10223 35826 10279 35840
rect 10143 35821 10152 35826
rect 10152 35821 10199 35826
rect 8002 35774 8054 35789
rect 8054 35774 8058 35789
rect 7921 35760 7977 35774
rect 8002 35760 8058 35774
rect 7921 35733 7936 35760
rect 7936 35733 7977 35760
rect 8002 35733 8054 35760
rect 8054 35733 8058 35760
rect 8083 35733 8139 35789
rect 8164 35733 8220 35789
rect 8245 35733 8301 35789
rect 8326 35733 8382 35789
rect 8407 35733 8463 35789
rect 8488 35774 8490 35789
rect 8490 35774 8542 35789
rect 8542 35774 8544 35789
rect 8569 35774 8608 35789
rect 8608 35774 8625 35789
rect 8488 35760 8544 35774
rect 8569 35760 8625 35774
rect 8488 35733 8490 35760
rect 8490 35733 8542 35760
rect 8542 35733 8544 35760
rect 8569 35733 8608 35760
rect 8608 35733 8625 35760
rect 8650 35733 8706 35789
rect 8731 35733 8787 35789
rect 8812 35733 8868 35789
rect 8893 35733 8949 35789
rect 8974 35733 9030 35789
rect 9055 35774 9096 35789
rect 9096 35774 9110 35789
rect 9110 35774 9111 35789
rect 9136 35774 9162 35789
rect 9162 35774 9192 35789
rect 9055 35760 9111 35774
rect 9136 35760 9192 35774
rect 9055 35733 9096 35760
rect 9096 35733 9110 35760
rect 9110 35733 9111 35760
rect 9136 35733 9162 35760
rect 9162 35733 9192 35760
rect 9217 35733 9273 35789
rect 9298 35733 9354 35789
rect 9379 35733 9435 35789
rect 9460 35733 9516 35789
rect 9541 35733 9597 35789
rect 9622 35774 9650 35789
rect 9650 35774 9664 35789
rect 9664 35774 9678 35789
rect 9703 35774 9716 35789
rect 9716 35774 9759 35789
rect 9622 35760 9678 35774
rect 9703 35760 9759 35774
rect 9622 35733 9650 35760
rect 9650 35733 9664 35760
rect 9664 35733 9678 35760
rect 9703 35733 9716 35760
rect 9716 35733 9759 35760
rect 9983 35733 10039 35789
rect 10063 35733 10119 35789
rect 10143 35774 10152 35789
rect 10152 35774 10199 35789
rect 10223 35821 10270 35826
rect 10270 35821 10279 35826
rect 10303 35821 10359 35877
rect 10383 35821 10439 35877
rect 10463 35821 10519 35877
rect 10544 35821 10600 35877
rect 10625 35821 10681 35877
rect 10706 35840 10758 35877
rect 10758 35840 10762 35877
rect 10787 35840 10824 35877
rect 10824 35840 10843 35877
rect 10706 35826 10762 35840
rect 10787 35826 10843 35840
rect 10706 35821 10758 35826
rect 10758 35821 10762 35826
rect 10787 35821 10824 35826
rect 10824 35821 10843 35826
rect 10868 35821 10924 35877
rect 10949 35821 11005 35877
rect 11030 35821 11086 35877
rect 11111 35821 11167 35877
rect 11192 35821 11248 35877
rect 11273 35840 11312 35877
rect 11312 35840 11326 35877
rect 11326 35840 11329 35877
rect 11354 35840 11378 35877
rect 11378 35840 11410 35877
rect 11273 35826 11329 35840
rect 11354 35826 11410 35840
rect 11273 35821 11312 35826
rect 11312 35821 11326 35826
rect 11326 35821 11329 35826
rect 11354 35821 11378 35826
rect 11378 35821 11410 35826
rect 11435 35821 11491 35877
rect 11516 35821 11572 35877
rect 11597 35821 11653 35877
rect 11678 35821 11734 35877
rect 11759 35840 11814 35877
rect 11814 35840 11815 35877
rect 11840 35840 11866 35877
rect 11866 35840 11880 35877
rect 11880 35840 11896 35877
rect 11921 35840 11932 35877
rect 11932 35840 11977 35877
rect 11759 35826 11815 35840
rect 11840 35826 11896 35840
rect 11921 35826 11977 35840
rect 11759 35821 11814 35826
rect 11814 35821 11815 35826
rect 11840 35821 11866 35826
rect 11866 35821 11880 35826
rect 11880 35821 11896 35826
rect 11921 35821 11932 35826
rect 11932 35821 11977 35826
rect 12002 35821 12058 35877
rect 10223 35774 10270 35789
rect 10270 35774 10279 35789
rect 10143 35760 10199 35774
rect 10223 35760 10279 35774
rect 10143 35733 10152 35760
rect 10152 35733 10199 35760
rect 10223 35733 10270 35760
rect 10270 35733 10279 35760
rect 10303 35733 10359 35789
rect 10383 35733 10439 35789
rect 10463 35733 10519 35789
rect 10544 35733 10600 35789
rect 10625 35733 10681 35789
rect 10706 35774 10758 35789
rect 10758 35774 10762 35789
rect 10787 35774 10824 35789
rect 10824 35774 10843 35789
rect 10706 35760 10762 35774
rect 10787 35760 10843 35774
rect 10706 35733 10758 35760
rect 10758 35733 10762 35760
rect 10787 35733 10824 35760
rect 10824 35733 10843 35760
rect 10868 35733 10924 35789
rect 10949 35733 11005 35789
rect 11030 35733 11086 35789
rect 11111 35733 11167 35789
rect 11192 35733 11248 35789
rect 11273 35774 11312 35789
rect 11312 35774 11326 35789
rect 11326 35774 11329 35789
rect 11354 35774 11378 35789
rect 11378 35774 11410 35789
rect 11273 35760 11329 35774
rect 11354 35760 11410 35774
rect 11273 35733 11312 35760
rect 11312 35733 11326 35760
rect 11326 35733 11329 35760
rect 11354 35733 11378 35760
rect 11378 35733 11410 35760
rect 11435 35733 11491 35789
rect 11516 35733 11572 35789
rect 11597 35733 11653 35789
rect 11678 35733 11734 35789
rect 11759 35774 11814 35789
rect 11814 35774 11815 35789
rect 11840 35774 11866 35789
rect 11866 35774 11880 35789
rect 11880 35774 11896 35789
rect 11921 35774 11932 35789
rect 11932 35774 11977 35789
rect 11759 35760 11815 35774
rect 11840 35760 11896 35774
rect 11921 35760 11977 35774
rect 11759 35733 11814 35760
rect 11814 35733 11815 35760
rect 11840 35733 11866 35760
rect 11866 35733 11880 35760
rect 11880 35733 11896 35760
rect 11921 35733 11932 35760
rect 11932 35733 11977 35760
rect 12002 35733 12058 35789
rect 3513 35694 3569 35708
rect 3593 35694 3649 35708
rect 3513 35652 3556 35694
rect 3556 35652 3569 35694
rect 3593 35652 3622 35694
rect 3622 35652 3649 35694
rect 3673 35652 3729 35708
rect 3753 35652 3809 35708
rect 3833 35652 3889 35708
rect 3913 35652 3969 35708
rect 3993 35652 4049 35708
rect 4073 35694 4129 35708
rect 4153 35694 4209 35708
rect 4073 35652 4110 35694
rect 4110 35652 4124 35694
rect 4124 35652 4129 35694
rect 4153 35652 4176 35694
rect 4176 35652 4209 35694
rect 4233 35652 4289 35708
rect 4314 35652 4370 35708
rect 4395 35652 4451 35708
rect 4476 35652 4532 35708
rect 4557 35694 4613 35708
rect 4638 35694 4694 35708
rect 4719 35694 4775 35708
rect 4557 35652 4612 35694
rect 4612 35652 4613 35694
rect 4638 35652 4664 35694
rect 4664 35652 4678 35694
rect 4678 35652 4694 35694
rect 4719 35652 4730 35694
rect 4730 35652 4775 35694
rect 4800 35652 4856 35708
rect 4881 35652 4937 35708
rect 4962 35652 5018 35708
rect 5215 35694 5271 35701
rect 5215 35645 5218 35694
rect 5218 35645 5232 35694
rect 5232 35645 5271 35694
rect 5296 35645 5352 35701
rect 5377 35645 5433 35701
rect 5458 35645 5514 35701
rect 5539 35645 5595 35701
rect 5620 35645 5676 35701
rect 5701 35694 5757 35701
rect 5782 35694 5838 35701
rect 5701 35645 5720 35694
rect 5720 35645 5757 35694
rect 5782 35645 5786 35694
rect 5786 35645 5838 35694
rect 5863 35645 5919 35701
rect 5944 35645 6000 35701
rect 6025 35645 6081 35701
rect 6106 35645 6162 35701
rect 6187 35645 6243 35701
rect 6268 35694 6324 35701
rect 6349 35694 6405 35701
rect 6268 35645 6274 35694
rect 6274 35645 6324 35694
rect 6349 35645 6392 35694
rect 6392 35645 6405 35694
rect 6430 35645 6486 35701
rect 6511 35645 6567 35701
rect 6592 35645 6648 35701
rect 6673 35645 6729 35701
rect 6754 35645 6810 35701
rect 6835 35694 6891 35701
rect 6916 35694 6972 35701
rect 6835 35645 6880 35694
rect 6880 35645 6891 35694
rect 6916 35645 6946 35694
rect 6946 35645 6972 35694
rect 6997 35645 7053 35701
rect 7078 35645 7134 35701
rect 7159 35645 7215 35701
rect 7240 35645 7296 35701
rect 7320 35645 7376 35701
rect 7598 35645 7654 35701
rect 7678 35645 7734 35701
rect 7759 35645 7815 35701
rect 7840 35645 7896 35701
rect 7921 35694 7977 35701
rect 8002 35694 8058 35701
rect 7921 35645 7936 35694
rect 7936 35645 7977 35694
rect 8002 35645 8054 35694
rect 8054 35645 8058 35694
rect 8083 35645 8139 35701
rect 8164 35645 8220 35701
rect 8245 35645 8301 35701
rect 8326 35645 8382 35701
rect 8407 35645 8463 35701
rect 8488 35694 8544 35701
rect 8569 35694 8625 35701
rect 8488 35645 8490 35694
rect 8490 35645 8542 35694
rect 8542 35645 8544 35694
rect 8569 35645 8608 35694
rect 8608 35645 8625 35694
rect 8650 35645 8706 35701
rect 8731 35645 8787 35701
rect 8812 35645 8868 35701
rect 8893 35645 8949 35701
rect 8974 35645 9030 35701
rect 9055 35694 9111 35701
rect 9136 35694 9192 35701
rect 9055 35645 9096 35694
rect 9096 35645 9110 35694
rect 9110 35645 9111 35694
rect 9136 35645 9162 35694
rect 9162 35645 9192 35694
rect 9217 35645 9273 35701
rect 9298 35645 9354 35701
rect 9379 35645 9435 35701
rect 9460 35645 9516 35701
rect 9541 35645 9597 35701
rect 9622 35694 9678 35701
rect 9703 35694 9759 35701
rect 9622 35645 9650 35694
rect 9650 35645 9664 35694
rect 9664 35645 9678 35694
rect 9703 35645 9716 35694
rect 9716 35645 9759 35694
rect 9983 35645 10039 35701
rect 10063 35645 10119 35701
rect 10143 35694 10199 35701
rect 10223 35694 10279 35701
rect 10143 35645 10152 35694
rect 10152 35645 10199 35694
rect 10223 35645 10270 35694
rect 10270 35645 10279 35694
rect 10303 35645 10359 35701
rect 10383 35645 10439 35701
rect 10463 35645 10519 35701
rect 10544 35645 10600 35701
rect 10625 35645 10681 35701
rect 10706 35694 10762 35701
rect 10787 35694 10843 35701
rect 10706 35645 10758 35694
rect 10758 35645 10762 35694
rect 10787 35645 10824 35694
rect 10824 35645 10843 35694
rect 10868 35645 10924 35701
rect 10949 35645 11005 35701
rect 11030 35645 11086 35701
rect 11111 35645 11167 35701
rect 11192 35645 11248 35701
rect 11273 35694 11329 35701
rect 11354 35694 11410 35701
rect 11273 35645 11312 35694
rect 11312 35645 11326 35694
rect 11326 35645 11329 35694
rect 11354 35645 11378 35694
rect 11378 35645 11410 35694
rect 11435 35645 11491 35701
rect 11516 35645 11572 35701
rect 11597 35645 11653 35701
rect 11678 35645 11734 35701
rect 11759 35694 11815 35701
rect 11840 35694 11896 35701
rect 11921 35694 11977 35701
rect 11759 35645 11814 35694
rect 11814 35645 11815 35694
rect 11840 35645 11866 35694
rect 11866 35645 11880 35694
rect 11880 35645 11896 35694
rect 11921 35645 11932 35694
rect 11932 35645 11977 35694
rect 12002 35645 12058 35701
rect 3513 35575 3556 35614
rect 3556 35575 3569 35614
rect 3593 35575 3622 35614
rect 3622 35575 3649 35614
rect 3513 35560 3569 35575
rect 3593 35560 3649 35575
rect 3513 35558 3556 35560
rect 3556 35558 3569 35560
rect 3593 35558 3622 35560
rect 3622 35558 3649 35560
rect 3673 35558 3729 35614
rect 3753 35558 3809 35614
rect 3833 35558 3889 35614
rect 3913 35558 3969 35614
rect 3993 35558 4049 35614
rect 4073 35575 4110 35614
rect 4110 35575 4124 35614
rect 4124 35575 4129 35614
rect 4153 35575 4176 35614
rect 4176 35575 4209 35614
rect 4073 35560 4129 35575
rect 4153 35560 4209 35575
rect 4073 35558 4110 35560
rect 4110 35558 4124 35560
rect 4124 35558 4129 35560
rect 4153 35558 4176 35560
rect 4176 35558 4209 35560
rect 4233 35558 4289 35614
rect 4314 35558 4370 35614
rect 4395 35558 4451 35614
rect 4476 35558 4532 35614
rect 4557 35575 4612 35614
rect 4612 35575 4613 35614
rect 4638 35575 4664 35614
rect 4664 35575 4678 35614
rect 4678 35575 4694 35614
rect 4719 35575 4730 35614
rect 4730 35575 4775 35614
rect 4557 35560 4613 35575
rect 4638 35560 4694 35575
rect 4719 35560 4775 35575
rect 4557 35558 4612 35560
rect 4612 35558 4613 35560
rect 4638 35558 4664 35560
rect 4664 35558 4678 35560
rect 4678 35558 4694 35560
rect 4719 35558 4730 35560
rect 4730 35558 4775 35560
rect 4800 35558 4856 35614
rect 4881 35558 4937 35614
rect 4962 35558 5018 35614
rect 5215 35575 5218 35613
rect 5218 35575 5232 35613
rect 5232 35575 5271 35613
rect 5215 35560 5271 35575
rect 5215 35557 5218 35560
rect 5218 35557 5232 35560
rect 5232 35557 5271 35560
rect 5296 35557 5352 35613
rect 5377 35557 5433 35613
rect 5458 35557 5514 35613
rect 5539 35557 5595 35613
rect 5620 35557 5676 35613
rect 5701 35575 5720 35613
rect 5720 35575 5757 35613
rect 5782 35575 5786 35613
rect 5786 35575 5838 35613
rect 5701 35560 5757 35575
rect 5782 35560 5838 35575
rect 5701 35557 5720 35560
rect 5720 35557 5757 35560
rect 5782 35557 5786 35560
rect 5786 35557 5838 35560
rect 5863 35557 5919 35613
rect 5944 35557 6000 35613
rect 6025 35557 6081 35613
rect 6106 35557 6162 35613
rect 6187 35557 6243 35613
rect 6268 35575 6274 35613
rect 6274 35575 6324 35613
rect 6349 35575 6392 35613
rect 6392 35575 6405 35613
rect 6268 35560 6324 35575
rect 6349 35560 6405 35575
rect 6268 35557 6274 35560
rect 6274 35557 6324 35560
rect 3513 35508 3556 35520
rect 3556 35508 3569 35520
rect 3593 35508 3622 35520
rect 3622 35508 3649 35520
rect 3513 35493 3569 35508
rect 3593 35493 3649 35508
rect 3513 35464 3556 35493
rect 3556 35464 3569 35493
rect 3593 35464 3622 35493
rect 3622 35464 3649 35493
rect 3673 35464 3729 35520
rect 3753 35464 3809 35520
rect 3833 35464 3889 35520
rect 3913 35464 3969 35520
rect 3993 35464 4049 35520
rect 4073 35508 4110 35520
rect 4110 35508 4124 35520
rect 4124 35508 4129 35520
rect 4153 35508 4176 35520
rect 4176 35508 4209 35520
rect 4073 35493 4129 35508
rect 4153 35493 4209 35508
rect 4073 35464 4110 35493
rect 4110 35464 4124 35493
rect 4124 35464 4129 35493
rect 4153 35464 4176 35493
rect 4176 35464 4209 35493
rect 4233 35464 4289 35520
rect 4314 35464 4370 35520
rect 4395 35464 4451 35520
rect 4476 35464 4532 35520
rect 4557 35508 4612 35520
rect 4612 35508 4613 35520
rect 4638 35508 4664 35520
rect 4664 35508 4678 35520
rect 4678 35508 4694 35520
rect 4719 35508 4730 35520
rect 4730 35508 4775 35520
rect 4557 35493 4613 35508
rect 4638 35493 4694 35508
rect 4719 35493 4775 35508
rect 4557 35464 4612 35493
rect 4612 35464 4613 35493
rect 4638 35464 4664 35493
rect 4664 35464 4678 35493
rect 4678 35464 4694 35493
rect 4719 35464 4730 35493
rect 4730 35464 4775 35493
rect 4800 35464 4856 35520
rect 4881 35464 4937 35520
rect 4962 35464 5018 35520
rect 5215 35508 5218 35525
rect 5218 35508 5232 35525
rect 5232 35508 5271 35525
rect 5215 35493 5271 35508
rect 5215 35469 5218 35493
rect 5218 35469 5232 35493
rect 5232 35469 5271 35493
rect 5296 35469 5352 35525
rect 5377 35469 5433 35525
rect 5458 35469 5514 35525
rect 5539 35469 5595 35525
rect 5620 35469 5676 35525
rect 5701 35508 5720 35525
rect 5720 35508 5757 35525
rect 5782 35508 5786 35525
rect 5786 35508 5838 35525
rect 5701 35493 5757 35508
rect 5782 35493 5838 35508
rect 5701 35469 5720 35493
rect 5720 35469 5757 35493
rect 5782 35469 5786 35493
rect 5786 35469 5838 35493
rect 5863 35469 5919 35525
rect 5944 35469 6000 35525
rect 6025 35469 6081 35525
rect 6106 35469 6162 35525
rect 6187 35469 6243 35525
rect 6268 35508 6274 35525
rect 6274 35508 6324 35525
rect 6349 35557 6392 35560
rect 6392 35557 6405 35560
rect 6430 35557 6486 35613
rect 6511 35557 6567 35613
rect 6592 35557 6648 35613
rect 6673 35557 6729 35613
rect 6754 35557 6810 35613
rect 6835 35575 6880 35613
rect 6880 35575 6891 35613
rect 6916 35575 6946 35613
rect 6946 35575 6972 35613
rect 6835 35560 6891 35575
rect 6916 35560 6972 35575
rect 6835 35557 6880 35560
rect 6880 35557 6891 35560
rect 6916 35557 6946 35560
rect 6946 35557 6972 35560
rect 6997 35557 7053 35613
rect 7078 35557 7134 35613
rect 7159 35557 7215 35613
rect 7240 35557 7296 35613
rect 7320 35557 7376 35613
rect 6349 35508 6392 35525
rect 6392 35508 6405 35525
rect 6268 35493 6324 35508
rect 6349 35493 6405 35508
rect 6268 35469 6274 35493
rect 6274 35469 6324 35493
rect 6349 35469 6392 35493
rect 6392 35469 6405 35493
rect 6430 35469 6486 35525
rect 6511 35469 6567 35525
rect 6592 35469 6648 35525
rect 6673 35469 6729 35525
rect 6754 35469 6810 35525
rect 6835 35508 6880 35525
rect 6880 35508 6891 35525
rect 6916 35508 6946 35525
rect 6946 35508 6972 35525
rect 6835 35493 6891 35508
rect 6916 35493 6972 35508
rect 6835 35469 6880 35493
rect 6880 35469 6891 35493
rect 6916 35469 6946 35493
rect 6946 35469 6972 35493
rect 6997 35469 7053 35525
rect 7078 35469 7134 35525
rect 7159 35469 7215 35525
rect 7240 35469 7296 35525
rect 7320 35469 7376 35525
rect 7598 35557 7654 35613
rect 7678 35557 7734 35613
rect 7759 35557 7815 35613
rect 7840 35557 7896 35613
rect 7921 35575 7936 35613
rect 7936 35575 7977 35613
rect 8002 35575 8054 35613
rect 8054 35575 8058 35613
rect 7921 35560 7977 35575
rect 8002 35560 8058 35575
rect 7921 35557 7936 35560
rect 7936 35557 7977 35560
rect 7598 35469 7654 35525
rect 7678 35469 7734 35525
rect 7759 35469 7815 35525
rect 7840 35469 7896 35525
rect 7921 35508 7936 35525
rect 7936 35508 7977 35525
rect 8002 35557 8054 35560
rect 8054 35557 8058 35560
rect 8083 35557 8139 35613
rect 8164 35557 8220 35613
rect 8245 35557 8301 35613
rect 8326 35557 8382 35613
rect 8407 35557 8463 35613
rect 8488 35575 8490 35613
rect 8490 35575 8542 35613
rect 8542 35575 8544 35613
rect 8569 35575 8608 35613
rect 8608 35575 8625 35613
rect 8488 35560 8544 35575
rect 8569 35560 8625 35575
rect 8488 35557 8490 35560
rect 8490 35557 8542 35560
rect 8542 35557 8544 35560
rect 8569 35557 8608 35560
rect 8608 35557 8625 35560
rect 8650 35557 8706 35613
rect 8731 35557 8787 35613
rect 8812 35557 8868 35613
rect 8893 35557 8949 35613
rect 8974 35557 9030 35613
rect 9055 35575 9096 35613
rect 9096 35575 9110 35613
rect 9110 35575 9111 35613
rect 9136 35575 9162 35613
rect 9162 35575 9192 35613
rect 9055 35560 9111 35575
rect 9136 35560 9192 35575
rect 9055 35557 9096 35560
rect 9096 35557 9110 35560
rect 9110 35557 9111 35560
rect 9136 35557 9162 35560
rect 9162 35557 9192 35560
rect 9217 35557 9273 35613
rect 9298 35557 9354 35613
rect 9379 35557 9435 35613
rect 9460 35557 9516 35613
rect 9541 35557 9597 35613
rect 9622 35575 9650 35613
rect 9650 35575 9664 35613
rect 9664 35575 9678 35613
rect 9703 35575 9716 35613
rect 9716 35575 9759 35613
rect 9622 35560 9678 35575
rect 9703 35560 9759 35575
rect 9622 35557 9650 35560
rect 9650 35557 9664 35560
rect 9664 35557 9678 35560
rect 9703 35557 9716 35560
rect 9716 35557 9759 35560
rect 9983 35557 10039 35613
rect 10063 35557 10119 35613
rect 10143 35575 10152 35613
rect 10152 35575 10199 35613
rect 10223 35575 10270 35613
rect 10270 35575 10279 35613
rect 10143 35560 10199 35575
rect 10223 35560 10279 35575
rect 10143 35557 10152 35560
rect 10152 35557 10199 35560
rect 8002 35508 8054 35525
rect 8054 35508 8058 35525
rect 7921 35493 7977 35508
rect 8002 35493 8058 35508
rect 7921 35469 7936 35493
rect 7936 35469 7977 35493
rect 8002 35469 8054 35493
rect 8054 35469 8058 35493
rect 8083 35469 8139 35525
rect 8164 35469 8220 35525
rect 8245 35469 8301 35525
rect 8326 35469 8382 35525
rect 8407 35469 8463 35525
rect 8488 35508 8490 35525
rect 8490 35508 8542 35525
rect 8542 35508 8544 35525
rect 8569 35508 8608 35525
rect 8608 35508 8625 35525
rect 8488 35493 8544 35508
rect 8569 35493 8625 35508
rect 8488 35469 8490 35493
rect 8490 35469 8542 35493
rect 8542 35469 8544 35493
rect 8569 35469 8608 35493
rect 8608 35469 8625 35493
rect 8650 35469 8706 35525
rect 8731 35469 8787 35525
rect 8812 35469 8868 35525
rect 8893 35469 8949 35525
rect 8974 35469 9030 35525
rect 9055 35508 9096 35525
rect 9096 35508 9110 35525
rect 9110 35508 9111 35525
rect 9136 35508 9162 35525
rect 9162 35508 9192 35525
rect 9055 35493 9111 35508
rect 9136 35493 9192 35508
rect 9055 35469 9096 35493
rect 9096 35469 9110 35493
rect 9110 35469 9111 35493
rect 9136 35469 9162 35493
rect 9162 35469 9192 35493
rect 9217 35469 9273 35525
rect 9298 35469 9354 35525
rect 9379 35469 9435 35525
rect 9460 35469 9516 35525
rect 9541 35469 9597 35525
rect 9622 35508 9650 35525
rect 9650 35508 9664 35525
rect 9664 35508 9678 35525
rect 9703 35508 9716 35525
rect 9716 35508 9759 35525
rect 9622 35493 9678 35508
rect 9703 35493 9759 35508
rect 9622 35469 9650 35493
rect 9650 35469 9664 35493
rect 9664 35469 9678 35493
rect 9703 35469 9716 35493
rect 9716 35469 9759 35493
rect 9983 35469 10039 35525
rect 10063 35469 10119 35525
rect 10143 35508 10152 35525
rect 10152 35508 10199 35525
rect 10223 35557 10270 35560
rect 10270 35557 10279 35560
rect 10303 35557 10359 35613
rect 10383 35557 10439 35613
rect 10463 35557 10519 35613
rect 10544 35557 10600 35613
rect 10625 35557 10681 35613
rect 10706 35575 10758 35613
rect 10758 35575 10762 35613
rect 10787 35575 10824 35613
rect 10824 35575 10843 35613
rect 10706 35560 10762 35575
rect 10787 35560 10843 35575
rect 10706 35557 10758 35560
rect 10758 35557 10762 35560
rect 10787 35557 10824 35560
rect 10824 35557 10843 35560
rect 10868 35557 10924 35613
rect 10949 35557 11005 35613
rect 11030 35557 11086 35613
rect 11111 35557 11167 35613
rect 11192 35557 11248 35613
rect 11273 35575 11312 35613
rect 11312 35575 11326 35613
rect 11326 35575 11329 35613
rect 11354 35575 11378 35613
rect 11378 35575 11410 35613
rect 11273 35560 11329 35575
rect 11354 35560 11410 35575
rect 11273 35557 11312 35560
rect 11312 35557 11326 35560
rect 11326 35557 11329 35560
rect 11354 35557 11378 35560
rect 11378 35557 11410 35560
rect 11435 35557 11491 35613
rect 11516 35557 11572 35613
rect 11597 35557 11653 35613
rect 11678 35557 11734 35613
rect 11759 35575 11814 35613
rect 11814 35575 11815 35613
rect 11840 35575 11866 35613
rect 11866 35575 11880 35613
rect 11880 35575 11896 35613
rect 11921 35575 11932 35613
rect 11932 35575 11977 35613
rect 11759 35560 11815 35575
rect 11840 35560 11896 35575
rect 11921 35560 11977 35575
rect 11759 35557 11814 35560
rect 11814 35557 11815 35560
rect 11840 35557 11866 35560
rect 11866 35557 11880 35560
rect 11880 35557 11896 35560
rect 11921 35557 11932 35560
rect 11932 35557 11977 35560
rect 12002 35557 12058 35613
rect 10223 35508 10270 35525
rect 10270 35508 10279 35525
rect 10143 35493 10199 35508
rect 10223 35493 10279 35508
rect 10143 35469 10152 35493
rect 10152 35469 10199 35493
rect 10223 35469 10270 35493
rect 10270 35469 10279 35493
rect 10303 35469 10359 35525
rect 10383 35469 10439 35525
rect 10463 35469 10519 35525
rect 10544 35469 10600 35525
rect 10625 35469 10681 35525
rect 10706 35508 10758 35525
rect 10758 35508 10762 35525
rect 10787 35508 10824 35525
rect 10824 35508 10843 35525
rect 10706 35493 10762 35508
rect 10787 35493 10843 35508
rect 10706 35469 10758 35493
rect 10758 35469 10762 35493
rect 10787 35469 10824 35493
rect 10824 35469 10843 35493
rect 10868 35469 10924 35525
rect 10949 35469 11005 35525
rect 11030 35469 11086 35525
rect 11111 35469 11167 35525
rect 11192 35469 11248 35525
rect 11273 35508 11312 35525
rect 11312 35508 11326 35525
rect 11326 35508 11329 35525
rect 11354 35508 11378 35525
rect 11378 35508 11410 35525
rect 11273 35493 11329 35508
rect 11354 35493 11410 35508
rect 11273 35469 11312 35493
rect 11312 35469 11326 35493
rect 11326 35469 11329 35493
rect 11354 35469 11378 35493
rect 11378 35469 11410 35493
rect 11435 35469 11491 35525
rect 11516 35469 11572 35525
rect 11597 35469 11653 35525
rect 11678 35469 11734 35525
rect 11759 35508 11814 35525
rect 11814 35508 11815 35525
rect 11840 35508 11866 35525
rect 11866 35508 11880 35525
rect 11880 35508 11896 35525
rect 11921 35508 11932 35525
rect 11932 35508 11977 35525
rect 11759 35493 11815 35508
rect 11840 35493 11896 35508
rect 11921 35493 11977 35508
rect 11759 35469 11814 35493
rect 11814 35469 11815 35493
rect 11840 35469 11866 35493
rect 11866 35469 11880 35493
rect 11880 35469 11896 35493
rect 11921 35469 11932 35493
rect 11932 35469 11977 35493
rect 12002 35469 12058 35525
rect 5215 35426 5271 35437
rect 3513 35374 3556 35426
rect 3556 35374 3569 35426
rect 3593 35374 3622 35426
rect 3622 35374 3649 35426
rect 3513 35370 3569 35374
rect 3593 35370 3649 35374
rect 3673 35370 3729 35426
rect 3753 35370 3809 35426
rect 3833 35370 3889 35426
rect 3913 35370 3969 35426
rect 3993 35370 4049 35426
rect 4073 35374 4110 35426
rect 4110 35374 4124 35426
rect 4124 35374 4129 35426
rect 4153 35374 4176 35426
rect 4176 35374 4209 35426
rect 4073 35370 4129 35374
rect 4153 35370 4209 35374
rect 4233 35370 4289 35426
rect 4314 35370 4370 35426
rect 4395 35370 4451 35426
rect 4476 35370 4532 35426
rect 4557 35374 4612 35426
rect 4612 35374 4613 35426
rect 4638 35374 4664 35426
rect 4664 35374 4678 35426
rect 4678 35374 4694 35426
rect 4719 35374 4730 35426
rect 4730 35374 4775 35426
rect 4557 35370 4613 35374
rect 4638 35370 4694 35374
rect 4719 35370 4775 35374
rect 4800 35370 4856 35426
rect 4881 35370 4937 35426
rect 4962 35370 5018 35426
rect 5215 35381 5218 35426
rect 5218 35381 5232 35426
rect 5232 35381 5271 35426
rect 5296 35381 5352 35437
rect 5377 35381 5433 35437
rect 5458 35381 5514 35437
rect 5539 35381 5595 35437
rect 5620 35381 5676 35437
rect 5701 35426 5757 35437
rect 5782 35426 5838 35437
rect 5701 35381 5720 35426
rect 5720 35381 5757 35426
rect 5782 35381 5786 35426
rect 5786 35381 5838 35426
rect 5863 35381 5919 35437
rect 5944 35381 6000 35437
rect 6025 35381 6081 35437
rect 6106 35381 6162 35437
rect 6187 35381 6243 35437
rect 6268 35426 6324 35437
rect 6349 35426 6405 35437
rect 6268 35381 6274 35426
rect 6274 35381 6324 35426
rect 6349 35381 6392 35426
rect 6392 35381 6405 35426
rect 6430 35381 6486 35437
rect 6511 35381 6567 35437
rect 6592 35381 6648 35437
rect 6673 35381 6729 35437
rect 6754 35381 6810 35437
rect 6835 35426 6891 35437
rect 6916 35426 6972 35437
rect 6835 35381 6880 35426
rect 6880 35381 6891 35426
rect 6916 35381 6946 35426
rect 6946 35381 6972 35426
rect 6997 35381 7053 35437
rect 7078 35381 7134 35437
rect 7159 35381 7215 35437
rect 7240 35381 7296 35437
rect 7320 35381 7376 35437
rect 7598 35381 7654 35437
rect 7678 35381 7734 35437
rect 7759 35381 7815 35437
rect 7840 35381 7896 35437
rect 7921 35426 7977 35437
rect 8002 35426 8058 35437
rect 7921 35381 7936 35426
rect 7936 35381 7977 35426
rect 8002 35381 8054 35426
rect 8054 35381 8058 35426
rect 8083 35381 8139 35437
rect 8164 35381 8220 35437
rect 8245 35381 8301 35437
rect 8326 35381 8382 35437
rect 8407 35381 8463 35437
rect 8488 35426 8544 35437
rect 8569 35426 8625 35437
rect 8488 35381 8490 35426
rect 8490 35381 8542 35426
rect 8542 35381 8544 35426
rect 8569 35381 8608 35426
rect 8608 35381 8625 35426
rect 8650 35381 8706 35437
rect 8731 35381 8787 35437
rect 8812 35381 8868 35437
rect 8893 35381 8949 35437
rect 8974 35381 9030 35437
rect 9055 35426 9111 35437
rect 9136 35426 9192 35437
rect 9055 35381 9096 35426
rect 9096 35381 9110 35426
rect 9110 35381 9111 35426
rect 9136 35381 9162 35426
rect 9162 35381 9192 35426
rect 9217 35381 9273 35437
rect 9298 35381 9354 35437
rect 9379 35381 9435 35437
rect 9460 35381 9516 35437
rect 9541 35381 9597 35437
rect 9622 35426 9678 35437
rect 9703 35426 9759 35437
rect 9622 35381 9650 35426
rect 9650 35381 9664 35426
rect 9664 35381 9678 35426
rect 9703 35381 9716 35426
rect 9716 35381 9759 35426
rect 9983 35381 10039 35437
rect 10063 35381 10119 35437
rect 10143 35426 10199 35437
rect 10223 35426 10279 35437
rect 10143 35381 10152 35426
rect 10152 35381 10199 35426
rect 10223 35381 10270 35426
rect 10270 35381 10279 35426
rect 10303 35381 10359 35437
rect 10383 35381 10439 35437
rect 10463 35381 10519 35437
rect 10544 35381 10600 35437
rect 10625 35381 10681 35437
rect 10706 35426 10762 35437
rect 10787 35426 10843 35437
rect 10706 35381 10758 35426
rect 10758 35381 10762 35426
rect 10787 35381 10824 35426
rect 10824 35381 10843 35426
rect 10868 35381 10924 35437
rect 10949 35381 11005 35437
rect 11030 35381 11086 35437
rect 11111 35381 11167 35437
rect 11192 35381 11248 35437
rect 11273 35426 11329 35437
rect 11354 35426 11410 35437
rect 11273 35381 11312 35426
rect 11312 35381 11326 35426
rect 11326 35381 11329 35426
rect 11354 35381 11378 35426
rect 11378 35381 11410 35426
rect 11435 35381 11491 35437
rect 11516 35381 11572 35437
rect 11597 35381 11653 35437
rect 11678 35381 11734 35437
rect 11759 35426 11815 35437
rect 11840 35426 11896 35437
rect 11921 35426 11977 35437
rect 11759 35381 11814 35426
rect 11814 35381 11815 35426
rect 11840 35381 11866 35426
rect 11866 35381 11880 35426
rect 11880 35381 11896 35426
rect 11921 35381 11932 35426
rect 11932 35381 11977 35426
rect 12002 35381 12058 35437
rect 3513 33840 3569 33896
rect 3594 33892 3650 33896
rect 3675 33892 3731 33896
rect 3594 33840 3637 33892
rect 3637 33840 3650 33892
rect 3675 33840 3703 33892
rect 3703 33840 3731 33892
rect 3757 33840 3813 33896
rect 3839 33840 3895 33896
rect 3921 33840 3977 33896
rect 4003 33840 4059 33896
rect 4085 33840 4141 33896
rect 4167 33840 4223 33896
rect 4249 33840 4305 33896
rect 4354 33824 4410 33880
rect 4446 33840 4473 33880
rect 4473 33840 4487 33880
rect 4487 33840 4502 33880
rect 4446 33826 4502 33840
rect 4556 33830 4612 33886
rect 5216 33840 5257 33878
rect 5257 33840 5272 33878
rect 5299 33840 5309 33878
rect 5309 33840 5323 33878
rect 5323 33840 5355 33878
rect 5216 33826 5272 33840
rect 5299 33826 5355 33840
rect 4446 33824 4473 33826
rect 4473 33824 4487 33826
rect 4487 33824 4502 33826
rect 3513 33746 3569 33802
rect 3594 33774 3637 33802
rect 3637 33774 3650 33802
rect 3675 33774 3703 33802
rect 3703 33774 3731 33802
rect 3594 33760 3650 33774
rect 3675 33760 3731 33774
rect 3594 33746 3637 33760
rect 3637 33746 3650 33760
rect 3675 33746 3703 33760
rect 3703 33746 3731 33760
rect 3757 33746 3813 33802
rect 3839 33746 3895 33802
rect 3921 33746 3977 33802
rect 4003 33746 4059 33802
rect 4085 33746 4141 33802
rect 4167 33746 4223 33802
rect 4249 33746 4305 33802
rect 5216 33822 5257 33826
rect 5257 33822 5272 33826
rect 5299 33822 5309 33826
rect 5309 33822 5323 33826
rect 5323 33822 5355 33826
rect 5382 33822 5438 33878
rect 5465 33822 5521 33878
rect 5548 33822 5604 33878
rect 5631 33822 5687 33878
rect 5714 33822 5770 33878
rect 5797 33822 5853 33878
rect 5880 33822 5936 33878
rect 5963 33822 6019 33878
rect 6046 33840 6093 33878
rect 6093 33840 6102 33878
rect 6129 33840 6145 33878
rect 6145 33840 6159 33878
rect 6159 33840 6185 33878
rect 6046 33826 6102 33840
rect 6129 33826 6185 33840
rect 6046 33822 6093 33826
rect 6093 33822 6102 33826
rect 6129 33822 6145 33826
rect 6145 33822 6159 33826
rect 6159 33822 6185 33826
rect 6211 33822 6267 33878
rect 6293 33822 6349 33878
rect 6375 33822 6431 33878
rect 6457 33822 6513 33878
rect 6539 33822 6595 33878
rect 6621 33822 6677 33878
rect 6703 33822 6759 33878
rect 6785 33822 6841 33878
rect 6867 33822 6923 33878
rect 6949 33840 6981 33878
rect 6981 33840 6995 33878
rect 6995 33840 7005 33878
rect 7031 33840 7047 33878
rect 7047 33840 7087 33878
rect 6949 33826 7005 33840
rect 7031 33826 7087 33840
rect 6949 33822 6981 33826
rect 6981 33822 6995 33826
rect 6995 33822 7005 33826
rect 7031 33822 7047 33826
rect 7047 33822 7087 33826
rect 7113 33822 7169 33878
rect 7195 33822 7251 33878
rect 4354 33724 4410 33780
rect 4446 33774 4473 33780
rect 4473 33774 4487 33780
rect 4487 33774 4502 33780
rect 4446 33760 4502 33774
rect 4446 33724 4473 33760
rect 4473 33724 4487 33760
rect 4487 33724 4502 33760
rect 4556 33748 4612 33804
rect 7636 33802 7692 33858
rect 7716 33840 7765 33858
rect 7765 33840 7772 33858
rect 7838 33840 7883 33881
rect 7883 33840 7894 33881
rect 7716 33826 7772 33840
rect 7838 33826 7894 33840
rect 7716 33802 7765 33826
rect 7765 33802 7772 33826
rect 5216 33774 5257 33790
rect 5257 33774 5272 33790
rect 5299 33774 5309 33790
rect 5309 33774 5323 33790
rect 5323 33774 5355 33790
rect 5216 33760 5272 33774
rect 5299 33760 5355 33774
rect 5216 33734 5257 33760
rect 5257 33734 5272 33760
rect 5299 33734 5309 33760
rect 5309 33734 5323 33760
rect 5323 33734 5355 33760
rect 5382 33734 5438 33790
rect 5465 33734 5521 33790
rect 5548 33734 5604 33790
rect 5631 33734 5687 33790
rect 5714 33734 5770 33790
rect 5797 33734 5853 33790
rect 5880 33734 5936 33790
rect 5963 33734 6019 33790
rect 6046 33774 6093 33790
rect 6093 33774 6102 33790
rect 6129 33774 6145 33790
rect 6145 33774 6159 33790
rect 6159 33774 6185 33790
rect 6046 33760 6102 33774
rect 6129 33760 6185 33774
rect 6046 33734 6093 33760
rect 6093 33734 6102 33760
rect 6129 33734 6145 33760
rect 6145 33734 6159 33760
rect 6159 33734 6185 33760
rect 6211 33734 6267 33790
rect 6293 33734 6349 33790
rect 6375 33734 6431 33790
rect 6457 33734 6513 33790
rect 6539 33734 6595 33790
rect 6621 33734 6677 33790
rect 6703 33734 6759 33790
rect 6785 33734 6841 33790
rect 6867 33734 6923 33790
rect 6949 33774 6981 33790
rect 6981 33774 6995 33790
rect 6995 33774 7005 33790
rect 7031 33774 7047 33790
rect 7047 33774 7087 33790
rect 6949 33760 7005 33774
rect 7031 33760 7087 33774
rect 6949 33734 6981 33760
rect 6981 33734 6995 33760
rect 6995 33734 7005 33760
rect 7031 33734 7047 33760
rect 7047 33734 7087 33760
rect 7113 33734 7169 33790
rect 7195 33734 7251 33790
rect 7838 33825 7883 33826
rect 7883 33825 7894 33826
rect 7922 33825 7978 33881
rect 8041 33822 8097 33878
rect 8124 33822 8180 33878
rect 8207 33822 8263 33878
rect 8290 33822 8346 33878
rect 8373 33822 8429 33878
rect 8456 33822 8512 33878
rect 8539 33822 8595 33878
rect 8622 33840 8653 33878
rect 8653 33840 8667 33878
rect 8667 33840 8678 33878
rect 8705 33840 8719 33878
rect 8719 33840 8761 33878
rect 8622 33826 8678 33840
rect 8705 33826 8761 33840
rect 8622 33822 8653 33826
rect 8653 33822 8667 33826
rect 8667 33822 8678 33826
rect 8705 33822 8719 33826
rect 8719 33822 8761 33826
rect 8788 33822 8844 33878
rect 8871 33822 8927 33878
rect 8954 33822 9010 33878
rect 9037 33822 9093 33878
rect 9120 33822 9176 33878
rect 9203 33822 9259 33878
rect 9286 33822 9342 33878
rect 9369 33822 9425 33878
rect 9452 33840 9489 33878
rect 9489 33840 9503 33878
rect 9503 33840 9508 33878
rect 9535 33840 9555 33878
rect 9555 33840 9591 33878
rect 9452 33826 9508 33840
rect 9535 33826 9591 33840
rect 9452 33822 9489 33826
rect 9489 33822 9503 33826
rect 9503 33822 9508 33826
rect 9535 33822 9555 33826
rect 9555 33822 9591 33826
rect 9618 33822 9674 33878
rect 9702 33822 9758 33878
rect 10000 33802 10056 33858
rect 10080 33802 10136 33858
rect 10202 33825 10258 33881
rect 10286 33840 10325 33881
rect 10325 33840 10339 33881
rect 10339 33840 10342 33881
rect 10286 33826 10342 33840
rect 10286 33825 10325 33826
rect 10325 33825 10339 33826
rect 10339 33825 10342 33826
rect 7838 33760 7894 33766
rect 7723 33708 7765 33751
rect 7765 33708 7779 33751
rect 7838 33710 7883 33760
rect 7883 33710 7894 33760
rect 7922 33710 7978 33766
rect 8041 33734 8097 33790
rect 8124 33734 8180 33790
rect 8207 33734 8263 33790
rect 8290 33734 8346 33790
rect 8373 33734 8429 33790
rect 8456 33734 8512 33790
rect 8539 33734 8595 33790
rect 8622 33774 8653 33790
rect 8653 33774 8667 33790
rect 8667 33774 8678 33790
rect 8705 33774 8719 33790
rect 8719 33774 8761 33790
rect 8622 33760 8678 33774
rect 8705 33760 8761 33774
rect 8622 33734 8653 33760
rect 8653 33734 8667 33760
rect 8667 33734 8678 33760
rect 8705 33734 8719 33760
rect 8719 33734 8761 33760
rect 8788 33734 8844 33790
rect 8871 33734 8927 33790
rect 8954 33734 9010 33790
rect 9037 33734 9093 33790
rect 9120 33734 9176 33790
rect 9203 33734 9259 33790
rect 9286 33734 9342 33790
rect 9369 33734 9425 33790
rect 9452 33774 9489 33790
rect 9489 33774 9503 33790
rect 9503 33774 9508 33790
rect 9535 33774 9555 33790
rect 9555 33774 9591 33790
rect 9452 33760 9508 33774
rect 9535 33760 9591 33774
rect 9452 33734 9489 33760
rect 9489 33734 9503 33760
rect 9503 33734 9508 33760
rect 9535 33734 9555 33760
rect 9555 33734 9591 33760
rect 9618 33734 9674 33790
rect 9702 33734 9758 33790
rect 10397 33822 10453 33878
rect 10477 33822 10533 33878
rect 10557 33822 10613 33878
rect 10637 33822 10693 33878
rect 10717 33822 10773 33878
rect 10797 33822 10853 33878
rect 10877 33822 10933 33878
rect 10957 33822 11013 33878
rect 11037 33822 11093 33878
rect 11117 33840 11161 33878
rect 11161 33840 11173 33878
rect 11197 33840 11227 33878
rect 11227 33840 11253 33878
rect 11117 33826 11173 33840
rect 11197 33826 11253 33840
rect 11117 33822 11161 33826
rect 11161 33822 11173 33826
rect 11197 33822 11227 33826
rect 11227 33822 11253 33826
rect 11277 33822 11333 33878
rect 11357 33822 11413 33878
rect 11437 33822 11493 33878
rect 11517 33822 11573 33878
rect 11597 33822 11653 33878
rect 11677 33822 11733 33878
rect 11758 33822 11814 33878
rect 11839 33822 11895 33878
rect 11920 33840 11945 33878
rect 11945 33840 11976 33878
rect 12001 33840 12011 33878
rect 12011 33840 12057 33878
rect 11920 33826 11976 33840
rect 12001 33826 12057 33840
rect 11920 33822 11945 33826
rect 11945 33822 11976 33826
rect 12001 33822 12011 33826
rect 12011 33822 12057 33826
rect 3513 33652 3569 33708
rect 3594 33694 3650 33708
rect 3675 33694 3731 33708
rect 3594 33652 3637 33694
rect 3637 33652 3650 33694
rect 3675 33652 3703 33694
rect 3703 33652 3731 33694
rect 3757 33652 3813 33708
rect 3839 33652 3895 33708
rect 3921 33652 3977 33708
rect 4003 33652 4059 33708
rect 4085 33652 4141 33708
rect 4167 33652 4223 33708
rect 4249 33652 4305 33708
rect 5216 33694 5272 33702
rect 5299 33694 5355 33702
rect 4354 33623 4410 33679
rect 4446 33642 4473 33679
rect 4473 33642 4487 33679
rect 4487 33642 4502 33679
rect 5216 33646 5257 33694
rect 5257 33646 5272 33694
rect 5299 33646 5309 33694
rect 5309 33646 5323 33694
rect 5323 33646 5355 33694
rect 5382 33646 5438 33702
rect 5465 33646 5521 33702
rect 5548 33646 5604 33702
rect 5631 33646 5687 33702
rect 5714 33646 5770 33702
rect 5797 33646 5853 33702
rect 5880 33646 5936 33702
rect 5963 33646 6019 33702
rect 6046 33694 6102 33702
rect 6129 33694 6185 33702
rect 6046 33646 6093 33694
rect 6093 33646 6102 33694
rect 6129 33646 6145 33694
rect 6145 33646 6159 33694
rect 6159 33646 6185 33694
rect 6211 33646 6267 33702
rect 6293 33646 6349 33702
rect 6375 33646 6431 33702
rect 6457 33646 6513 33702
rect 6539 33646 6595 33702
rect 6621 33646 6677 33702
rect 6703 33646 6759 33702
rect 6785 33646 6841 33702
rect 6867 33646 6923 33702
rect 6949 33694 7005 33702
rect 7031 33694 7087 33702
rect 6949 33646 6981 33694
rect 6981 33646 6995 33694
rect 6995 33646 7005 33694
rect 7031 33646 7047 33694
rect 7047 33646 7087 33694
rect 7113 33646 7169 33702
rect 7195 33646 7251 33702
rect 7723 33695 7779 33708
rect 7838 33642 7883 33650
rect 7883 33642 7894 33650
rect 4446 33627 4502 33642
rect 7838 33627 7894 33642
rect 4446 33623 4473 33627
rect 4473 33623 4487 33627
rect 4487 33623 4502 33627
rect 3513 33558 3569 33614
rect 3594 33575 3637 33614
rect 3637 33575 3650 33614
rect 3675 33575 3703 33614
rect 3703 33575 3731 33614
rect 3594 33560 3650 33575
rect 3675 33560 3731 33575
rect 3594 33558 3637 33560
rect 3637 33558 3650 33560
rect 3675 33558 3703 33560
rect 3703 33558 3731 33560
rect 3757 33558 3813 33614
rect 3839 33558 3895 33614
rect 3921 33558 3977 33614
rect 4003 33558 4059 33614
rect 4085 33558 4141 33614
rect 4167 33558 4223 33614
rect 4249 33558 4305 33614
rect 5216 33575 5257 33614
rect 5257 33575 5272 33614
rect 5299 33575 5309 33614
rect 5309 33575 5323 33614
rect 5323 33575 5355 33614
rect 5216 33560 5272 33575
rect 5299 33560 5355 33575
rect 3513 33464 3569 33520
rect 3594 33508 3637 33520
rect 3637 33508 3650 33520
rect 3675 33508 3703 33520
rect 3703 33508 3731 33520
rect 3594 33493 3650 33508
rect 3675 33493 3731 33508
rect 3594 33464 3637 33493
rect 3637 33464 3650 33493
rect 3675 33464 3703 33493
rect 3703 33464 3731 33493
rect 3757 33464 3813 33520
rect 3839 33464 3895 33520
rect 3921 33464 3977 33520
rect 4003 33464 4059 33520
rect 4085 33464 4141 33520
rect 4167 33464 4223 33520
rect 4249 33464 4305 33520
rect 5216 33558 5257 33560
rect 5257 33558 5272 33560
rect 5299 33558 5309 33560
rect 5309 33558 5323 33560
rect 5323 33558 5355 33560
rect 5382 33558 5438 33614
rect 5465 33558 5521 33614
rect 5548 33558 5604 33614
rect 5631 33558 5687 33614
rect 5714 33558 5770 33614
rect 5797 33558 5853 33614
rect 5880 33558 5936 33614
rect 5963 33558 6019 33614
rect 6046 33575 6093 33614
rect 6093 33575 6102 33614
rect 6129 33575 6145 33614
rect 6145 33575 6159 33614
rect 6159 33575 6185 33614
rect 6046 33560 6102 33575
rect 6129 33560 6185 33575
rect 6046 33558 6093 33560
rect 6093 33558 6102 33560
rect 6129 33558 6145 33560
rect 6145 33558 6159 33560
rect 6159 33558 6185 33560
rect 6211 33558 6267 33614
rect 6293 33558 6349 33614
rect 6375 33558 6431 33614
rect 6457 33558 6513 33614
rect 6539 33558 6595 33614
rect 6621 33558 6677 33614
rect 6703 33558 6759 33614
rect 6785 33558 6841 33614
rect 6867 33558 6923 33614
rect 6949 33575 6981 33614
rect 6981 33575 6995 33614
rect 6995 33575 7005 33614
rect 7031 33575 7047 33614
rect 7047 33575 7087 33614
rect 6949 33560 7005 33575
rect 7031 33560 7087 33575
rect 6949 33558 6981 33560
rect 6981 33558 6995 33560
rect 6995 33558 7005 33560
rect 7031 33558 7047 33560
rect 7047 33558 7087 33560
rect 7113 33558 7169 33614
rect 7195 33558 7251 33614
rect 7838 33594 7883 33627
rect 7883 33594 7894 33627
rect 7922 33594 7978 33650
rect 8041 33646 8097 33702
rect 8124 33646 8180 33702
rect 8207 33646 8263 33702
rect 8290 33646 8346 33702
rect 8373 33646 8429 33702
rect 8456 33646 8512 33702
rect 8539 33646 8595 33702
rect 8622 33694 8678 33702
rect 8705 33694 8761 33702
rect 8622 33646 8653 33694
rect 8653 33646 8667 33694
rect 8667 33646 8678 33694
rect 8705 33646 8719 33694
rect 8719 33646 8761 33694
rect 8788 33646 8844 33702
rect 8871 33646 8927 33702
rect 8954 33646 9010 33702
rect 9037 33646 9093 33702
rect 9120 33646 9176 33702
rect 9203 33646 9259 33702
rect 9286 33646 9342 33702
rect 9369 33646 9425 33702
rect 9452 33694 9508 33702
rect 9535 33694 9591 33702
rect 9452 33646 9489 33694
rect 9489 33646 9503 33694
rect 9503 33646 9508 33694
rect 9535 33646 9555 33694
rect 9555 33646 9591 33694
rect 9618 33646 9674 33702
rect 9702 33646 9758 33702
rect 10087 33695 10143 33751
rect 10202 33710 10258 33766
rect 10286 33760 10342 33766
rect 10286 33710 10325 33760
rect 10325 33710 10339 33760
rect 10339 33710 10342 33760
rect 10397 33734 10453 33790
rect 10477 33734 10533 33790
rect 10557 33734 10613 33790
rect 10637 33734 10693 33790
rect 10717 33734 10773 33790
rect 10797 33734 10853 33790
rect 10877 33734 10933 33790
rect 10957 33734 11013 33790
rect 11037 33734 11093 33790
rect 11117 33774 11161 33790
rect 11161 33774 11173 33790
rect 11197 33774 11227 33790
rect 11227 33774 11253 33790
rect 11117 33760 11173 33774
rect 11197 33760 11253 33774
rect 11117 33734 11161 33760
rect 11161 33734 11173 33760
rect 11197 33734 11227 33760
rect 11227 33734 11253 33760
rect 11277 33734 11333 33790
rect 11357 33734 11413 33790
rect 11437 33734 11493 33790
rect 11517 33734 11573 33790
rect 11597 33734 11653 33790
rect 11677 33734 11733 33790
rect 11758 33734 11814 33790
rect 11839 33734 11895 33790
rect 11920 33774 11945 33790
rect 11945 33774 11976 33790
rect 12001 33774 12011 33790
rect 12011 33774 12057 33790
rect 11920 33760 11976 33774
rect 12001 33760 12057 33774
rect 11920 33734 11945 33760
rect 11945 33734 11976 33760
rect 12001 33734 12011 33760
rect 12011 33734 12057 33760
rect 5216 33508 5257 33526
rect 5257 33508 5272 33526
rect 5299 33508 5309 33526
rect 5309 33508 5323 33526
rect 5323 33508 5355 33526
rect 5216 33493 5272 33508
rect 5299 33493 5355 33508
rect 5216 33470 5257 33493
rect 5257 33470 5272 33493
rect 5299 33470 5309 33493
rect 5309 33470 5323 33493
rect 5323 33470 5355 33493
rect 5382 33470 5438 33526
rect 5465 33470 5521 33526
rect 5548 33470 5604 33526
rect 5631 33470 5687 33526
rect 5714 33470 5770 33526
rect 5797 33470 5853 33526
rect 5880 33470 5936 33526
rect 5963 33470 6019 33526
rect 6046 33508 6093 33526
rect 6093 33508 6102 33526
rect 6129 33508 6145 33526
rect 6145 33508 6159 33526
rect 6159 33508 6185 33526
rect 6046 33493 6102 33508
rect 6129 33493 6185 33508
rect 6046 33470 6093 33493
rect 6093 33470 6102 33493
rect 6129 33470 6145 33493
rect 6145 33470 6159 33493
rect 6159 33470 6185 33493
rect 6211 33470 6267 33526
rect 6293 33470 6349 33526
rect 6375 33470 6431 33526
rect 6457 33470 6513 33526
rect 6539 33470 6595 33526
rect 6621 33470 6677 33526
rect 6703 33470 6759 33526
rect 6785 33470 6841 33526
rect 6867 33470 6923 33526
rect 6949 33508 6981 33526
rect 6981 33508 6995 33526
rect 6995 33508 7005 33526
rect 7031 33508 7047 33526
rect 7047 33508 7087 33526
rect 6949 33493 7005 33508
rect 7031 33493 7087 33508
rect 6949 33470 6981 33493
rect 6981 33470 6995 33493
rect 6995 33470 7005 33493
rect 7031 33470 7047 33493
rect 7047 33470 7087 33493
rect 7113 33470 7169 33526
rect 7195 33470 7251 33526
rect 8041 33558 8097 33614
rect 8124 33558 8180 33614
rect 8207 33558 8263 33614
rect 8290 33558 8346 33614
rect 8373 33558 8429 33614
rect 8456 33558 8512 33614
rect 8539 33558 8595 33614
rect 8622 33575 8653 33614
rect 8653 33575 8667 33614
rect 8667 33575 8678 33614
rect 8705 33575 8719 33614
rect 8719 33575 8761 33614
rect 8622 33560 8678 33575
rect 8705 33560 8761 33575
rect 8622 33558 8653 33560
rect 8653 33558 8667 33560
rect 8667 33558 8678 33560
rect 8705 33558 8719 33560
rect 8719 33558 8761 33560
rect 8788 33558 8844 33614
rect 8871 33558 8927 33614
rect 8954 33558 9010 33614
rect 9037 33558 9093 33614
rect 9120 33558 9176 33614
rect 9203 33558 9259 33614
rect 9286 33558 9342 33614
rect 9369 33558 9425 33614
rect 9452 33575 9489 33614
rect 9489 33575 9503 33614
rect 9503 33575 9508 33614
rect 9535 33575 9555 33614
rect 9555 33575 9591 33614
rect 9452 33560 9508 33575
rect 9535 33560 9591 33575
rect 9452 33558 9489 33560
rect 9489 33558 9503 33560
rect 9503 33558 9508 33560
rect 9535 33558 9555 33560
rect 9555 33558 9591 33560
rect 9618 33558 9674 33614
rect 9702 33558 9758 33614
rect 10202 33594 10258 33650
rect 10286 33642 10325 33650
rect 10325 33642 10339 33650
rect 10339 33642 10342 33650
rect 10397 33646 10453 33702
rect 10477 33646 10533 33702
rect 10557 33646 10613 33702
rect 10637 33646 10693 33702
rect 10717 33646 10773 33702
rect 10797 33646 10853 33702
rect 10877 33646 10933 33702
rect 10957 33646 11013 33702
rect 11037 33646 11093 33702
rect 11117 33694 11173 33702
rect 11197 33694 11253 33702
rect 11117 33646 11161 33694
rect 11161 33646 11173 33694
rect 11197 33646 11227 33694
rect 11227 33646 11253 33694
rect 11277 33646 11333 33702
rect 11357 33646 11413 33702
rect 11437 33646 11493 33702
rect 11517 33646 11573 33702
rect 11597 33646 11653 33702
rect 11677 33646 11733 33702
rect 11758 33646 11814 33702
rect 11839 33646 11895 33702
rect 11920 33694 11976 33702
rect 12001 33694 12057 33702
rect 11920 33646 11945 33694
rect 11945 33646 11976 33694
rect 12001 33646 12011 33694
rect 12011 33646 12057 33694
rect 10286 33627 10342 33642
rect 10286 33594 10325 33627
rect 10325 33594 10339 33627
rect 10339 33594 10342 33627
rect 7943 33479 7999 33535
rect 10397 33558 10453 33614
rect 10477 33558 10533 33614
rect 10557 33558 10613 33614
rect 10637 33558 10693 33614
rect 10717 33558 10773 33614
rect 10797 33558 10853 33614
rect 10877 33558 10933 33614
rect 10957 33558 11013 33614
rect 11037 33558 11093 33614
rect 11117 33575 11161 33614
rect 11161 33575 11173 33614
rect 11197 33575 11227 33614
rect 11227 33575 11253 33614
rect 11117 33560 11173 33575
rect 11197 33560 11253 33575
rect 11117 33558 11161 33560
rect 11161 33558 11173 33560
rect 11197 33558 11227 33560
rect 11227 33558 11253 33560
rect 11277 33558 11333 33614
rect 11357 33558 11413 33614
rect 11437 33558 11493 33614
rect 11517 33558 11573 33614
rect 11597 33558 11653 33614
rect 11677 33558 11733 33614
rect 11758 33558 11814 33614
rect 11839 33558 11895 33614
rect 11920 33575 11945 33614
rect 11945 33575 11976 33614
rect 12001 33575 12011 33614
rect 12011 33575 12057 33614
rect 11920 33560 11976 33575
rect 12001 33560 12057 33575
rect 11920 33558 11945 33560
rect 11945 33558 11976 33560
rect 12001 33558 12011 33560
rect 12011 33558 12057 33560
rect 8041 33470 8097 33526
rect 8124 33470 8180 33526
rect 8207 33470 8263 33526
rect 8290 33470 8346 33526
rect 8373 33470 8429 33526
rect 8456 33470 8512 33526
rect 8539 33470 8595 33526
rect 8622 33508 8653 33526
rect 8653 33508 8667 33526
rect 8667 33508 8678 33526
rect 8705 33508 8719 33526
rect 8719 33508 8761 33526
rect 8622 33493 8678 33508
rect 8705 33493 8761 33508
rect 8622 33470 8653 33493
rect 8653 33470 8667 33493
rect 8667 33470 8678 33493
rect 8705 33470 8719 33493
rect 8719 33470 8761 33493
rect 8788 33470 8844 33526
rect 8871 33470 8927 33526
rect 8954 33470 9010 33526
rect 9037 33470 9093 33526
rect 9120 33470 9176 33526
rect 9203 33470 9259 33526
rect 9286 33470 9342 33526
rect 9369 33470 9425 33526
rect 9452 33508 9489 33526
rect 9489 33508 9503 33526
rect 9503 33508 9508 33526
rect 9535 33508 9555 33526
rect 9555 33508 9591 33526
rect 9452 33493 9508 33508
rect 9535 33493 9591 33508
rect 9452 33470 9489 33493
rect 9489 33470 9503 33493
rect 9503 33470 9508 33493
rect 9535 33470 9555 33493
rect 9555 33470 9591 33493
rect 9618 33470 9674 33526
rect 9702 33470 9758 33526
rect 10307 33508 10325 33535
rect 10325 33508 10339 33535
rect 10339 33508 10363 33535
rect 10307 33493 10363 33508
rect 10307 33479 10325 33493
rect 10325 33479 10339 33493
rect 10339 33479 10363 33493
rect 10397 33470 10453 33526
rect 10477 33470 10533 33526
rect 10557 33470 10613 33526
rect 10637 33470 10693 33526
rect 10717 33470 10773 33526
rect 10797 33470 10853 33526
rect 10877 33470 10933 33526
rect 10957 33470 11013 33526
rect 11037 33470 11093 33526
rect 11117 33508 11161 33526
rect 11161 33508 11173 33526
rect 11197 33508 11227 33526
rect 11227 33508 11253 33526
rect 11117 33493 11173 33508
rect 11197 33493 11253 33508
rect 11117 33470 11161 33493
rect 11161 33470 11173 33493
rect 11197 33470 11227 33493
rect 11227 33470 11253 33493
rect 11277 33470 11333 33526
rect 11357 33470 11413 33526
rect 11437 33470 11493 33526
rect 11517 33470 11573 33526
rect 11597 33470 11653 33526
rect 11677 33470 11733 33526
rect 11758 33470 11814 33526
rect 11839 33470 11895 33526
rect 11920 33508 11945 33526
rect 11945 33508 11976 33526
rect 12001 33508 12011 33526
rect 12011 33508 12057 33526
rect 11920 33493 11976 33508
rect 12001 33493 12057 33508
rect 11920 33470 11945 33493
rect 11945 33470 11976 33493
rect 12001 33470 12011 33493
rect 12011 33470 12057 33493
rect 5216 33426 5272 33438
rect 5299 33426 5355 33438
rect 3513 33370 3569 33426
rect 3594 33374 3637 33426
rect 3637 33374 3650 33426
rect 3675 33374 3703 33426
rect 3703 33374 3731 33426
rect 3594 33370 3650 33374
rect 3675 33370 3731 33374
rect 3757 33370 3813 33426
rect 3839 33370 3895 33426
rect 3921 33370 3977 33426
rect 4003 33370 4059 33426
rect 4085 33370 4141 33426
rect 4167 33370 4223 33426
rect 4249 33370 4305 33426
rect 5216 33382 5257 33426
rect 5257 33382 5272 33426
rect 5299 33382 5309 33426
rect 5309 33382 5323 33426
rect 5323 33382 5355 33426
rect 5382 33382 5438 33438
rect 5465 33382 5521 33438
rect 5548 33382 5604 33438
rect 5631 33382 5687 33438
rect 5714 33382 5770 33438
rect 5797 33382 5853 33438
rect 5880 33382 5936 33438
rect 5963 33382 6019 33438
rect 6046 33426 6102 33438
rect 6129 33426 6185 33438
rect 6046 33382 6093 33426
rect 6093 33382 6102 33426
rect 6129 33382 6145 33426
rect 6145 33382 6159 33426
rect 6159 33382 6185 33426
rect 6211 33382 6267 33438
rect 6293 33382 6349 33438
rect 6375 33382 6431 33438
rect 6457 33382 6513 33438
rect 6539 33382 6595 33438
rect 6621 33382 6677 33438
rect 6703 33382 6759 33438
rect 6785 33382 6841 33438
rect 6867 33382 6923 33438
rect 6949 33426 7005 33438
rect 7031 33426 7087 33438
rect 6949 33382 6981 33426
rect 6981 33382 6995 33426
rect 6995 33382 7005 33426
rect 7031 33382 7047 33426
rect 7047 33382 7087 33426
rect 7113 33382 7169 33438
rect 7195 33382 7251 33438
rect 8041 33382 8097 33438
rect 8124 33382 8180 33438
rect 8207 33382 8263 33438
rect 8290 33382 8346 33438
rect 8373 33382 8429 33438
rect 8456 33382 8512 33438
rect 8539 33382 8595 33438
rect 8622 33426 8678 33438
rect 8705 33426 8761 33438
rect 8622 33382 8653 33426
rect 8653 33382 8667 33426
rect 8667 33382 8678 33426
rect 8705 33382 8719 33426
rect 8719 33382 8761 33426
rect 8788 33382 8844 33438
rect 8871 33382 8927 33438
rect 8954 33382 9010 33438
rect 9037 33382 9093 33438
rect 9120 33382 9176 33438
rect 9203 33382 9259 33438
rect 9286 33382 9342 33438
rect 9369 33382 9425 33438
rect 9452 33426 9508 33438
rect 9535 33426 9591 33438
rect 9452 33382 9489 33426
rect 9489 33382 9503 33426
rect 9503 33382 9508 33426
rect 9535 33382 9555 33426
rect 9555 33382 9591 33426
rect 9618 33382 9674 33438
rect 9702 33382 9758 33438
rect 10397 33382 10453 33438
rect 10477 33382 10533 33438
rect 10557 33382 10613 33438
rect 10637 33382 10693 33438
rect 10717 33382 10773 33438
rect 10797 33382 10853 33438
rect 10877 33382 10933 33438
rect 10957 33382 11013 33438
rect 11037 33382 11093 33438
rect 11117 33426 11173 33438
rect 11197 33426 11253 33438
rect 11117 33382 11161 33426
rect 11161 33382 11173 33426
rect 11197 33382 11227 33426
rect 11227 33382 11253 33426
rect 11277 33382 11333 33438
rect 11357 33382 11413 33438
rect 11437 33382 11493 33438
rect 11517 33382 11573 33438
rect 11597 33382 11653 33438
rect 11677 33382 11733 33438
rect 11758 33382 11814 33438
rect 11839 33382 11895 33438
rect 11920 33426 11976 33438
rect 12001 33426 12057 33438
rect 11920 33382 11945 33426
rect 11945 33382 11976 33426
rect 12001 33382 12011 33426
rect 12011 33382 12057 33426
rect 3513 31840 3569 31896
rect 3596 31892 3652 31896
rect 3679 31892 3735 31896
rect 3596 31840 3637 31892
rect 3637 31840 3651 31892
rect 3651 31840 3652 31892
rect 3679 31840 3703 31892
rect 3703 31840 3735 31892
rect 3762 31840 3818 31896
rect 3845 31840 3901 31896
rect 3928 31840 3984 31896
rect 4011 31840 4067 31896
rect 4094 31840 4150 31896
rect 4177 31840 4233 31896
rect 4260 31840 4316 31896
rect 5215 31840 5257 31883
rect 5257 31840 5271 31883
rect 5296 31840 5309 31883
rect 5309 31840 5323 31883
rect 5323 31840 5352 31883
rect 5215 31827 5271 31840
rect 5296 31827 5352 31840
rect 5377 31827 5433 31883
rect 5458 31827 5514 31883
rect 5539 31827 5595 31883
rect 5620 31827 5676 31883
rect 5701 31827 5757 31883
rect 5782 31827 5838 31883
rect 5863 31827 5919 31883
rect 5944 31827 6000 31883
rect 6025 31827 6081 31883
rect 6106 31840 6145 31883
rect 6145 31840 6159 31883
rect 6159 31840 6162 31883
rect 6186 31840 6211 31883
rect 6211 31840 6242 31883
rect 6106 31827 6162 31840
rect 6186 31827 6242 31840
rect 6266 31827 6322 31883
rect 6346 31827 6402 31883
rect 8572 31840 8601 31883
rect 8601 31840 8628 31883
rect 8652 31840 8653 31883
rect 8653 31840 8667 31883
rect 8667 31840 8708 31883
rect 8572 31827 8628 31840
rect 8652 31827 8708 31840
rect 8732 31827 8788 31883
rect 8812 31827 8868 31883
rect 8893 31827 8949 31883
rect 8974 31827 9030 31883
rect 9055 31827 9111 31883
rect 9136 31827 9192 31883
rect 9217 31827 9273 31883
rect 9298 31827 9354 31883
rect 9379 31827 9435 31883
rect 9460 31840 9489 31883
rect 9489 31840 9503 31883
rect 9503 31840 9516 31883
rect 9541 31840 9555 31883
rect 9555 31840 9597 31883
rect 9460 31827 9516 31840
rect 9541 31827 9597 31840
rect 9622 31827 9678 31883
rect 9703 31827 9759 31883
rect 10871 31827 10927 31883
rect 10951 31827 11007 31883
rect 11031 31827 11087 31883
rect 11111 31840 11161 31883
rect 11161 31840 11167 31883
rect 11192 31840 11227 31883
rect 11227 31840 11248 31883
rect 11111 31827 11167 31840
rect 11192 31827 11248 31840
rect 11273 31827 11329 31883
rect 11354 31827 11410 31883
rect 11435 31827 11491 31883
rect 11516 31827 11572 31883
rect 11597 31827 11653 31883
rect 11678 31827 11734 31883
rect 11759 31827 11815 31883
rect 11840 31827 11896 31883
rect 11921 31840 11945 31883
rect 11945 31840 11977 31883
rect 12002 31840 12011 31883
rect 12011 31840 12058 31883
rect 11921 31827 11977 31840
rect 12002 31827 12058 31840
rect 3513 31746 3569 31802
rect 3596 31774 3637 31802
rect 3637 31774 3651 31802
rect 3651 31774 3652 31802
rect 3679 31774 3703 31802
rect 3703 31774 3735 31802
rect 3596 31760 3652 31774
rect 3679 31760 3735 31774
rect 3596 31746 3637 31760
rect 3637 31746 3651 31760
rect 3651 31746 3652 31760
rect 3679 31746 3703 31760
rect 3703 31746 3735 31760
rect 3762 31746 3818 31802
rect 3845 31746 3901 31802
rect 3928 31746 3984 31802
rect 4011 31746 4067 31802
rect 4094 31746 4150 31802
rect 4177 31746 4233 31802
rect 4260 31746 4316 31802
rect 5215 31774 5257 31795
rect 5257 31774 5271 31795
rect 5296 31774 5309 31795
rect 5309 31774 5323 31795
rect 5323 31774 5352 31795
rect 5215 31760 5271 31774
rect 5296 31760 5352 31774
rect 5215 31739 5257 31760
rect 5257 31739 5271 31760
rect 5296 31739 5309 31760
rect 5309 31739 5323 31760
rect 5323 31739 5352 31760
rect 5377 31739 5433 31795
rect 5458 31739 5514 31795
rect 5539 31739 5595 31795
rect 5620 31739 5676 31795
rect 5701 31739 5757 31795
rect 5782 31739 5838 31795
rect 5863 31739 5919 31795
rect 5944 31739 6000 31795
rect 6025 31739 6081 31795
rect 6106 31774 6145 31795
rect 6145 31774 6159 31795
rect 6159 31774 6162 31795
rect 6186 31774 6211 31795
rect 6211 31774 6242 31795
rect 6106 31760 6162 31774
rect 6186 31760 6242 31774
rect 6106 31739 6145 31760
rect 6145 31739 6159 31760
rect 6159 31739 6162 31760
rect 6186 31739 6211 31760
rect 6211 31739 6242 31760
rect 6266 31739 6322 31795
rect 6346 31739 6402 31795
rect 8572 31774 8601 31795
rect 8601 31774 8628 31795
rect 8652 31774 8653 31795
rect 8653 31774 8667 31795
rect 8667 31774 8708 31795
rect 8572 31760 8628 31774
rect 8652 31760 8708 31774
rect 8572 31739 8601 31760
rect 8601 31739 8628 31760
rect 8652 31739 8653 31760
rect 8653 31739 8667 31760
rect 8667 31739 8708 31760
rect 8732 31739 8788 31795
rect 8812 31739 8868 31795
rect 8893 31739 8949 31795
rect 8974 31739 9030 31795
rect 9055 31739 9111 31795
rect 9136 31739 9192 31795
rect 9217 31739 9273 31795
rect 9298 31739 9354 31795
rect 9379 31739 9435 31795
rect 9460 31774 9489 31795
rect 9489 31774 9503 31795
rect 9503 31774 9516 31795
rect 9541 31774 9555 31795
rect 9555 31774 9597 31795
rect 9460 31760 9516 31774
rect 9541 31760 9597 31774
rect 9460 31739 9489 31760
rect 9489 31739 9503 31760
rect 9503 31739 9516 31760
rect 9541 31739 9555 31760
rect 9555 31739 9597 31760
rect 9622 31739 9678 31795
rect 9703 31739 9759 31795
rect 10871 31739 10927 31795
rect 10951 31739 11007 31795
rect 11031 31739 11087 31795
rect 11111 31774 11161 31795
rect 11161 31774 11167 31795
rect 11192 31774 11227 31795
rect 11227 31774 11248 31795
rect 11111 31760 11167 31774
rect 11192 31760 11248 31774
rect 11111 31739 11161 31760
rect 11161 31739 11167 31760
rect 11192 31739 11227 31760
rect 11227 31739 11248 31760
rect 11273 31739 11329 31795
rect 11354 31739 11410 31795
rect 11435 31739 11491 31795
rect 11516 31739 11572 31795
rect 11597 31739 11653 31795
rect 11678 31739 11734 31795
rect 11759 31739 11815 31795
rect 11840 31739 11896 31795
rect 11921 31774 11945 31795
rect 11945 31774 11977 31795
rect 12002 31774 12011 31795
rect 12011 31774 12058 31795
rect 11921 31760 11977 31774
rect 12002 31760 12058 31774
rect 11921 31739 11945 31760
rect 11945 31739 11977 31760
rect 12002 31739 12011 31760
rect 12011 31739 12058 31760
rect 3513 31652 3569 31708
rect 3596 31694 3652 31708
rect 3679 31694 3735 31708
rect 3596 31652 3637 31694
rect 3637 31652 3651 31694
rect 3651 31652 3652 31694
rect 3679 31652 3703 31694
rect 3703 31652 3735 31694
rect 3762 31652 3818 31708
rect 3845 31652 3901 31708
rect 3928 31652 3984 31708
rect 4011 31652 4067 31708
rect 4094 31652 4150 31708
rect 4177 31652 4233 31708
rect 4260 31652 4316 31708
rect 5215 31694 5271 31707
rect 5296 31694 5352 31707
rect 5215 31651 5257 31694
rect 5257 31651 5271 31694
rect 5296 31651 5309 31694
rect 5309 31651 5323 31694
rect 5323 31651 5352 31694
rect 5377 31651 5433 31707
rect 5458 31651 5514 31707
rect 5539 31651 5595 31707
rect 5620 31651 5676 31707
rect 5701 31651 5757 31707
rect 5782 31651 5838 31707
rect 5863 31651 5919 31707
rect 5944 31651 6000 31707
rect 6025 31651 6081 31707
rect 6106 31694 6162 31707
rect 6186 31694 6242 31707
rect 6106 31651 6145 31694
rect 6145 31651 6159 31694
rect 6159 31651 6162 31694
rect 6186 31651 6211 31694
rect 6211 31651 6242 31694
rect 6266 31651 6322 31707
rect 6346 31651 6402 31707
rect 8572 31694 8628 31707
rect 8652 31694 8708 31707
rect 8572 31651 8601 31694
rect 8601 31651 8628 31694
rect 8652 31651 8653 31694
rect 8653 31651 8667 31694
rect 8667 31651 8708 31694
rect 8732 31651 8788 31707
rect 8812 31651 8868 31707
rect 8893 31651 8949 31707
rect 8974 31651 9030 31707
rect 9055 31651 9111 31707
rect 9136 31651 9192 31707
rect 9217 31651 9273 31707
rect 9298 31651 9354 31707
rect 9379 31651 9435 31707
rect 9460 31694 9516 31707
rect 9541 31694 9597 31707
rect 9460 31651 9489 31694
rect 9489 31651 9503 31694
rect 9503 31651 9516 31694
rect 9541 31651 9555 31694
rect 9555 31651 9597 31694
rect 9622 31651 9678 31707
rect 9703 31651 9759 31707
rect 10871 31651 10927 31707
rect 10951 31651 11007 31707
rect 11031 31651 11087 31707
rect 11111 31694 11167 31707
rect 11192 31694 11248 31707
rect 11111 31651 11161 31694
rect 11161 31651 11167 31694
rect 11192 31651 11227 31694
rect 11227 31651 11248 31694
rect 11273 31651 11329 31707
rect 11354 31651 11410 31707
rect 11435 31651 11491 31707
rect 11516 31651 11572 31707
rect 11597 31651 11653 31707
rect 11678 31651 11734 31707
rect 11759 31651 11815 31707
rect 11840 31651 11896 31707
rect 11921 31694 11977 31707
rect 12002 31694 12058 31707
rect 11921 31651 11945 31694
rect 11945 31651 11977 31694
rect 12002 31651 12011 31694
rect 12011 31651 12058 31694
rect 3513 31558 3569 31614
rect 3596 31575 3637 31614
rect 3637 31575 3651 31614
rect 3651 31575 3652 31614
rect 3679 31575 3703 31614
rect 3703 31575 3735 31614
rect 3596 31560 3652 31575
rect 3679 31560 3735 31575
rect 3596 31558 3637 31560
rect 3637 31558 3651 31560
rect 3651 31558 3652 31560
rect 3679 31558 3703 31560
rect 3703 31558 3735 31560
rect 3762 31558 3818 31614
rect 3845 31558 3901 31614
rect 3928 31558 3984 31614
rect 4011 31558 4067 31614
rect 4094 31558 4150 31614
rect 4177 31558 4233 31614
rect 4260 31558 4316 31614
rect 5215 31575 5257 31619
rect 5257 31575 5271 31619
rect 5296 31575 5309 31619
rect 5309 31575 5323 31619
rect 5323 31575 5352 31619
rect 5215 31563 5271 31575
rect 5296 31563 5352 31575
rect 5377 31563 5433 31619
rect 5458 31563 5514 31619
rect 5539 31563 5595 31619
rect 5620 31563 5676 31619
rect 5701 31563 5757 31619
rect 5782 31563 5838 31619
rect 5863 31563 5919 31619
rect 5944 31563 6000 31619
rect 6025 31563 6081 31619
rect 6106 31575 6145 31619
rect 6145 31575 6159 31619
rect 6159 31575 6162 31619
rect 6186 31575 6211 31619
rect 6211 31575 6242 31619
rect 6106 31563 6162 31575
rect 6186 31563 6242 31575
rect 6266 31563 6322 31619
rect 6346 31563 6402 31619
rect 8572 31575 8601 31619
rect 8601 31575 8628 31619
rect 8652 31575 8653 31619
rect 8653 31575 8667 31619
rect 8667 31575 8708 31619
rect 8572 31563 8628 31575
rect 8652 31563 8708 31575
rect 8732 31563 8788 31619
rect 8812 31563 8868 31619
rect 8893 31563 8949 31619
rect 8974 31563 9030 31619
rect 9055 31563 9111 31619
rect 9136 31563 9192 31619
rect 9217 31563 9273 31619
rect 9298 31563 9354 31619
rect 9379 31563 9435 31619
rect 9460 31575 9489 31619
rect 9489 31575 9503 31619
rect 9503 31575 9516 31619
rect 9541 31575 9555 31619
rect 9555 31575 9597 31619
rect 9460 31563 9516 31575
rect 9541 31563 9597 31575
rect 9622 31563 9678 31619
rect 9703 31563 9759 31619
rect 10871 31563 10927 31619
rect 10951 31563 11007 31619
rect 11031 31563 11087 31619
rect 11111 31575 11161 31619
rect 11161 31575 11167 31619
rect 11192 31575 11227 31619
rect 11227 31575 11248 31619
rect 11111 31563 11167 31575
rect 11192 31563 11248 31575
rect 11273 31563 11329 31619
rect 11354 31563 11410 31619
rect 11435 31563 11491 31619
rect 11516 31563 11572 31619
rect 11597 31563 11653 31619
rect 11678 31563 11734 31619
rect 11759 31563 11815 31619
rect 11840 31563 11896 31619
rect 11921 31575 11945 31619
rect 11945 31575 11977 31619
rect 12002 31575 12011 31619
rect 12011 31575 12058 31619
rect 11921 31563 11977 31575
rect 12002 31563 12058 31575
rect 3513 31464 3569 31520
rect 3596 31508 3637 31520
rect 3637 31508 3651 31520
rect 3651 31508 3652 31520
rect 3679 31508 3703 31520
rect 3703 31508 3735 31520
rect 3596 31493 3652 31508
rect 3679 31493 3735 31508
rect 3596 31464 3637 31493
rect 3637 31464 3651 31493
rect 3651 31464 3652 31493
rect 3679 31464 3703 31493
rect 3703 31464 3735 31493
rect 3762 31464 3818 31520
rect 3845 31464 3901 31520
rect 3928 31464 3984 31520
rect 4011 31464 4067 31520
rect 4094 31464 4150 31520
rect 4177 31464 4233 31520
rect 4260 31464 4316 31520
rect 5215 31508 5257 31531
rect 5257 31508 5271 31531
rect 5296 31508 5309 31531
rect 5309 31508 5323 31531
rect 5323 31508 5352 31531
rect 5215 31493 5271 31508
rect 5296 31493 5352 31508
rect 5215 31475 5257 31493
rect 5257 31475 5271 31493
rect 5296 31475 5309 31493
rect 5309 31475 5323 31493
rect 5323 31475 5352 31493
rect 5377 31475 5433 31531
rect 5458 31475 5514 31531
rect 5539 31475 5595 31531
rect 5620 31475 5676 31531
rect 5701 31475 5757 31531
rect 5782 31475 5838 31531
rect 5863 31475 5919 31531
rect 5944 31475 6000 31531
rect 6025 31475 6081 31531
rect 6106 31508 6145 31531
rect 6145 31508 6159 31531
rect 6159 31508 6162 31531
rect 6186 31508 6211 31531
rect 6211 31508 6242 31531
rect 6106 31493 6162 31508
rect 6186 31493 6242 31508
rect 6106 31475 6145 31493
rect 6145 31475 6159 31493
rect 6159 31475 6162 31493
rect 6186 31475 6211 31493
rect 6211 31475 6242 31493
rect 6266 31475 6322 31531
rect 6346 31475 6402 31531
rect 8572 31508 8601 31531
rect 8601 31508 8628 31531
rect 8652 31508 8653 31531
rect 8653 31508 8667 31531
rect 8667 31508 8708 31531
rect 8572 31493 8628 31508
rect 8652 31493 8708 31508
rect 5215 31441 5257 31443
rect 5257 31441 5271 31443
rect 5296 31441 5309 31443
rect 5309 31441 5323 31443
rect 5323 31441 5352 31443
rect 5215 31426 5271 31441
rect 5296 31426 5352 31441
rect 3513 31370 3569 31426
rect 3596 31374 3637 31426
rect 3637 31374 3651 31426
rect 3651 31374 3652 31426
rect 3679 31374 3703 31426
rect 3703 31374 3735 31426
rect 3596 31370 3652 31374
rect 3679 31370 3735 31374
rect 3762 31370 3818 31426
rect 3845 31370 3901 31426
rect 3928 31370 3984 31426
rect 4011 31370 4067 31426
rect 4094 31370 4150 31426
rect 4177 31370 4233 31426
rect 4260 31370 4316 31426
rect 5215 31387 5257 31426
rect 5257 31387 5271 31426
rect 5296 31387 5309 31426
rect 5309 31387 5323 31426
rect 5323 31387 5352 31426
rect 5377 31387 5433 31443
rect 5458 31387 5514 31443
rect 5539 31387 5595 31443
rect 5620 31387 5676 31443
rect 5701 31387 5757 31443
rect 5782 31387 5838 31443
rect 5863 31387 5919 31443
rect 5944 31387 6000 31443
rect 6025 31387 6081 31443
rect 6106 31441 6145 31443
rect 6145 31441 6159 31443
rect 6159 31441 6162 31443
rect 6186 31441 6211 31443
rect 6211 31441 6242 31443
rect 6106 31426 6162 31441
rect 6186 31426 6242 31441
rect 6106 31387 6145 31426
rect 6145 31387 6159 31426
rect 6159 31387 6162 31426
rect 6186 31387 6211 31426
rect 6211 31387 6242 31426
rect 6266 31387 6322 31443
rect 6346 31387 6402 31443
rect 8572 31475 8601 31493
rect 8601 31475 8628 31493
rect 8652 31475 8653 31493
rect 8653 31475 8667 31493
rect 8667 31475 8708 31493
rect 8732 31475 8788 31531
rect 8812 31475 8868 31531
rect 8893 31475 8949 31531
rect 8974 31475 9030 31531
rect 9055 31475 9111 31531
rect 9136 31475 9192 31531
rect 9217 31475 9273 31531
rect 9298 31475 9354 31531
rect 9379 31475 9435 31531
rect 9460 31508 9489 31531
rect 9489 31508 9503 31531
rect 9503 31508 9516 31531
rect 9541 31508 9555 31531
rect 9555 31508 9597 31531
rect 9460 31493 9516 31508
rect 9541 31493 9597 31508
rect 9460 31475 9489 31493
rect 9489 31475 9503 31493
rect 9503 31475 9516 31493
rect 9541 31475 9555 31493
rect 9555 31475 9597 31493
rect 9622 31475 9678 31531
rect 9703 31475 9759 31531
rect 8572 31441 8601 31443
rect 8601 31441 8628 31443
rect 8652 31441 8653 31443
rect 8653 31441 8667 31443
rect 8667 31441 8708 31443
rect 8572 31426 8628 31441
rect 8652 31426 8708 31441
rect 8572 31387 8601 31426
rect 8601 31387 8628 31426
rect 8652 31387 8653 31426
rect 8653 31387 8667 31426
rect 8667 31387 8708 31426
rect 8732 31387 8788 31443
rect 8812 31387 8868 31443
rect 8893 31387 8949 31443
rect 8974 31387 9030 31443
rect 9055 31387 9111 31443
rect 9136 31387 9192 31443
rect 9217 31387 9273 31443
rect 9298 31387 9354 31443
rect 9379 31387 9435 31443
rect 9460 31441 9489 31443
rect 9489 31441 9503 31443
rect 9503 31441 9516 31443
rect 9541 31441 9555 31443
rect 9555 31441 9597 31443
rect 9460 31426 9516 31441
rect 9541 31426 9597 31441
rect 9460 31387 9489 31426
rect 9489 31387 9503 31426
rect 9503 31387 9516 31426
rect 9541 31387 9555 31426
rect 9555 31387 9597 31426
rect 9622 31387 9678 31443
rect 9703 31387 9759 31443
rect 10871 31475 10927 31531
rect 10951 31475 11007 31531
rect 11031 31475 11087 31531
rect 11111 31508 11161 31531
rect 11161 31508 11167 31531
rect 11192 31508 11227 31531
rect 11227 31508 11248 31531
rect 11111 31493 11167 31508
rect 11192 31493 11248 31508
rect 11111 31475 11161 31493
rect 11161 31475 11167 31493
rect 11192 31475 11227 31493
rect 11227 31475 11248 31493
rect 11273 31475 11329 31531
rect 11354 31475 11410 31531
rect 11435 31475 11491 31531
rect 11516 31475 11572 31531
rect 11597 31475 11653 31531
rect 11678 31475 11734 31531
rect 11759 31475 11815 31531
rect 11840 31475 11896 31531
rect 11921 31508 11945 31531
rect 11945 31508 11977 31531
rect 12002 31508 12011 31531
rect 12011 31508 12058 31531
rect 11921 31493 11977 31508
rect 12002 31493 12058 31508
rect 11921 31475 11945 31493
rect 11945 31475 11977 31493
rect 12002 31475 12011 31493
rect 12011 31475 12058 31493
rect 10871 31387 10927 31443
rect 10951 31387 11007 31443
rect 11031 31387 11087 31443
rect 11111 31441 11161 31443
rect 11161 31441 11167 31443
rect 11192 31441 11227 31443
rect 11227 31441 11248 31443
rect 11111 31426 11167 31441
rect 11192 31426 11248 31441
rect 11111 31387 11161 31426
rect 11161 31387 11167 31426
rect 11192 31387 11227 31426
rect 11227 31387 11248 31426
rect 11273 31387 11329 31443
rect 11354 31387 11410 31443
rect 11435 31387 11491 31443
rect 11516 31387 11572 31443
rect 11597 31387 11653 31443
rect 11678 31387 11734 31443
rect 11759 31387 11815 31443
rect 11840 31387 11896 31443
rect 11921 31441 11945 31443
rect 11945 31441 11977 31443
rect 12002 31441 12011 31443
rect 12011 31441 12058 31443
rect 11921 31426 11977 31441
rect 12002 31426 12058 31441
rect 11921 31387 11945 31426
rect 11945 31387 11977 31426
rect 12002 31387 12011 31426
rect 12011 31387 12058 31426
rect 3513 29840 3569 29896
rect 3596 29892 3652 29896
rect 3679 29892 3735 29896
rect 3596 29840 3637 29892
rect 3637 29840 3651 29892
rect 3651 29840 3652 29892
rect 3679 29840 3703 29892
rect 3703 29840 3735 29892
rect 3762 29840 3818 29896
rect 3845 29840 3901 29896
rect 3928 29840 3984 29896
rect 4011 29840 4067 29896
rect 4094 29840 4150 29896
rect 4177 29840 4233 29896
rect 4260 29840 4316 29896
rect 5215 29840 5257 29883
rect 5257 29840 5271 29883
rect 5296 29840 5309 29883
rect 5309 29840 5323 29883
rect 5323 29840 5352 29883
rect 5215 29827 5271 29840
rect 5296 29827 5352 29840
rect 5377 29827 5433 29883
rect 5458 29827 5514 29883
rect 5539 29827 5595 29883
rect 5620 29827 5676 29883
rect 5701 29827 5757 29883
rect 5782 29827 5838 29883
rect 5863 29827 5919 29883
rect 5944 29827 6000 29883
rect 6025 29827 6081 29883
rect 6106 29840 6145 29883
rect 6145 29840 6159 29883
rect 6159 29840 6162 29883
rect 6186 29840 6211 29883
rect 6211 29840 6242 29883
rect 6106 29827 6162 29840
rect 6186 29827 6242 29840
rect 6266 29827 6322 29883
rect 6346 29827 6402 29883
rect 8572 29840 8601 29883
rect 8601 29840 8628 29883
rect 8652 29840 8653 29883
rect 8653 29840 8667 29883
rect 8667 29840 8708 29883
rect 8572 29827 8628 29840
rect 8652 29827 8708 29840
rect 8732 29827 8788 29883
rect 8812 29827 8868 29883
rect 8893 29827 8949 29883
rect 8974 29827 9030 29883
rect 9055 29827 9111 29883
rect 9136 29827 9192 29883
rect 9217 29827 9273 29883
rect 9298 29827 9354 29883
rect 9379 29827 9435 29883
rect 9460 29840 9489 29883
rect 9489 29840 9503 29883
rect 9503 29840 9516 29883
rect 9541 29840 9555 29883
rect 9555 29840 9597 29883
rect 9460 29827 9516 29840
rect 9541 29827 9597 29840
rect 9622 29827 9678 29883
rect 9703 29827 9759 29883
rect 10871 29827 10927 29883
rect 10951 29827 11007 29883
rect 11031 29827 11087 29883
rect 11111 29840 11161 29883
rect 11161 29840 11167 29883
rect 11192 29840 11227 29883
rect 11227 29840 11248 29883
rect 11111 29827 11167 29840
rect 11192 29827 11248 29840
rect 11273 29827 11329 29883
rect 11354 29827 11410 29883
rect 11435 29827 11491 29883
rect 11516 29827 11572 29883
rect 11597 29827 11653 29883
rect 11678 29827 11734 29883
rect 11759 29827 11815 29883
rect 11840 29827 11896 29883
rect 11921 29840 11945 29883
rect 11945 29840 11977 29883
rect 12002 29840 12011 29883
rect 12011 29840 12058 29883
rect 11921 29827 11977 29840
rect 12002 29827 12058 29840
rect 3513 29746 3569 29802
rect 3596 29774 3637 29802
rect 3637 29774 3651 29802
rect 3651 29774 3652 29802
rect 3679 29774 3703 29802
rect 3703 29774 3735 29802
rect 3596 29760 3652 29774
rect 3679 29760 3735 29774
rect 3596 29746 3637 29760
rect 3637 29746 3651 29760
rect 3651 29746 3652 29760
rect 3679 29746 3703 29760
rect 3703 29746 3735 29760
rect 3762 29746 3818 29802
rect 3845 29746 3901 29802
rect 3928 29746 3984 29802
rect 4011 29746 4067 29802
rect 4094 29746 4150 29802
rect 4177 29746 4233 29802
rect 4260 29746 4316 29802
rect 5215 29774 5257 29795
rect 5257 29774 5271 29795
rect 5296 29774 5309 29795
rect 5309 29774 5323 29795
rect 5323 29774 5352 29795
rect 5215 29760 5271 29774
rect 5296 29760 5352 29774
rect 5215 29739 5257 29760
rect 5257 29739 5271 29760
rect 5296 29739 5309 29760
rect 5309 29739 5323 29760
rect 5323 29739 5352 29760
rect 5377 29739 5433 29795
rect 5458 29739 5514 29795
rect 5539 29739 5595 29795
rect 5620 29739 5676 29795
rect 5701 29739 5757 29795
rect 5782 29739 5838 29795
rect 5863 29739 5919 29795
rect 5944 29739 6000 29795
rect 6025 29739 6081 29795
rect 6106 29774 6145 29795
rect 6145 29774 6159 29795
rect 6159 29774 6162 29795
rect 6186 29774 6211 29795
rect 6211 29774 6242 29795
rect 6106 29760 6162 29774
rect 6186 29760 6242 29774
rect 6106 29739 6145 29760
rect 6145 29739 6159 29760
rect 6159 29739 6162 29760
rect 6186 29739 6211 29760
rect 6211 29739 6242 29760
rect 6266 29739 6322 29795
rect 6346 29739 6402 29795
rect 8572 29774 8601 29795
rect 8601 29774 8628 29795
rect 8652 29774 8653 29795
rect 8653 29774 8667 29795
rect 8667 29774 8708 29795
rect 8572 29760 8628 29774
rect 8652 29760 8708 29774
rect 8572 29739 8601 29760
rect 8601 29739 8628 29760
rect 8652 29739 8653 29760
rect 8653 29739 8667 29760
rect 8667 29739 8708 29760
rect 8732 29739 8788 29795
rect 8812 29739 8868 29795
rect 8893 29739 8949 29795
rect 8974 29739 9030 29795
rect 9055 29739 9111 29795
rect 9136 29739 9192 29795
rect 9217 29739 9273 29795
rect 9298 29739 9354 29795
rect 9379 29739 9435 29795
rect 9460 29774 9489 29795
rect 9489 29774 9503 29795
rect 9503 29774 9516 29795
rect 9541 29774 9555 29795
rect 9555 29774 9597 29795
rect 9460 29760 9516 29774
rect 9541 29760 9597 29774
rect 9460 29739 9489 29760
rect 9489 29739 9503 29760
rect 9503 29739 9516 29760
rect 9541 29739 9555 29760
rect 9555 29739 9597 29760
rect 9622 29739 9678 29795
rect 9703 29739 9759 29795
rect 10871 29739 10927 29795
rect 10951 29739 11007 29795
rect 11031 29739 11087 29795
rect 11111 29774 11161 29795
rect 11161 29774 11167 29795
rect 11192 29774 11227 29795
rect 11227 29774 11248 29795
rect 11111 29760 11167 29774
rect 11192 29760 11248 29774
rect 11111 29739 11161 29760
rect 11161 29739 11167 29760
rect 11192 29739 11227 29760
rect 11227 29739 11248 29760
rect 11273 29739 11329 29795
rect 11354 29739 11410 29795
rect 11435 29739 11491 29795
rect 11516 29739 11572 29795
rect 11597 29739 11653 29795
rect 11678 29739 11734 29795
rect 11759 29739 11815 29795
rect 11840 29739 11896 29795
rect 11921 29774 11945 29795
rect 11945 29774 11977 29795
rect 12002 29774 12011 29795
rect 12011 29774 12058 29795
rect 11921 29760 11977 29774
rect 12002 29760 12058 29774
rect 11921 29739 11945 29760
rect 11945 29739 11977 29760
rect 12002 29739 12011 29760
rect 12011 29739 12058 29760
rect 3513 29652 3569 29708
rect 3596 29694 3652 29708
rect 3679 29694 3735 29708
rect 3596 29652 3637 29694
rect 3637 29652 3651 29694
rect 3651 29652 3652 29694
rect 3679 29652 3703 29694
rect 3703 29652 3735 29694
rect 3762 29652 3818 29708
rect 3845 29652 3901 29708
rect 3928 29652 3984 29708
rect 4011 29652 4067 29708
rect 4094 29652 4150 29708
rect 4177 29652 4233 29708
rect 4260 29652 4316 29708
rect 5215 29694 5271 29707
rect 5296 29694 5352 29707
rect 5215 29651 5257 29694
rect 5257 29651 5271 29694
rect 5296 29651 5309 29694
rect 5309 29651 5323 29694
rect 5323 29651 5352 29694
rect 5377 29651 5433 29707
rect 5458 29651 5514 29707
rect 5539 29651 5595 29707
rect 5620 29651 5676 29707
rect 5701 29651 5757 29707
rect 5782 29651 5838 29707
rect 5863 29651 5919 29707
rect 5944 29651 6000 29707
rect 6025 29651 6081 29707
rect 6106 29694 6162 29707
rect 6186 29694 6242 29707
rect 6106 29651 6145 29694
rect 6145 29651 6159 29694
rect 6159 29651 6162 29694
rect 6186 29651 6211 29694
rect 6211 29651 6242 29694
rect 6266 29651 6322 29707
rect 6346 29651 6402 29707
rect 8572 29694 8628 29707
rect 8652 29694 8708 29707
rect 8572 29651 8601 29694
rect 8601 29651 8628 29694
rect 8652 29651 8653 29694
rect 8653 29651 8667 29694
rect 8667 29651 8708 29694
rect 8732 29651 8788 29707
rect 8812 29651 8868 29707
rect 8893 29651 8949 29707
rect 8974 29651 9030 29707
rect 9055 29651 9111 29707
rect 9136 29651 9192 29707
rect 9217 29651 9273 29707
rect 9298 29651 9354 29707
rect 9379 29651 9435 29707
rect 9460 29694 9516 29707
rect 9541 29694 9597 29707
rect 9460 29651 9489 29694
rect 9489 29651 9503 29694
rect 9503 29651 9516 29694
rect 9541 29651 9555 29694
rect 9555 29651 9597 29694
rect 9622 29651 9678 29707
rect 9703 29651 9759 29707
rect 10871 29651 10927 29707
rect 10951 29651 11007 29707
rect 11031 29651 11087 29707
rect 11111 29694 11167 29707
rect 11192 29694 11248 29707
rect 11111 29651 11161 29694
rect 11161 29651 11167 29694
rect 11192 29651 11227 29694
rect 11227 29651 11248 29694
rect 11273 29651 11329 29707
rect 11354 29651 11410 29707
rect 11435 29651 11491 29707
rect 11516 29651 11572 29707
rect 11597 29651 11653 29707
rect 11678 29651 11734 29707
rect 11759 29651 11815 29707
rect 11840 29651 11896 29707
rect 11921 29694 11977 29707
rect 12002 29694 12058 29707
rect 11921 29651 11945 29694
rect 11945 29651 11977 29694
rect 12002 29651 12011 29694
rect 12011 29651 12058 29694
rect 3513 29558 3569 29614
rect 3596 29575 3637 29614
rect 3637 29575 3651 29614
rect 3651 29575 3652 29614
rect 3679 29575 3703 29614
rect 3703 29575 3735 29614
rect 3596 29560 3652 29575
rect 3679 29560 3735 29575
rect 3596 29558 3637 29560
rect 3637 29558 3651 29560
rect 3651 29558 3652 29560
rect 3679 29558 3703 29560
rect 3703 29558 3735 29560
rect 3762 29558 3818 29614
rect 3845 29558 3901 29614
rect 3928 29558 3984 29614
rect 4011 29558 4067 29614
rect 4094 29558 4150 29614
rect 4177 29558 4233 29614
rect 4260 29558 4316 29614
rect 5215 29575 5257 29619
rect 5257 29575 5271 29619
rect 5296 29575 5309 29619
rect 5309 29575 5323 29619
rect 5323 29575 5352 29619
rect 5215 29563 5271 29575
rect 5296 29563 5352 29575
rect 5377 29563 5433 29619
rect 5458 29563 5514 29619
rect 5539 29563 5595 29619
rect 5620 29563 5676 29619
rect 5701 29563 5757 29619
rect 5782 29563 5838 29619
rect 5863 29563 5919 29619
rect 5944 29563 6000 29619
rect 6025 29563 6081 29619
rect 6106 29575 6145 29619
rect 6145 29575 6159 29619
rect 6159 29575 6162 29619
rect 6186 29575 6211 29619
rect 6211 29575 6242 29619
rect 6106 29563 6162 29575
rect 6186 29563 6242 29575
rect 6266 29563 6322 29619
rect 6346 29563 6402 29619
rect 8572 29575 8601 29619
rect 8601 29575 8628 29619
rect 8652 29575 8653 29619
rect 8653 29575 8667 29619
rect 8667 29575 8708 29619
rect 8572 29563 8628 29575
rect 8652 29563 8708 29575
rect 8732 29563 8788 29619
rect 8812 29563 8868 29619
rect 8893 29563 8949 29619
rect 8974 29563 9030 29619
rect 9055 29563 9111 29619
rect 9136 29563 9192 29619
rect 9217 29563 9273 29619
rect 9298 29563 9354 29619
rect 9379 29563 9435 29619
rect 9460 29575 9489 29619
rect 9489 29575 9503 29619
rect 9503 29575 9516 29619
rect 9541 29575 9555 29619
rect 9555 29575 9597 29619
rect 9460 29563 9516 29575
rect 9541 29563 9597 29575
rect 9622 29563 9678 29619
rect 9703 29563 9759 29619
rect 10871 29563 10927 29619
rect 10951 29563 11007 29619
rect 11031 29563 11087 29619
rect 11111 29575 11161 29619
rect 11161 29575 11167 29619
rect 11192 29575 11227 29619
rect 11227 29575 11248 29619
rect 11111 29563 11167 29575
rect 11192 29563 11248 29575
rect 11273 29563 11329 29619
rect 11354 29563 11410 29619
rect 11435 29563 11491 29619
rect 11516 29563 11572 29619
rect 11597 29563 11653 29619
rect 11678 29563 11734 29619
rect 11759 29563 11815 29619
rect 11840 29563 11896 29619
rect 11921 29575 11945 29619
rect 11945 29575 11977 29619
rect 12002 29575 12011 29619
rect 12011 29575 12058 29619
rect 11921 29563 11977 29575
rect 12002 29563 12058 29575
rect 3513 29464 3569 29520
rect 3596 29508 3637 29520
rect 3637 29508 3651 29520
rect 3651 29508 3652 29520
rect 3679 29508 3703 29520
rect 3703 29508 3735 29520
rect 3596 29493 3652 29508
rect 3679 29493 3735 29508
rect 3596 29464 3637 29493
rect 3637 29464 3651 29493
rect 3651 29464 3652 29493
rect 3679 29464 3703 29493
rect 3703 29464 3735 29493
rect 3762 29464 3818 29520
rect 3845 29464 3901 29520
rect 3928 29464 3984 29520
rect 4011 29464 4067 29520
rect 4094 29464 4150 29520
rect 4177 29464 4233 29520
rect 4260 29464 4316 29520
rect 5215 29508 5257 29531
rect 5257 29508 5271 29531
rect 5296 29508 5309 29531
rect 5309 29508 5323 29531
rect 5323 29508 5352 29531
rect 5215 29493 5271 29508
rect 5296 29493 5352 29508
rect 5215 29475 5257 29493
rect 5257 29475 5271 29493
rect 5296 29475 5309 29493
rect 5309 29475 5323 29493
rect 5323 29475 5352 29493
rect 5377 29475 5433 29531
rect 5458 29475 5514 29531
rect 5539 29475 5595 29531
rect 5620 29475 5676 29531
rect 5701 29475 5757 29531
rect 5782 29475 5838 29531
rect 5863 29475 5919 29531
rect 5944 29475 6000 29531
rect 6025 29475 6081 29531
rect 6106 29508 6145 29531
rect 6145 29508 6159 29531
rect 6159 29508 6162 29531
rect 6186 29508 6211 29531
rect 6211 29508 6242 29531
rect 6106 29493 6162 29508
rect 6186 29493 6242 29508
rect 6106 29475 6145 29493
rect 6145 29475 6159 29493
rect 6159 29475 6162 29493
rect 6186 29475 6211 29493
rect 6211 29475 6242 29493
rect 6266 29475 6322 29531
rect 6346 29475 6402 29531
rect 8572 29508 8601 29531
rect 8601 29508 8628 29531
rect 8652 29508 8653 29531
rect 8653 29508 8667 29531
rect 8667 29508 8708 29531
rect 8572 29493 8628 29508
rect 8652 29493 8708 29508
rect 5215 29441 5257 29443
rect 5257 29441 5271 29443
rect 5296 29441 5309 29443
rect 5309 29441 5323 29443
rect 5323 29441 5352 29443
rect 5215 29426 5271 29441
rect 5296 29426 5352 29441
rect 3513 29370 3569 29426
rect 3596 29374 3637 29426
rect 3637 29374 3651 29426
rect 3651 29374 3652 29426
rect 3679 29374 3703 29426
rect 3703 29374 3735 29426
rect 3596 29370 3652 29374
rect 3679 29370 3735 29374
rect 3762 29370 3818 29426
rect 3845 29370 3901 29426
rect 3928 29370 3984 29426
rect 4011 29370 4067 29426
rect 4094 29370 4150 29426
rect 4177 29370 4233 29426
rect 4260 29370 4316 29426
rect 5215 29387 5257 29426
rect 5257 29387 5271 29426
rect 5296 29387 5309 29426
rect 5309 29387 5323 29426
rect 5323 29387 5352 29426
rect 5377 29387 5433 29443
rect 5458 29387 5514 29443
rect 5539 29387 5595 29443
rect 5620 29387 5676 29443
rect 5701 29387 5757 29443
rect 5782 29387 5838 29443
rect 5863 29387 5919 29443
rect 5944 29387 6000 29443
rect 6025 29387 6081 29443
rect 6106 29441 6145 29443
rect 6145 29441 6159 29443
rect 6159 29441 6162 29443
rect 6186 29441 6211 29443
rect 6211 29441 6242 29443
rect 6106 29426 6162 29441
rect 6186 29426 6242 29441
rect 6106 29387 6145 29426
rect 6145 29387 6159 29426
rect 6159 29387 6162 29426
rect 6186 29387 6211 29426
rect 6211 29387 6242 29426
rect 6266 29387 6322 29443
rect 6346 29387 6402 29443
rect 8572 29475 8601 29493
rect 8601 29475 8628 29493
rect 8652 29475 8653 29493
rect 8653 29475 8667 29493
rect 8667 29475 8708 29493
rect 8732 29475 8788 29531
rect 8812 29475 8868 29531
rect 8893 29475 8949 29531
rect 8974 29475 9030 29531
rect 9055 29475 9111 29531
rect 9136 29475 9192 29531
rect 9217 29475 9273 29531
rect 9298 29475 9354 29531
rect 9379 29475 9435 29531
rect 9460 29508 9489 29531
rect 9489 29508 9503 29531
rect 9503 29508 9516 29531
rect 9541 29508 9555 29531
rect 9555 29508 9597 29531
rect 9460 29493 9516 29508
rect 9541 29493 9597 29508
rect 9460 29475 9489 29493
rect 9489 29475 9503 29493
rect 9503 29475 9516 29493
rect 9541 29475 9555 29493
rect 9555 29475 9597 29493
rect 9622 29475 9678 29531
rect 9703 29475 9759 29531
rect 8572 29441 8601 29443
rect 8601 29441 8628 29443
rect 8652 29441 8653 29443
rect 8653 29441 8667 29443
rect 8667 29441 8708 29443
rect 8572 29426 8628 29441
rect 8652 29426 8708 29441
rect 8572 29387 8601 29426
rect 8601 29387 8628 29426
rect 8652 29387 8653 29426
rect 8653 29387 8667 29426
rect 8667 29387 8708 29426
rect 8732 29387 8788 29443
rect 8812 29387 8868 29443
rect 8893 29387 8949 29443
rect 8974 29387 9030 29443
rect 9055 29387 9111 29443
rect 9136 29387 9192 29443
rect 9217 29387 9273 29443
rect 9298 29387 9354 29443
rect 9379 29387 9435 29443
rect 9460 29441 9489 29443
rect 9489 29441 9503 29443
rect 9503 29441 9516 29443
rect 9541 29441 9555 29443
rect 9555 29441 9597 29443
rect 9460 29426 9516 29441
rect 9541 29426 9597 29441
rect 9460 29387 9489 29426
rect 9489 29387 9503 29426
rect 9503 29387 9516 29426
rect 9541 29387 9555 29426
rect 9555 29387 9597 29426
rect 9622 29387 9678 29443
rect 9703 29387 9759 29443
rect 10871 29475 10927 29531
rect 10951 29475 11007 29531
rect 11031 29475 11087 29531
rect 11111 29508 11161 29531
rect 11161 29508 11167 29531
rect 11192 29508 11227 29531
rect 11227 29508 11248 29531
rect 11111 29493 11167 29508
rect 11192 29493 11248 29508
rect 11111 29475 11161 29493
rect 11161 29475 11167 29493
rect 11192 29475 11227 29493
rect 11227 29475 11248 29493
rect 11273 29475 11329 29531
rect 11354 29475 11410 29531
rect 11435 29475 11491 29531
rect 11516 29475 11572 29531
rect 11597 29475 11653 29531
rect 11678 29475 11734 29531
rect 11759 29475 11815 29531
rect 11840 29475 11896 29531
rect 11921 29508 11945 29531
rect 11945 29508 11977 29531
rect 12002 29508 12011 29531
rect 12011 29508 12058 29531
rect 11921 29493 11977 29508
rect 12002 29493 12058 29508
rect 11921 29475 11945 29493
rect 11945 29475 11977 29493
rect 12002 29475 12011 29493
rect 12011 29475 12058 29493
rect 10871 29387 10927 29443
rect 10951 29387 11007 29443
rect 11031 29387 11087 29443
rect 11111 29441 11161 29443
rect 11161 29441 11167 29443
rect 11192 29441 11227 29443
rect 11227 29441 11248 29443
rect 11111 29426 11167 29441
rect 11192 29426 11248 29441
rect 11111 29387 11161 29426
rect 11161 29387 11167 29426
rect 11192 29387 11227 29426
rect 11227 29387 11248 29426
rect 11273 29387 11329 29443
rect 11354 29387 11410 29443
rect 11435 29387 11491 29443
rect 11516 29387 11572 29443
rect 11597 29387 11653 29443
rect 11678 29387 11734 29443
rect 11759 29387 11815 29443
rect 11840 29387 11896 29443
rect 11921 29441 11945 29443
rect 11945 29441 11977 29443
rect 12002 29441 12011 29443
rect 12011 29441 12058 29443
rect 11921 29426 11977 29441
rect 12002 29426 12058 29441
rect 11921 29387 11945 29426
rect 11945 29387 11977 29426
rect 12002 29387 12011 29426
rect 12011 29387 12058 29426
rect 3452 27840 3508 27896
rect 3532 27840 3588 27896
rect 3612 27840 3668 27896
rect 3693 27840 3749 27896
rect 3774 27840 3830 27896
rect 3855 27840 3911 27896
rect 3936 27840 3992 27896
rect 4017 27840 4073 27896
rect 4098 27840 4154 27896
rect 4179 27840 4235 27896
rect 4260 27840 4316 27896
rect 5215 27840 5257 27883
rect 5257 27840 5271 27883
rect 5296 27840 5309 27883
rect 5309 27840 5323 27883
rect 5323 27840 5352 27883
rect 5215 27827 5271 27840
rect 5296 27827 5352 27840
rect 5377 27827 5433 27883
rect 5458 27827 5514 27883
rect 5539 27827 5595 27883
rect 5620 27827 5676 27883
rect 5701 27827 5757 27883
rect 5782 27827 5838 27883
rect 5863 27827 5919 27883
rect 5944 27827 6000 27883
rect 6025 27827 6081 27883
rect 6106 27840 6145 27883
rect 6145 27840 6159 27883
rect 6159 27840 6162 27883
rect 6186 27840 6211 27883
rect 6211 27840 6242 27883
rect 6106 27827 6162 27840
rect 6186 27827 6242 27840
rect 6266 27827 6322 27883
rect 6346 27827 6402 27883
rect 8572 27840 8601 27883
rect 8601 27840 8628 27883
rect 8652 27840 8653 27883
rect 8653 27840 8667 27883
rect 8667 27840 8708 27883
rect 8572 27827 8628 27840
rect 8652 27827 8708 27840
rect 8732 27827 8788 27883
rect 8812 27827 8868 27883
rect 8893 27827 8949 27883
rect 8974 27827 9030 27883
rect 9055 27827 9111 27883
rect 9136 27827 9192 27883
rect 9217 27827 9273 27883
rect 9298 27827 9354 27883
rect 9379 27827 9435 27883
rect 9460 27840 9489 27883
rect 9489 27840 9503 27883
rect 9503 27840 9516 27883
rect 9541 27840 9555 27883
rect 9555 27840 9597 27883
rect 9460 27827 9516 27840
rect 9541 27827 9597 27840
rect 9622 27827 9678 27883
rect 9703 27827 9759 27883
rect 10871 27827 10927 27883
rect 10951 27827 11007 27883
rect 11031 27827 11087 27883
rect 11111 27840 11161 27883
rect 11161 27840 11167 27883
rect 11192 27840 11227 27883
rect 11227 27840 11248 27883
rect 11111 27827 11167 27840
rect 11192 27827 11248 27840
rect 11273 27827 11329 27883
rect 11354 27827 11410 27883
rect 11435 27827 11491 27883
rect 11516 27827 11572 27883
rect 11597 27827 11653 27883
rect 11678 27827 11734 27883
rect 11759 27827 11815 27883
rect 11840 27827 11896 27883
rect 11921 27840 11945 27883
rect 11945 27840 11977 27883
rect 12002 27840 12011 27883
rect 12011 27840 12058 27883
rect 11921 27827 11977 27840
rect 12002 27827 12058 27840
rect 3452 27746 3508 27802
rect 3532 27746 3588 27802
rect 3612 27746 3668 27802
rect 3693 27746 3749 27802
rect 3774 27746 3830 27802
rect 3855 27746 3911 27802
rect 3936 27746 3992 27802
rect 4017 27746 4073 27802
rect 4098 27746 4154 27802
rect 4179 27746 4235 27802
rect 4260 27746 4316 27802
rect 5215 27774 5257 27795
rect 5257 27774 5271 27795
rect 5296 27774 5309 27795
rect 5309 27774 5323 27795
rect 5323 27774 5352 27795
rect 5215 27760 5271 27774
rect 5296 27760 5352 27774
rect 5215 27739 5257 27760
rect 5257 27739 5271 27760
rect 5296 27739 5309 27760
rect 5309 27739 5323 27760
rect 5323 27739 5352 27760
rect 5377 27739 5433 27795
rect 5458 27739 5514 27795
rect 5539 27739 5595 27795
rect 5620 27739 5676 27795
rect 5701 27739 5757 27795
rect 5782 27739 5838 27795
rect 5863 27739 5919 27795
rect 5944 27739 6000 27795
rect 6025 27739 6081 27795
rect 6106 27774 6145 27795
rect 6145 27774 6159 27795
rect 6159 27774 6162 27795
rect 6186 27774 6211 27795
rect 6211 27774 6242 27795
rect 6106 27760 6162 27774
rect 6186 27760 6242 27774
rect 6106 27739 6145 27760
rect 6145 27739 6159 27760
rect 6159 27739 6162 27760
rect 6186 27739 6211 27760
rect 6211 27739 6242 27760
rect 6266 27739 6322 27795
rect 6346 27739 6402 27795
rect 8572 27774 8601 27795
rect 8601 27774 8628 27795
rect 8652 27774 8653 27795
rect 8653 27774 8667 27795
rect 8667 27774 8708 27795
rect 8572 27760 8628 27774
rect 8652 27760 8708 27774
rect 8572 27739 8601 27760
rect 8601 27739 8628 27760
rect 8652 27739 8653 27760
rect 8653 27739 8667 27760
rect 8667 27739 8708 27760
rect 8732 27739 8788 27795
rect 8812 27739 8868 27795
rect 8893 27739 8949 27795
rect 8974 27739 9030 27795
rect 9055 27739 9111 27795
rect 9136 27739 9192 27795
rect 9217 27739 9273 27795
rect 9298 27739 9354 27795
rect 9379 27739 9435 27795
rect 9460 27774 9489 27795
rect 9489 27774 9503 27795
rect 9503 27774 9516 27795
rect 9541 27774 9555 27795
rect 9555 27774 9597 27795
rect 9460 27760 9516 27774
rect 9541 27760 9597 27774
rect 9460 27739 9489 27760
rect 9489 27739 9503 27760
rect 9503 27739 9516 27760
rect 9541 27739 9555 27760
rect 9555 27739 9597 27760
rect 9622 27739 9678 27795
rect 9703 27739 9759 27795
rect 10871 27739 10927 27795
rect 10951 27739 11007 27795
rect 11031 27739 11087 27795
rect 11111 27774 11161 27795
rect 11161 27774 11167 27795
rect 11192 27774 11227 27795
rect 11227 27774 11248 27795
rect 11111 27760 11167 27774
rect 11192 27760 11248 27774
rect 11111 27739 11161 27760
rect 11161 27739 11167 27760
rect 11192 27739 11227 27760
rect 11227 27739 11248 27760
rect 11273 27739 11329 27795
rect 11354 27739 11410 27795
rect 11435 27739 11491 27795
rect 11516 27739 11572 27795
rect 11597 27739 11653 27795
rect 11678 27739 11734 27795
rect 11759 27739 11815 27795
rect 11840 27739 11896 27795
rect 11921 27774 11945 27795
rect 11945 27774 11977 27795
rect 12002 27774 12011 27795
rect 12011 27774 12058 27795
rect 11921 27760 11977 27774
rect 12002 27760 12058 27774
rect 11921 27739 11945 27760
rect 11945 27739 11977 27760
rect 12002 27739 12011 27760
rect 12011 27739 12058 27760
rect 3452 27652 3508 27708
rect 3532 27652 3588 27708
rect 3612 27652 3668 27708
rect 3693 27652 3749 27708
rect 3774 27652 3830 27708
rect 3855 27652 3911 27708
rect 3936 27652 3992 27708
rect 4017 27652 4073 27708
rect 4098 27652 4154 27708
rect 4179 27652 4235 27708
rect 4260 27652 4316 27708
rect 5215 27694 5271 27707
rect 5296 27694 5352 27707
rect 5215 27651 5257 27694
rect 5257 27651 5271 27694
rect 5296 27651 5309 27694
rect 5309 27651 5323 27694
rect 5323 27651 5352 27694
rect 5377 27651 5433 27707
rect 5458 27651 5514 27707
rect 5539 27651 5595 27707
rect 5620 27651 5676 27707
rect 5701 27651 5757 27707
rect 5782 27651 5838 27707
rect 5863 27651 5919 27707
rect 5944 27651 6000 27707
rect 6025 27651 6081 27707
rect 6106 27694 6162 27707
rect 6186 27694 6242 27707
rect 6106 27651 6145 27694
rect 6145 27651 6159 27694
rect 6159 27651 6162 27694
rect 6186 27651 6211 27694
rect 6211 27651 6242 27694
rect 6266 27651 6322 27707
rect 6346 27651 6402 27707
rect 8572 27694 8628 27707
rect 8652 27694 8708 27707
rect 8572 27651 8601 27694
rect 8601 27651 8628 27694
rect 8652 27651 8653 27694
rect 8653 27651 8667 27694
rect 8667 27651 8708 27694
rect 8732 27651 8788 27707
rect 8812 27651 8868 27707
rect 8893 27651 8949 27707
rect 8974 27651 9030 27707
rect 9055 27651 9111 27707
rect 9136 27651 9192 27707
rect 9217 27651 9273 27707
rect 9298 27651 9354 27707
rect 9379 27651 9435 27707
rect 9460 27694 9516 27707
rect 9541 27694 9597 27707
rect 9460 27651 9489 27694
rect 9489 27651 9503 27694
rect 9503 27651 9516 27694
rect 9541 27651 9555 27694
rect 9555 27651 9597 27694
rect 9622 27651 9678 27707
rect 9703 27651 9759 27707
rect 10871 27651 10927 27707
rect 10951 27651 11007 27707
rect 11031 27651 11087 27707
rect 11111 27694 11167 27707
rect 11192 27694 11248 27707
rect 11111 27651 11161 27694
rect 11161 27651 11167 27694
rect 11192 27651 11227 27694
rect 11227 27651 11248 27694
rect 11273 27651 11329 27707
rect 11354 27651 11410 27707
rect 11435 27651 11491 27707
rect 11516 27651 11572 27707
rect 11597 27651 11653 27707
rect 11678 27651 11734 27707
rect 11759 27651 11815 27707
rect 11840 27651 11896 27707
rect 11921 27694 11977 27707
rect 12002 27694 12058 27707
rect 11921 27651 11945 27694
rect 11945 27651 11977 27694
rect 12002 27651 12011 27694
rect 12011 27651 12058 27694
rect 3452 27558 3508 27614
rect 3532 27558 3588 27614
rect 3612 27558 3668 27614
rect 3693 27558 3749 27614
rect 3774 27558 3830 27614
rect 3855 27558 3911 27614
rect 3936 27558 3992 27614
rect 4017 27558 4073 27614
rect 4098 27558 4154 27614
rect 4179 27558 4235 27614
rect 4260 27558 4316 27614
rect 5215 27575 5257 27619
rect 5257 27575 5271 27619
rect 5296 27575 5309 27619
rect 5309 27575 5323 27619
rect 5323 27575 5352 27619
rect 5215 27563 5271 27575
rect 5296 27563 5352 27575
rect 5377 27563 5433 27619
rect 5458 27563 5514 27619
rect 5539 27563 5595 27619
rect 5620 27563 5676 27619
rect 5701 27563 5757 27619
rect 5782 27563 5838 27619
rect 5863 27563 5919 27619
rect 5944 27563 6000 27619
rect 6025 27563 6081 27619
rect 6106 27575 6145 27619
rect 6145 27575 6159 27619
rect 6159 27575 6162 27619
rect 6186 27575 6211 27619
rect 6211 27575 6242 27619
rect 6106 27563 6162 27575
rect 6186 27563 6242 27575
rect 6266 27563 6322 27619
rect 6346 27563 6402 27619
rect 8572 27575 8601 27619
rect 8601 27575 8628 27619
rect 8652 27575 8653 27619
rect 8653 27575 8667 27619
rect 8667 27575 8708 27619
rect 8572 27563 8628 27575
rect 8652 27563 8708 27575
rect 8732 27563 8788 27619
rect 8812 27563 8868 27619
rect 8893 27563 8949 27619
rect 8974 27563 9030 27619
rect 9055 27563 9111 27619
rect 9136 27563 9192 27619
rect 9217 27563 9273 27619
rect 9298 27563 9354 27619
rect 9379 27563 9435 27619
rect 9460 27575 9489 27619
rect 9489 27575 9503 27619
rect 9503 27575 9516 27619
rect 9541 27575 9555 27619
rect 9555 27575 9597 27619
rect 9460 27563 9516 27575
rect 9541 27563 9597 27575
rect 9622 27563 9678 27619
rect 9703 27563 9759 27619
rect 10871 27563 10927 27619
rect 10951 27563 11007 27619
rect 11031 27563 11087 27619
rect 11111 27575 11161 27619
rect 11161 27575 11167 27619
rect 11192 27575 11227 27619
rect 11227 27575 11248 27619
rect 11111 27563 11167 27575
rect 11192 27563 11248 27575
rect 11273 27563 11329 27619
rect 11354 27563 11410 27619
rect 11435 27563 11491 27619
rect 11516 27563 11572 27619
rect 11597 27563 11653 27619
rect 11678 27563 11734 27619
rect 11759 27563 11815 27619
rect 11840 27563 11896 27619
rect 11921 27575 11945 27619
rect 11945 27575 11977 27619
rect 12002 27575 12011 27619
rect 12011 27575 12058 27619
rect 11921 27563 11977 27575
rect 12002 27563 12058 27575
rect 3452 27464 3508 27520
rect 3532 27464 3588 27520
rect 3612 27464 3668 27520
rect 3693 27464 3749 27520
rect 3774 27464 3830 27520
rect 3855 27464 3911 27520
rect 3936 27464 3992 27520
rect 4017 27464 4073 27520
rect 4098 27464 4154 27520
rect 4179 27464 4235 27520
rect 4260 27464 4316 27520
rect 5215 27508 5257 27531
rect 5257 27508 5271 27531
rect 5296 27508 5309 27531
rect 5309 27508 5323 27531
rect 5323 27508 5352 27531
rect 5215 27493 5271 27508
rect 5296 27493 5352 27508
rect 5215 27475 5257 27493
rect 5257 27475 5271 27493
rect 5296 27475 5309 27493
rect 5309 27475 5323 27493
rect 5323 27475 5352 27493
rect 5377 27475 5433 27531
rect 5458 27475 5514 27531
rect 5539 27475 5595 27531
rect 5620 27475 5676 27531
rect 5701 27475 5757 27531
rect 5782 27475 5838 27531
rect 5863 27475 5919 27531
rect 5944 27475 6000 27531
rect 6025 27475 6081 27531
rect 6106 27508 6145 27531
rect 6145 27508 6159 27531
rect 6159 27508 6162 27531
rect 6186 27508 6211 27531
rect 6211 27508 6242 27531
rect 6106 27493 6162 27508
rect 6186 27493 6242 27508
rect 6106 27475 6145 27493
rect 6145 27475 6159 27493
rect 6159 27475 6162 27493
rect 6186 27475 6211 27493
rect 6211 27475 6242 27493
rect 6266 27475 6322 27531
rect 6346 27475 6402 27531
rect 8572 27508 8601 27531
rect 8601 27508 8628 27531
rect 8652 27508 8653 27531
rect 8653 27508 8667 27531
rect 8667 27508 8708 27531
rect 8572 27493 8628 27508
rect 8652 27493 8708 27508
rect 5215 27441 5257 27443
rect 5257 27441 5271 27443
rect 5296 27441 5309 27443
rect 5309 27441 5323 27443
rect 5323 27441 5352 27443
rect 5215 27426 5271 27441
rect 5296 27426 5352 27441
rect 3452 27370 3508 27426
rect 3532 27370 3588 27426
rect 3612 27370 3668 27426
rect 3693 27370 3749 27426
rect 3774 27370 3830 27426
rect 3855 27370 3911 27426
rect 3936 27370 3992 27426
rect 4017 27370 4073 27426
rect 4098 27370 4154 27426
rect 4179 27370 4235 27426
rect 4260 27370 4316 27426
rect 5215 27387 5257 27426
rect 5257 27387 5271 27426
rect 5296 27387 5309 27426
rect 5309 27387 5323 27426
rect 5323 27387 5352 27426
rect 5377 27387 5433 27443
rect 5458 27387 5514 27443
rect 5539 27387 5595 27443
rect 5620 27387 5676 27443
rect 5701 27387 5757 27443
rect 5782 27387 5838 27443
rect 5863 27387 5919 27443
rect 5944 27387 6000 27443
rect 6025 27387 6081 27443
rect 6106 27441 6145 27443
rect 6145 27441 6159 27443
rect 6159 27441 6162 27443
rect 6186 27441 6211 27443
rect 6211 27441 6242 27443
rect 6106 27426 6162 27441
rect 6186 27426 6242 27441
rect 6106 27387 6145 27426
rect 6145 27387 6159 27426
rect 6159 27387 6162 27426
rect 6186 27387 6211 27426
rect 6211 27387 6242 27426
rect 6266 27387 6322 27443
rect 6346 27387 6402 27443
rect 8572 27475 8601 27493
rect 8601 27475 8628 27493
rect 8652 27475 8653 27493
rect 8653 27475 8667 27493
rect 8667 27475 8708 27493
rect 8732 27475 8788 27531
rect 8812 27475 8868 27531
rect 8893 27475 8949 27531
rect 8974 27475 9030 27531
rect 9055 27475 9111 27531
rect 9136 27475 9192 27531
rect 9217 27475 9273 27531
rect 9298 27475 9354 27531
rect 9379 27475 9435 27531
rect 9460 27508 9489 27531
rect 9489 27508 9503 27531
rect 9503 27508 9516 27531
rect 9541 27508 9555 27531
rect 9555 27508 9597 27531
rect 9460 27493 9516 27508
rect 9541 27493 9597 27508
rect 9460 27475 9489 27493
rect 9489 27475 9503 27493
rect 9503 27475 9516 27493
rect 9541 27475 9555 27493
rect 9555 27475 9597 27493
rect 9622 27475 9678 27531
rect 9703 27475 9759 27531
rect 8572 27441 8601 27443
rect 8601 27441 8628 27443
rect 8652 27441 8653 27443
rect 8653 27441 8667 27443
rect 8667 27441 8708 27443
rect 8572 27426 8628 27441
rect 8652 27426 8708 27441
rect 8572 27387 8601 27426
rect 8601 27387 8628 27426
rect 8652 27387 8653 27426
rect 8653 27387 8667 27426
rect 8667 27387 8708 27426
rect 8732 27387 8788 27443
rect 8812 27387 8868 27443
rect 8893 27387 8949 27443
rect 8974 27387 9030 27443
rect 9055 27387 9111 27443
rect 9136 27387 9192 27443
rect 9217 27387 9273 27443
rect 9298 27387 9354 27443
rect 9379 27387 9435 27443
rect 9460 27441 9489 27443
rect 9489 27441 9503 27443
rect 9503 27441 9516 27443
rect 9541 27441 9555 27443
rect 9555 27441 9597 27443
rect 9460 27426 9516 27441
rect 9541 27426 9597 27441
rect 9460 27387 9489 27426
rect 9489 27387 9503 27426
rect 9503 27387 9516 27426
rect 9541 27387 9555 27426
rect 9555 27387 9597 27426
rect 9622 27387 9678 27443
rect 9703 27387 9759 27443
rect 10871 27475 10927 27531
rect 10951 27475 11007 27531
rect 11031 27475 11087 27531
rect 11111 27508 11161 27531
rect 11161 27508 11167 27531
rect 11192 27508 11227 27531
rect 11227 27508 11248 27531
rect 11111 27493 11167 27508
rect 11192 27493 11248 27508
rect 11111 27475 11161 27493
rect 11161 27475 11167 27493
rect 11192 27475 11227 27493
rect 11227 27475 11248 27493
rect 11273 27475 11329 27531
rect 11354 27475 11410 27531
rect 11435 27475 11491 27531
rect 11516 27475 11572 27531
rect 11597 27475 11653 27531
rect 11678 27475 11734 27531
rect 11759 27475 11815 27531
rect 11840 27475 11896 27531
rect 11921 27508 11945 27531
rect 11945 27508 11977 27531
rect 12002 27508 12011 27531
rect 12011 27508 12058 27531
rect 11921 27493 11977 27508
rect 12002 27493 12058 27508
rect 11921 27475 11945 27493
rect 11945 27475 11977 27493
rect 12002 27475 12011 27493
rect 12011 27475 12058 27493
rect 10871 27387 10927 27443
rect 10951 27387 11007 27443
rect 11031 27387 11087 27443
rect 11111 27441 11161 27443
rect 11161 27441 11167 27443
rect 11192 27441 11227 27443
rect 11227 27441 11248 27443
rect 11111 27426 11167 27441
rect 11192 27426 11248 27441
rect 11111 27387 11161 27426
rect 11161 27387 11167 27426
rect 11192 27387 11227 27426
rect 11227 27387 11248 27426
rect 11273 27387 11329 27443
rect 11354 27387 11410 27443
rect 11435 27387 11491 27443
rect 11516 27387 11572 27443
rect 11597 27387 11653 27443
rect 11678 27387 11734 27443
rect 11759 27387 11815 27443
rect 11840 27387 11896 27443
rect 11921 27441 11945 27443
rect 11945 27441 11977 27443
rect 12002 27441 12011 27443
rect 12011 27441 12058 27443
rect 11921 27426 11977 27441
rect 12002 27426 12058 27441
rect 11921 27387 11945 27426
rect 11945 27387 11977 27426
rect 12002 27387 12011 27426
rect 12011 27387 12058 27426
rect 3443 25826 3499 25882
rect 3525 25826 3581 25882
rect 3607 25826 3663 25882
rect 3689 25826 3745 25882
rect 3771 25826 3827 25882
rect 3853 25826 3909 25882
rect 3935 25826 3991 25882
rect 4017 25826 4073 25882
rect 4098 25826 4154 25882
rect 4179 25826 4235 25882
rect 4260 25826 4316 25882
rect 5215 25839 5257 25882
rect 5257 25839 5271 25882
rect 5296 25839 5309 25882
rect 5309 25839 5323 25882
rect 5323 25839 5352 25882
rect 5215 25826 5271 25839
rect 5296 25826 5352 25839
rect 5377 25826 5433 25882
rect 5458 25826 5514 25882
rect 5539 25826 5595 25882
rect 5620 25826 5676 25882
rect 5701 25826 5757 25882
rect 5782 25826 5838 25882
rect 5863 25826 5919 25882
rect 5944 25826 6000 25882
rect 6025 25826 6081 25882
rect 6106 25839 6145 25882
rect 6145 25839 6159 25882
rect 6159 25839 6162 25882
rect 6186 25839 6211 25882
rect 6211 25839 6242 25882
rect 6106 25826 6162 25839
rect 6186 25826 6242 25839
rect 6266 25826 6322 25882
rect 6346 25826 6402 25882
rect 8572 25839 8601 25882
rect 8601 25839 8628 25882
rect 8652 25839 8653 25882
rect 8653 25839 8667 25882
rect 8667 25839 8708 25882
rect 8572 25826 8628 25839
rect 8652 25826 8708 25839
rect 8732 25826 8788 25882
rect 8812 25826 8868 25882
rect 8893 25826 8949 25882
rect 8974 25826 9030 25882
rect 9055 25826 9111 25882
rect 9136 25826 9192 25882
rect 9217 25826 9273 25882
rect 9298 25826 9354 25882
rect 9379 25826 9435 25882
rect 9460 25839 9489 25882
rect 9489 25839 9503 25882
rect 9503 25839 9516 25882
rect 9541 25839 9555 25882
rect 9555 25839 9597 25882
rect 9460 25826 9516 25839
rect 9541 25826 9597 25839
rect 9622 25826 9678 25882
rect 9703 25826 9759 25882
rect 10871 25826 10927 25882
rect 10951 25826 11007 25882
rect 11031 25826 11087 25882
rect 11111 25839 11161 25882
rect 11161 25839 11167 25882
rect 11192 25839 11227 25882
rect 11227 25839 11248 25882
rect 11111 25826 11167 25839
rect 11192 25826 11248 25839
rect 11273 25826 11329 25882
rect 11354 25826 11410 25882
rect 11435 25826 11491 25882
rect 11516 25826 11572 25882
rect 11597 25826 11653 25882
rect 11678 25826 11734 25882
rect 11759 25826 11815 25882
rect 11840 25826 11896 25882
rect 11921 25839 11945 25882
rect 11945 25839 11977 25882
rect 12002 25839 12011 25882
rect 12011 25839 12058 25882
rect 11921 25826 11977 25839
rect 12002 25826 12058 25839
rect 3443 25738 3499 25794
rect 3525 25738 3581 25794
rect 3607 25738 3663 25794
rect 3689 25738 3745 25794
rect 3771 25738 3827 25794
rect 3853 25738 3909 25794
rect 3935 25738 3991 25794
rect 4017 25738 4073 25794
rect 4098 25738 4154 25794
rect 4179 25738 4235 25794
rect 4260 25738 4316 25794
rect 5215 25773 5257 25794
rect 5257 25773 5271 25794
rect 5296 25773 5309 25794
rect 5309 25773 5323 25794
rect 5323 25773 5352 25794
rect 5215 25759 5271 25773
rect 5296 25759 5352 25773
rect 5215 25738 5257 25759
rect 5257 25738 5271 25759
rect 5296 25738 5309 25759
rect 5309 25738 5323 25759
rect 5323 25738 5352 25759
rect 5377 25738 5433 25794
rect 5458 25738 5514 25794
rect 5539 25738 5595 25794
rect 5620 25738 5676 25794
rect 5701 25738 5757 25794
rect 5782 25738 5838 25794
rect 5863 25738 5919 25794
rect 5944 25738 6000 25794
rect 6025 25738 6081 25794
rect 6106 25773 6145 25794
rect 6145 25773 6159 25794
rect 6159 25773 6162 25794
rect 6186 25773 6211 25794
rect 6211 25773 6242 25794
rect 6106 25759 6162 25773
rect 6186 25759 6242 25773
rect 6106 25738 6145 25759
rect 6145 25738 6159 25759
rect 6159 25738 6162 25759
rect 6186 25738 6211 25759
rect 6211 25738 6242 25759
rect 6266 25738 6322 25794
rect 6346 25738 6402 25794
rect 8572 25773 8601 25794
rect 8601 25773 8628 25794
rect 8652 25773 8653 25794
rect 8653 25773 8667 25794
rect 8667 25773 8708 25794
rect 8572 25759 8628 25773
rect 8652 25759 8708 25773
rect 8572 25738 8601 25759
rect 8601 25738 8628 25759
rect 8652 25738 8653 25759
rect 8653 25738 8667 25759
rect 8667 25738 8708 25759
rect 8732 25738 8788 25794
rect 8812 25738 8868 25794
rect 8893 25738 8949 25794
rect 8974 25738 9030 25794
rect 9055 25738 9111 25794
rect 9136 25738 9192 25794
rect 9217 25738 9273 25794
rect 9298 25738 9354 25794
rect 9379 25738 9435 25794
rect 9460 25773 9489 25794
rect 9489 25773 9503 25794
rect 9503 25773 9516 25794
rect 9541 25773 9555 25794
rect 9555 25773 9597 25794
rect 9460 25759 9516 25773
rect 9541 25759 9597 25773
rect 9460 25738 9489 25759
rect 9489 25738 9503 25759
rect 9503 25738 9516 25759
rect 9541 25738 9555 25759
rect 9555 25738 9597 25759
rect 9622 25738 9678 25794
rect 9703 25738 9759 25794
rect 10871 25738 10927 25794
rect 10951 25738 11007 25794
rect 11031 25738 11087 25794
rect 11111 25773 11161 25794
rect 11161 25773 11167 25794
rect 11192 25773 11227 25794
rect 11227 25773 11248 25794
rect 11111 25759 11167 25773
rect 11192 25759 11248 25773
rect 11111 25738 11161 25759
rect 11161 25738 11167 25759
rect 11192 25738 11227 25759
rect 11227 25738 11248 25759
rect 11273 25738 11329 25794
rect 11354 25738 11410 25794
rect 11435 25738 11491 25794
rect 11516 25738 11572 25794
rect 11597 25738 11653 25794
rect 11678 25738 11734 25794
rect 11759 25738 11815 25794
rect 11840 25738 11896 25794
rect 11921 25773 11945 25794
rect 11945 25773 11977 25794
rect 12002 25773 12011 25794
rect 12011 25773 12058 25794
rect 11921 25759 11977 25773
rect 12002 25759 12058 25773
rect 11921 25738 11945 25759
rect 11945 25738 11977 25759
rect 12002 25738 12011 25759
rect 12011 25738 12058 25759
rect 3443 25650 3499 25706
rect 3525 25650 3581 25706
rect 3607 25650 3663 25706
rect 3689 25650 3745 25706
rect 3771 25650 3827 25706
rect 3853 25650 3909 25706
rect 3935 25650 3991 25706
rect 4017 25650 4073 25706
rect 4098 25650 4154 25706
rect 4179 25650 4235 25706
rect 4260 25650 4316 25706
rect 5215 25693 5271 25706
rect 5296 25693 5352 25706
rect 5215 25650 5257 25693
rect 5257 25650 5271 25693
rect 5296 25650 5309 25693
rect 5309 25650 5323 25693
rect 5323 25650 5352 25693
rect 5377 25650 5433 25706
rect 5458 25650 5514 25706
rect 5539 25650 5595 25706
rect 5620 25650 5676 25706
rect 5701 25650 5757 25706
rect 5782 25650 5838 25706
rect 5863 25650 5919 25706
rect 5944 25650 6000 25706
rect 6025 25650 6081 25706
rect 6106 25693 6162 25706
rect 6186 25693 6242 25706
rect 6106 25650 6145 25693
rect 6145 25650 6159 25693
rect 6159 25650 6162 25693
rect 6186 25650 6211 25693
rect 6211 25650 6242 25693
rect 6266 25650 6322 25706
rect 6346 25650 6402 25706
rect 8572 25693 8628 25706
rect 8652 25693 8708 25706
rect 8572 25650 8601 25693
rect 8601 25650 8628 25693
rect 8652 25650 8653 25693
rect 8653 25650 8667 25693
rect 8667 25650 8708 25693
rect 8732 25650 8788 25706
rect 8812 25650 8868 25706
rect 8893 25650 8949 25706
rect 8974 25650 9030 25706
rect 9055 25650 9111 25706
rect 9136 25650 9192 25706
rect 9217 25650 9273 25706
rect 9298 25650 9354 25706
rect 9379 25650 9435 25706
rect 9460 25693 9516 25706
rect 9541 25693 9597 25706
rect 9460 25650 9489 25693
rect 9489 25650 9503 25693
rect 9503 25650 9516 25693
rect 9541 25650 9555 25693
rect 9555 25650 9597 25693
rect 9622 25650 9678 25706
rect 9703 25650 9759 25706
rect 10871 25650 10927 25706
rect 10951 25650 11007 25706
rect 11031 25650 11087 25706
rect 11111 25693 11167 25706
rect 11192 25693 11248 25706
rect 11111 25650 11161 25693
rect 11161 25650 11167 25693
rect 11192 25650 11227 25693
rect 11227 25650 11248 25693
rect 11273 25650 11329 25706
rect 11354 25650 11410 25706
rect 11435 25650 11491 25706
rect 11516 25650 11572 25706
rect 11597 25650 11653 25706
rect 11678 25650 11734 25706
rect 11759 25650 11815 25706
rect 11840 25650 11896 25706
rect 11921 25693 11977 25706
rect 12002 25693 12058 25706
rect 11921 25650 11945 25693
rect 11945 25650 11977 25693
rect 12002 25650 12011 25693
rect 12011 25650 12058 25693
rect 3443 25562 3499 25618
rect 3525 25562 3581 25618
rect 3607 25562 3663 25618
rect 3689 25562 3745 25618
rect 3771 25562 3827 25618
rect 3853 25562 3909 25618
rect 3935 25562 3991 25618
rect 4017 25562 4073 25618
rect 4098 25562 4154 25618
rect 4179 25562 4235 25618
rect 4260 25562 4316 25618
rect 5215 25574 5257 25618
rect 5257 25574 5271 25618
rect 5296 25574 5309 25618
rect 5309 25574 5323 25618
rect 5323 25574 5352 25618
rect 5215 25562 5271 25574
rect 5296 25562 5352 25574
rect 5377 25562 5433 25618
rect 5458 25562 5514 25618
rect 5539 25562 5595 25618
rect 5620 25562 5676 25618
rect 5701 25562 5757 25618
rect 5782 25562 5838 25618
rect 5863 25562 5919 25618
rect 5944 25562 6000 25618
rect 6025 25562 6081 25618
rect 6106 25574 6145 25618
rect 6145 25574 6159 25618
rect 6159 25574 6162 25618
rect 6186 25574 6211 25618
rect 6211 25574 6242 25618
rect 6106 25562 6162 25574
rect 6186 25562 6242 25574
rect 6266 25562 6322 25618
rect 6346 25562 6402 25618
rect 8572 25574 8601 25618
rect 8601 25574 8628 25618
rect 8652 25574 8653 25618
rect 8653 25574 8667 25618
rect 8667 25574 8708 25618
rect 8572 25562 8628 25574
rect 8652 25562 8708 25574
rect 8732 25562 8788 25618
rect 8812 25562 8868 25618
rect 8893 25562 8949 25618
rect 8974 25562 9030 25618
rect 9055 25562 9111 25618
rect 9136 25562 9192 25618
rect 9217 25562 9273 25618
rect 9298 25562 9354 25618
rect 9379 25562 9435 25618
rect 9460 25574 9489 25618
rect 9489 25574 9503 25618
rect 9503 25574 9516 25618
rect 9541 25574 9555 25618
rect 9555 25574 9597 25618
rect 9460 25562 9516 25574
rect 9541 25562 9597 25574
rect 9622 25562 9678 25618
rect 9703 25562 9759 25618
rect 10871 25562 10927 25618
rect 10951 25562 11007 25618
rect 11031 25562 11087 25618
rect 11111 25574 11161 25618
rect 11161 25574 11167 25618
rect 11192 25574 11227 25618
rect 11227 25574 11248 25618
rect 11111 25562 11167 25574
rect 11192 25562 11248 25574
rect 11273 25562 11329 25618
rect 11354 25562 11410 25618
rect 11435 25562 11491 25618
rect 11516 25562 11572 25618
rect 11597 25562 11653 25618
rect 11678 25562 11734 25618
rect 11759 25562 11815 25618
rect 11840 25562 11896 25618
rect 11921 25574 11945 25618
rect 11945 25574 11977 25618
rect 12002 25574 12011 25618
rect 12011 25574 12058 25618
rect 11921 25562 11977 25574
rect 12002 25562 12058 25574
rect 3443 25474 3499 25530
rect 3525 25474 3581 25530
rect 3607 25474 3663 25530
rect 3689 25474 3745 25530
rect 3771 25474 3827 25530
rect 3853 25474 3909 25530
rect 3935 25474 3991 25530
rect 4017 25474 4073 25530
rect 4098 25474 4154 25530
rect 4179 25474 4235 25530
rect 4260 25474 4316 25530
rect 5215 25507 5257 25530
rect 5257 25507 5271 25530
rect 5296 25507 5309 25530
rect 5309 25507 5323 25530
rect 5323 25507 5352 25530
rect 5215 25492 5271 25507
rect 5296 25492 5352 25507
rect 5215 25474 5257 25492
rect 5257 25474 5271 25492
rect 5296 25474 5309 25492
rect 5309 25474 5323 25492
rect 5323 25474 5352 25492
rect 5377 25474 5433 25530
rect 5458 25474 5514 25530
rect 5539 25474 5595 25530
rect 5620 25474 5676 25530
rect 5701 25474 5757 25530
rect 5782 25474 5838 25530
rect 5863 25474 5919 25530
rect 5944 25474 6000 25530
rect 6025 25474 6081 25530
rect 6106 25507 6145 25530
rect 6145 25507 6159 25530
rect 6159 25507 6162 25530
rect 6186 25507 6211 25530
rect 6211 25507 6242 25530
rect 6106 25492 6162 25507
rect 6186 25492 6242 25507
rect 6106 25474 6145 25492
rect 6145 25474 6159 25492
rect 6159 25474 6162 25492
rect 6186 25474 6211 25492
rect 6211 25474 6242 25492
rect 6266 25474 6322 25530
rect 6346 25474 6402 25530
rect 8572 25507 8601 25530
rect 8601 25507 8628 25530
rect 8652 25507 8653 25530
rect 8653 25507 8667 25530
rect 8667 25507 8708 25530
rect 8572 25492 8628 25507
rect 8652 25492 8708 25507
rect 3443 25386 3499 25442
rect 3525 25386 3581 25442
rect 3607 25386 3663 25442
rect 3689 25386 3745 25442
rect 3771 25386 3827 25442
rect 3853 25386 3909 25442
rect 3935 25386 3991 25442
rect 4017 25386 4073 25442
rect 4098 25386 4154 25442
rect 4179 25386 4235 25442
rect 4260 25386 4316 25442
rect 5215 25440 5257 25442
rect 5257 25440 5271 25442
rect 5296 25440 5309 25442
rect 5309 25440 5323 25442
rect 5323 25440 5352 25442
rect 5215 25425 5271 25440
rect 5296 25425 5352 25440
rect 5215 25386 5257 25425
rect 5257 25386 5271 25425
rect 5296 25386 5309 25425
rect 5309 25386 5323 25425
rect 5323 25386 5352 25425
rect 5377 25386 5433 25442
rect 5458 25386 5514 25442
rect 5539 25386 5595 25442
rect 5620 25386 5676 25442
rect 5701 25386 5757 25442
rect 5782 25386 5838 25442
rect 5863 25386 5919 25442
rect 5944 25386 6000 25442
rect 6025 25386 6081 25442
rect 6106 25440 6145 25442
rect 6145 25440 6159 25442
rect 6159 25440 6162 25442
rect 6186 25440 6211 25442
rect 6211 25440 6242 25442
rect 6106 25425 6162 25440
rect 6186 25425 6242 25440
rect 6106 25386 6145 25425
rect 6145 25386 6159 25425
rect 6159 25386 6162 25425
rect 6186 25386 6211 25425
rect 6211 25386 6242 25425
rect 6266 25386 6322 25442
rect 6346 25386 6402 25442
rect 8572 25474 8601 25492
rect 8601 25474 8628 25492
rect 8652 25474 8653 25492
rect 8653 25474 8667 25492
rect 8667 25474 8708 25492
rect 8732 25474 8788 25530
rect 8812 25474 8868 25530
rect 8893 25474 8949 25530
rect 8974 25474 9030 25530
rect 9055 25474 9111 25530
rect 9136 25474 9192 25530
rect 9217 25474 9273 25530
rect 9298 25474 9354 25530
rect 9379 25474 9435 25530
rect 9460 25507 9489 25530
rect 9489 25507 9503 25530
rect 9503 25507 9516 25530
rect 9541 25507 9555 25530
rect 9555 25507 9597 25530
rect 9460 25492 9516 25507
rect 9541 25492 9597 25507
rect 9460 25474 9489 25492
rect 9489 25474 9503 25492
rect 9503 25474 9516 25492
rect 9541 25474 9555 25492
rect 9555 25474 9597 25492
rect 9622 25474 9678 25530
rect 9703 25474 9759 25530
rect 8572 25440 8601 25442
rect 8601 25440 8628 25442
rect 8652 25440 8653 25442
rect 8653 25440 8667 25442
rect 8667 25440 8708 25442
rect 8572 25425 8628 25440
rect 8652 25425 8708 25440
rect 8572 25386 8601 25425
rect 8601 25386 8628 25425
rect 8652 25386 8653 25425
rect 8653 25386 8667 25425
rect 8667 25386 8708 25425
rect 8732 25386 8788 25442
rect 8812 25386 8868 25442
rect 8893 25386 8949 25442
rect 8974 25386 9030 25442
rect 9055 25386 9111 25442
rect 9136 25386 9192 25442
rect 9217 25386 9273 25442
rect 9298 25386 9354 25442
rect 9379 25386 9435 25442
rect 9460 25440 9489 25442
rect 9489 25440 9503 25442
rect 9503 25440 9516 25442
rect 9541 25440 9555 25442
rect 9555 25440 9597 25442
rect 9460 25425 9516 25440
rect 9541 25425 9597 25440
rect 9460 25386 9489 25425
rect 9489 25386 9503 25425
rect 9503 25386 9516 25425
rect 9541 25386 9555 25425
rect 9555 25386 9597 25425
rect 9622 25386 9678 25442
rect 9703 25386 9759 25442
rect 10871 25474 10927 25530
rect 10951 25474 11007 25530
rect 11031 25474 11087 25530
rect 11111 25507 11161 25530
rect 11161 25507 11167 25530
rect 11192 25507 11227 25530
rect 11227 25507 11248 25530
rect 11111 25492 11167 25507
rect 11192 25492 11248 25507
rect 11111 25474 11161 25492
rect 11161 25474 11167 25492
rect 11192 25474 11227 25492
rect 11227 25474 11248 25492
rect 11273 25474 11329 25530
rect 11354 25474 11410 25530
rect 11435 25474 11491 25530
rect 11516 25474 11572 25530
rect 11597 25474 11653 25530
rect 11678 25474 11734 25530
rect 11759 25474 11815 25530
rect 11840 25474 11896 25530
rect 11921 25507 11945 25530
rect 11945 25507 11977 25530
rect 12002 25507 12011 25530
rect 12011 25507 12058 25530
rect 11921 25492 11977 25507
rect 12002 25492 12058 25507
rect 11921 25474 11945 25492
rect 11945 25474 11977 25492
rect 12002 25474 12011 25492
rect 12011 25474 12058 25492
rect 10871 25386 10927 25442
rect 10951 25386 11007 25442
rect 11031 25386 11087 25442
rect 11111 25440 11161 25442
rect 11161 25440 11167 25442
rect 11192 25440 11227 25442
rect 11227 25440 11248 25442
rect 11111 25425 11167 25440
rect 11192 25425 11248 25440
rect 11111 25386 11161 25425
rect 11161 25386 11167 25425
rect 11192 25386 11227 25425
rect 11227 25386 11248 25425
rect 11273 25386 11329 25442
rect 11354 25386 11410 25442
rect 11435 25386 11491 25442
rect 11516 25386 11572 25442
rect 11597 25386 11653 25442
rect 11678 25386 11734 25442
rect 11759 25386 11815 25442
rect 11840 25386 11896 25442
rect 11921 25440 11945 25442
rect 11945 25440 11977 25442
rect 12002 25440 12011 25442
rect 12011 25440 12058 25442
rect 11921 25425 11977 25440
rect 12002 25425 12058 25440
rect 11921 25386 11945 25425
rect 11945 25386 11977 25425
rect 12002 25386 12011 25425
rect 12011 25386 12058 25425
rect 7691 13821 7747 13877
rect 7775 13821 7831 13877
rect 7858 13821 7914 13877
rect 7941 13840 7988 13877
rect 7988 13840 7997 13877
rect 8024 13840 8054 13877
rect 8054 13840 8080 13877
rect 7941 13826 7997 13840
rect 8024 13826 8080 13840
rect 7941 13821 7988 13826
rect 7988 13821 7997 13826
rect 8024 13821 8054 13826
rect 8054 13821 8080 13826
rect 8107 13821 8163 13877
rect 8190 13821 8246 13877
rect 8273 13821 8329 13877
rect 8356 13821 8412 13877
rect 8439 13840 8490 13877
rect 8490 13840 8495 13877
rect 8522 13840 8542 13877
rect 8542 13840 8556 13877
rect 8556 13840 8578 13877
rect 8605 13840 8608 13877
rect 8608 13840 8661 13877
rect 8439 13826 8495 13840
rect 8522 13826 8578 13840
rect 8605 13826 8661 13840
rect 8439 13821 8490 13826
rect 8490 13821 8495 13826
rect 8522 13821 8542 13826
rect 8542 13821 8556 13826
rect 8556 13821 8578 13826
rect 8605 13821 8608 13826
rect 8608 13821 8661 13826
rect 8688 13821 8744 13877
rect 8771 13821 8827 13877
rect 8854 13821 8910 13877
rect 8937 13821 8993 13877
rect 9020 13840 9044 13877
rect 9044 13840 9076 13877
rect 9103 13840 9110 13877
rect 9110 13840 9159 13877
rect 9020 13826 9076 13840
rect 9103 13826 9159 13840
rect 9020 13821 9044 13826
rect 9044 13821 9076 13826
rect 9103 13821 9110 13826
rect 9110 13821 9159 13826
rect 9186 13821 9242 13877
rect 9269 13821 9325 13877
rect 9352 13821 9408 13877
rect 9435 13821 9491 13877
rect 9518 13821 9574 13877
rect 9601 13840 9650 13877
rect 9650 13840 9657 13877
rect 9684 13840 9716 13877
rect 9716 13840 9740 13877
rect 9601 13826 9657 13840
rect 9684 13826 9740 13840
rect 9601 13821 9650 13826
rect 9650 13821 9657 13826
rect 9684 13821 9716 13826
rect 9716 13821 9740 13826
rect 9767 13821 9823 13877
rect 7691 13733 7747 13789
rect 7775 13733 7831 13789
rect 7858 13733 7914 13789
rect 7941 13774 7988 13789
rect 7988 13774 7997 13789
rect 8024 13774 8054 13789
rect 8054 13774 8080 13789
rect 7941 13760 7997 13774
rect 8024 13760 8080 13774
rect 7941 13733 7988 13760
rect 7988 13733 7997 13760
rect 8024 13733 8054 13760
rect 8054 13733 8080 13760
rect 8107 13733 8163 13789
rect 8190 13733 8246 13789
rect 8273 13733 8329 13789
rect 8356 13733 8412 13789
rect 8439 13774 8490 13789
rect 8490 13774 8495 13789
rect 8522 13774 8542 13789
rect 8542 13774 8556 13789
rect 8556 13774 8578 13789
rect 8605 13774 8608 13789
rect 8608 13774 8661 13789
rect 8439 13760 8495 13774
rect 8522 13760 8578 13774
rect 8605 13760 8661 13774
rect 8439 13733 8490 13760
rect 8490 13733 8495 13760
rect 8522 13733 8542 13760
rect 8542 13733 8556 13760
rect 8556 13733 8578 13760
rect 8605 13733 8608 13760
rect 8608 13733 8661 13760
rect 8688 13733 8744 13789
rect 8771 13733 8827 13789
rect 8854 13733 8910 13789
rect 8937 13733 8993 13789
rect 9020 13774 9044 13789
rect 9044 13774 9076 13789
rect 9103 13774 9110 13789
rect 9110 13774 9159 13789
rect 9020 13760 9076 13774
rect 9103 13760 9159 13774
rect 9020 13733 9044 13760
rect 9044 13733 9076 13760
rect 9103 13733 9110 13760
rect 9110 13733 9159 13760
rect 9186 13733 9242 13789
rect 9269 13733 9325 13789
rect 9352 13733 9408 13789
rect 9435 13733 9491 13789
rect 9518 13733 9574 13789
rect 9601 13774 9650 13789
rect 9650 13774 9657 13789
rect 9684 13774 9716 13789
rect 9716 13774 9740 13789
rect 9601 13760 9657 13774
rect 9684 13760 9740 13774
rect 9601 13733 9650 13760
rect 9650 13733 9657 13760
rect 9684 13733 9716 13760
rect 9716 13733 9740 13760
rect 9767 13733 9823 13789
rect 7691 13645 7747 13701
rect 7775 13645 7831 13701
rect 7858 13645 7914 13701
rect 7941 13694 7997 13701
rect 8024 13694 8080 13701
rect 7941 13645 7988 13694
rect 7988 13645 7997 13694
rect 8024 13645 8054 13694
rect 8054 13645 8080 13694
rect 8107 13645 8163 13701
rect 8190 13645 8246 13701
rect 8273 13645 8329 13701
rect 8356 13645 8412 13701
rect 8439 13694 8495 13701
rect 8522 13694 8578 13701
rect 8605 13694 8661 13701
rect 8439 13645 8490 13694
rect 8490 13645 8495 13694
rect 8522 13645 8542 13694
rect 8542 13645 8556 13694
rect 8556 13645 8578 13694
rect 8605 13645 8608 13694
rect 8608 13645 8661 13694
rect 8688 13645 8744 13701
rect 8771 13645 8827 13701
rect 8854 13645 8910 13701
rect 8937 13645 8993 13701
rect 9020 13694 9076 13701
rect 9103 13694 9159 13701
rect 9020 13645 9044 13694
rect 9044 13645 9076 13694
rect 9103 13645 9110 13694
rect 9110 13645 9159 13694
rect 9186 13645 9242 13701
rect 9269 13645 9325 13701
rect 9352 13645 9408 13701
rect 9435 13645 9491 13701
rect 9518 13645 9574 13701
rect 9601 13694 9657 13701
rect 9684 13694 9740 13701
rect 9601 13645 9650 13694
rect 9650 13645 9657 13694
rect 9684 13645 9716 13694
rect 9716 13645 9740 13694
rect 9767 13645 9823 13701
rect 7691 13557 7747 13613
rect 7775 13557 7831 13613
rect 7858 13557 7914 13613
rect 7941 13576 7988 13613
rect 7988 13576 7997 13613
rect 8024 13576 8054 13613
rect 8054 13576 8080 13613
rect 7941 13562 7997 13576
rect 8024 13562 8080 13576
rect 7941 13557 7988 13562
rect 7988 13557 7997 13562
rect 8024 13557 8054 13562
rect 8054 13557 8080 13562
rect 8107 13557 8163 13613
rect 8190 13557 8246 13613
rect 8273 13557 8329 13613
rect 8356 13557 8412 13613
rect 8439 13576 8490 13613
rect 8490 13576 8495 13613
rect 8522 13576 8542 13613
rect 8542 13576 8556 13613
rect 8556 13576 8578 13613
rect 8605 13576 8608 13613
rect 8608 13576 8661 13613
rect 8439 13562 8495 13576
rect 8522 13562 8578 13576
rect 8605 13562 8661 13576
rect 8439 13557 8490 13562
rect 8490 13557 8495 13562
rect 8522 13557 8542 13562
rect 8542 13557 8556 13562
rect 8556 13557 8578 13562
rect 8605 13557 8608 13562
rect 8608 13557 8661 13562
rect 8688 13557 8744 13613
rect 8771 13557 8827 13613
rect 8854 13557 8910 13613
rect 8937 13557 8993 13613
rect 9020 13576 9044 13613
rect 9044 13576 9076 13613
rect 9103 13576 9110 13613
rect 9110 13576 9159 13613
rect 9020 13562 9076 13576
rect 9103 13562 9159 13576
rect 9020 13557 9044 13562
rect 9044 13557 9076 13562
rect 9103 13557 9110 13562
rect 9110 13557 9159 13562
rect 9186 13557 9242 13613
rect 9269 13557 9325 13613
rect 9352 13557 9408 13613
rect 9435 13557 9491 13613
rect 9518 13557 9574 13613
rect 9601 13576 9650 13613
rect 9650 13576 9657 13613
rect 9684 13576 9716 13613
rect 9716 13576 9740 13613
rect 9601 13562 9657 13576
rect 9684 13562 9740 13576
rect 9601 13557 9650 13562
rect 9650 13557 9657 13562
rect 9684 13557 9716 13562
rect 9716 13557 9740 13562
rect 9767 13557 9823 13613
rect 7691 13469 7747 13525
rect 7775 13469 7831 13525
rect 7858 13469 7914 13525
rect 7941 13510 7988 13525
rect 7988 13510 7997 13525
rect 8024 13510 8054 13525
rect 8054 13510 8080 13525
rect 7941 13495 7997 13510
rect 8024 13495 8080 13510
rect 7941 13469 7988 13495
rect 7988 13469 7997 13495
rect 8024 13469 8054 13495
rect 8054 13469 8080 13495
rect 8107 13469 8163 13525
rect 8190 13469 8246 13525
rect 8273 13469 8329 13525
rect 8356 13469 8412 13525
rect 8439 13510 8490 13525
rect 8490 13510 8495 13525
rect 8522 13510 8542 13525
rect 8542 13510 8556 13525
rect 8556 13510 8578 13525
rect 8605 13510 8608 13525
rect 8608 13510 8661 13525
rect 8439 13495 8495 13510
rect 8522 13495 8578 13510
rect 8605 13495 8661 13510
rect 8439 13469 8490 13495
rect 8490 13469 8495 13495
rect 8522 13469 8542 13495
rect 8542 13469 8556 13495
rect 8556 13469 8578 13495
rect 8605 13469 8608 13495
rect 8608 13469 8661 13495
rect 8688 13469 8744 13525
rect 8771 13469 8827 13525
rect 8854 13469 8910 13525
rect 8937 13469 8993 13525
rect 9020 13510 9044 13525
rect 9044 13510 9076 13525
rect 9103 13510 9110 13525
rect 9110 13510 9159 13525
rect 9020 13495 9076 13510
rect 9103 13495 9159 13510
rect 9020 13469 9044 13495
rect 9044 13469 9076 13495
rect 9103 13469 9110 13495
rect 9110 13469 9159 13495
rect 9186 13469 9242 13525
rect 9269 13469 9325 13525
rect 9352 13469 9408 13525
rect 9435 13469 9491 13525
rect 9518 13469 9574 13525
rect 9601 13510 9650 13525
rect 9650 13510 9657 13525
rect 9684 13510 9716 13525
rect 9716 13510 9740 13525
rect 9601 13495 9657 13510
rect 9684 13495 9740 13510
rect 9601 13469 9650 13495
rect 9650 13469 9657 13495
rect 9684 13469 9716 13495
rect 9716 13469 9740 13495
rect 9767 13469 9823 13525
rect 7691 13381 7747 13437
rect 7775 13381 7831 13437
rect 7858 13381 7914 13437
rect 7941 13428 7997 13437
rect 8024 13428 8080 13437
rect 7941 13381 7988 13428
rect 7988 13381 7997 13428
rect 8024 13381 8054 13428
rect 8054 13381 8080 13428
rect 8107 13381 8163 13437
rect 8190 13381 8246 13437
rect 8273 13381 8329 13437
rect 8356 13381 8412 13437
rect 8439 13428 8495 13437
rect 8522 13428 8578 13437
rect 8605 13428 8661 13437
rect 8439 13381 8490 13428
rect 8490 13381 8495 13428
rect 8522 13381 8542 13428
rect 8542 13381 8556 13428
rect 8556 13381 8578 13428
rect 8605 13381 8608 13428
rect 8608 13381 8661 13428
rect 8688 13381 8744 13437
rect 8771 13381 8827 13437
rect 8854 13381 8910 13437
rect 8937 13381 8993 13437
rect 9020 13428 9076 13437
rect 9103 13428 9159 13437
rect 9020 13381 9044 13428
rect 9044 13381 9076 13428
rect 9103 13381 9110 13428
rect 9110 13381 9159 13428
rect 9186 13381 9242 13437
rect 9269 13381 9325 13437
rect 9352 13381 9408 13437
rect 9435 13381 9491 13437
rect 9518 13381 9574 13437
rect 9601 13428 9657 13437
rect 9684 13428 9740 13437
rect 9601 13381 9650 13428
rect 9650 13381 9657 13428
rect 9684 13381 9716 13428
rect 9716 13381 9740 13428
rect 9767 13381 9823 13437
rect 7691 11826 7747 11882
rect 7775 11826 7831 11882
rect 7858 11826 7914 11882
rect 7941 11840 7988 11882
rect 7988 11840 7997 11882
rect 8024 11840 8054 11882
rect 8054 11840 8080 11882
rect 7941 11826 7997 11840
rect 8024 11826 8080 11840
rect 8107 11826 8163 11882
rect 8190 11826 8246 11882
rect 8273 11826 8329 11882
rect 8356 11826 8412 11882
rect 8439 11840 8490 11882
rect 8490 11840 8495 11882
rect 8522 11840 8542 11882
rect 8542 11840 8556 11882
rect 8556 11840 8578 11882
rect 8605 11840 8608 11882
rect 8608 11840 8661 11882
rect 8439 11826 8495 11840
rect 8522 11826 8578 11840
rect 8605 11826 8661 11840
rect 8688 11826 8744 11882
rect 8771 11826 8827 11882
rect 8854 11826 8910 11882
rect 8937 11826 8993 11882
rect 9020 11840 9044 11882
rect 9044 11840 9076 11882
rect 9103 11840 9110 11882
rect 9110 11840 9159 11882
rect 9020 11826 9076 11840
rect 9103 11826 9159 11840
rect 9186 11826 9242 11882
rect 9269 11826 9325 11882
rect 9352 11826 9408 11882
rect 9435 11826 9491 11882
rect 9518 11826 9574 11882
rect 9601 11840 9650 11882
rect 9650 11840 9657 11882
rect 9684 11840 9716 11882
rect 9716 11840 9740 11882
rect 9601 11826 9657 11840
rect 9684 11826 9740 11840
rect 9767 11826 9823 11882
rect 7691 11738 7747 11794
rect 7775 11738 7831 11794
rect 7858 11738 7914 11794
rect 7941 11774 7988 11794
rect 7988 11774 7997 11794
rect 8024 11774 8054 11794
rect 8054 11774 8080 11794
rect 7941 11760 7997 11774
rect 8024 11760 8080 11774
rect 7941 11738 7988 11760
rect 7988 11738 7997 11760
rect 8024 11738 8054 11760
rect 8054 11738 8080 11760
rect 8107 11738 8163 11794
rect 8190 11738 8246 11794
rect 8273 11738 8329 11794
rect 8356 11738 8412 11794
rect 8439 11774 8490 11794
rect 8490 11774 8495 11794
rect 8522 11774 8542 11794
rect 8542 11774 8556 11794
rect 8556 11774 8578 11794
rect 8605 11774 8608 11794
rect 8608 11774 8661 11794
rect 8439 11760 8495 11774
rect 8522 11760 8578 11774
rect 8605 11760 8661 11774
rect 8439 11738 8490 11760
rect 8490 11738 8495 11760
rect 8522 11738 8542 11760
rect 8542 11738 8556 11760
rect 8556 11738 8578 11760
rect 8605 11738 8608 11760
rect 8608 11738 8661 11760
rect 8688 11738 8744 11794
rect 8771 11738 8827 11794
rect 8854 11738 8910 11794
rect 8937 11738 8993 11794
rect 9020 11774 9044 11794
rect 9044 11774 9076 11794
rect 9103 11774 9110 11794
rect 9110 11774 9159 11794
rect 9020 11760 9076 11774
rect 9103 11760 9159 11774
rect 9020 11738 9044 11760
rect 9044 11738 9076 11760
rect 9103 11738 9110 11760
rect 9110 11738 9159 11760
rect 9186 11738 9242 11794
rect 9269 11738 9325 11794
rect 9352 11738 9408 11794
rect 9435 11738 9491 11794
rect 9518 11738 9574 11794
rect 9601 11774 9650 11794
rect 9650 11774 9657 11794
rect 9684 11774 9716 11794
rect 9716 11774 9740 11794
rect 9601 11760 9657 11774
rect 9684 11760 9740 11774
rect 9601 11738 9650 11760
rect 9650 11738 9657 11760
rect 9684 11738 9716 11760
rect 9716 11738 9740 11760
rect 9767 11738 9823 11794
rect 7691 11650 7747 11706
rect 7775 11650 7831 11706
rect 7858 11650 7914 11706
rect 7941 11694 7997 11706
rect 8024 11694 8080 11706
rect 7941 11650 7988 11694
rect 7988 11650 7997 11694
rect 8024 11650 8054 11694
rect 8054 11650 8080 11694
rect 8107 11650 8163 11706
rect 8190 11650 8246 11706
rect 8273 11650 8329 11706
rect 8356 11650 8412 11706
rect 8439 11694 8495 11706
rect 8522 11694 8578 11706
rect 8605 11694 8661 11706
rect 8439 11650 8490 11694
rect 8490 11650 8495 11694
rect 8522 11650 8542 11694
rect 8542 11650 8556 11694
rect 8556 11650 8578 11694
rect 8605 11650 8608 11694
rect 8608 11650 8661 11694
rect 8688 11650 8744 11706
rect 8771 11650 8827 11706
rect 8854 11650 8910 11706
rect 8937 11650 8993 11706
rect 9020 11694 9076 11706
rect 9103 11694 9159 11706
rect 9020 11650 9044 11694
rect 9044 11650 9076 11694
rect 9103 11650 9110 11694
rect 9110 11650 9159 11694
rect 9186 11650 9242 11706
rect 9269 11650 9325 11706
rect 9352 11650 9408 11706
rect 9435 11650 9491 11706
rect 9518 11650 9574 11706
rect 9601 11694 9657 11706
rect 9684 11694 9740 11706
rect 9601 11650 9650 11694
rect 9650 11650 9657 11694
rect 9684 11650 9716 11694
rect 9716 11650 9740 11694
rect 9767 11650 9823 11706
rect 7691 11562 7747 11618
rect 7775 11562 7831 11618
rect 7858 11562 7914 11618
rect 7941 11576 7988 11618
rect 7988 11576 7997 11618
rect 8024 11576 8054 11618
rect 8054 11576 8080 11618
rect 7941 11562 7997 11576
rect 8024 11562 8080 11576
rect 8107 11562 8163 11618
rect 8190 11562 8246 11618
rect 8273 11562 8329 11618
rect 8356 11562 8412 11618
rect 8439 11576 8490 11618
rect 8490 11576 8495 11618
rect 8522 11576 8542 11618
rect 8542 11576 8556 11618
rect 8556 11576 8578 11618
rect 8605 11576 8608 11618
rect 8608 11576 8661 11618
rect 8439 11562 8495 11576
rect 8522 11562 8578 11576
rect 8605 11562 8661 11576
rect 8688 11562 8744 11618
rect 8771 11562 8827 11618
rect 8854 11562 8910 11618
rect 8937 11562 8993 11618
rect 9020 11576 9044 11618
rect 9044 11576 9076 11618
rect 9103 11576 9110 11618
rect 9110 11576 9159 11618
rect 9020 11562 9076 11576
rect 9103 11562 9159 11576
rect 9186 11562 9242 11618
rect 9269 11562 9325 11618
rect 9352 11562 9408 11618
rect 9435 11562 9491 11618
rect 9518 11562 9574 11618
rect 9601 11576 9650 11618
rect 9650 11576 9657 11618
rect 9684 11576 9716 11618
rect 9716 11576 9740 11618
rect 9601 11562 9657 11576
rect 9684 11562 9740 11576
rect 9767 11562 9823 11618
rect 7691 11474 7747 11530
rect 7775 11474 7831 11530
rect 7858 11474 7914 11530
rect 7941 11510 7988 11530
rect 7988 11510 7997 11530
rect 8024 11510 8054 11530
rect 8054 11510 8080 11530
rect 7941 11495 7997 11510
rect 8024 11495 8080 11510
rect 7941 11474 7988 11495
rect 7988 11474 7997 11495
rect 8024 11474 8054 11495
rect 8054 11474 8080 11495
rect 8107 11474 8163 11530
rect 8190 11474 8246 11530
rect 8273 11474 8329 11530
rect 8356 11474 8412 11530
rect 8439 11510 8490 11530
rect 8490 11510 8495 11530
rect 8522 11510 8542 11530
rect 8542 11510 8556 11530
rect 8556 11510 8578 11530
rect 8605 11510 8608 11530
rect 8608 11510 8661 11530
rect 8439 11495 8495 11510
rect 8522 11495 8578 11510
rect 8605 11495 8661 11510
rect 8439 11474 8490 11495
rect 8490 11474 8495 11495
rect 8522 11474 8542 11495
rect 8542 11474 8556 11495
rect 8556 11474 8578 11495
rect 8605 11474 8608 11495
rect 8608 11474 8661 11495
rect 8688 11474 8744 11530
rect 8771 11474 8827 11530
rect 8854 11474 8910 11530
rect 8937 11474 8993 11530
rect 9020 11510 9044 11530
rect 9044 11510 9076 11530
rect 9103 11510 9110 11530
rect 9110 11510 9159 11530
rect 9020 11495 9076 11510
rect 9103 11495 9159 11510
rect 9020 11474 9044 11495
rect 9044 11474 9076 11495
rect 9103 11474 9110 11495
rect 9110 11474 9159 11495
rect 9186 11474 9242 11530
rect 9269 11474 9325 11530
rect 9352 11474 9408 11530
rect 9435 11474 9491 11530
rect 9518 11474 9574 11530
rect 9601 11510 9650 11530
rect 9650 11510 9657 11530
rect 9684 11510 9716 11530
rect 9716 11510 9740 11530
rect 9601 11495 9657 11510
rect 9684 11495 9740 11510
rect 9601 11474 9650 11495
rect 9650 11474 9657 11495
rect 9684 11474 9716 11495
rect 9716 11474 9740 11495
rect 9767 11474 9823 11530
rect 7691 11386 7747 11442
rect 7775 11386 7831 11442
rect 7858 11386 7914 11442
rect 7941 11428 7997 11442
rect 8024 11428 8080 11442
rect 7941 11386 7988 11428
rect 7988 11386 7997 11428
rect 8024 11386 8054 11428
rect 8054 11386 8080 11428
rect 8107 11386 8163 11442
rect 8190 11386 8246 11442
rect 8273 11386 8329 11442
rect 8356 11386 8412 11442
rect 8439 11428 8495 11442
rect 8522 11428 8578 11442
rect 8605 11428 8661 11442
rect 8439 11386 8490 11428
rect 8490 11386 8495 11428
rect 8522 11386 8542 11428
rect 8542 11386 8556 11428
rect 8556 11386 8578 11428
rect 8605 11386 8608 11428
rect 8608 11386 8661 11428
rect 8688 11386 8744 11442
rect 8771 11386 8827 11442
rect 8854 11386 8910 11442
rect 8937 11386 8993 11442
rect 9020 11428 9076 11442
rect 9103 11428 9159 11442
rect 9020 11386 9044 11428
rect 9044 11386 9076 11428
rect 9103 11386 9110 11428
rect 9110 11386 9159 11428
rect 9186 11386 9242 11442
rect 9269 11386 9325 11442
rect 9352 11386 9408 11442
rect 9435 11386 9491 11442
rect 9518 11386 9574 11442
rect 9601 11428 9657 11442
rect 9684 11428 9740 11442
rect 9601 11386 9650 11428
rect 9650 11386 9657 11428
rect 9684 11386 9716 11428
rect 9716 11386 9740 11428
rect 9767 11386 9823 11442
rect 7691 9821 7747 9877
rect 7775 9821 7831 9877
rect 7858 9821 7914 9877
rect 7941 9844 7988 9877
rect 7988 9844 7997 9877
rect 8024 9844 8054 9877
rect 8054 9844 8080 9877
rect 7941 9830 7997 9844
rect 8024 9830 8080 9844
rect 7941 9821 7988 9830
rect 7988 9821 7997 9830
rect 8024 9821 8054 9830
rect 8054 9821 8080 9830
rect 8107 9821 8163 9877
rect 8190 9821 8246 9877
rect 8273 9821 8329 9877
rect 8356 9821 8412 9877
rect 8439 9844 8490 9877
rect 8490 9844 8495 9877
rect 8522 9844 8542 9877
rect 8542 9844 8556 9877
rect 8556 9844 8578 9877
rect 8605 9844 8608 9877
rect 8608 9844 8661 9877
rect 8439 9830 8495 9844
rect 8522 9830 8578 9844
rect 8605 9830 8661 9844
rect 8439 9821 8490 9830
rect 8490 9821 8495 9830
rect 8522 9821 8542 9830
rect 8542 9821 8556 9830
rect 8556 9821 8578 9830
rect 8605 9821 8608 9830
rect 8608 9821 8661 9830
rect 8688 9821 8744 9877
rect 8771 9821 8827 9877
rect 8854 9821 8910 9877
rect 8937 9821 8993 9877
rect 9020 9844 9044 9877
rect 9044 9844 9076 9877
rect 9103 9844 9110 9877
rect 9110 9844 9159 9877
rect 9020 9830 9076 9844
rect 9103 9830 9159 9844
rect 9020 9821 9044 9830
rect 9044 9821 9076 9830
rect 9103 9821 9110 9830
rect 9110 9821 9159 9830
rect 9186 9821 9242 9877
rect 9269 9821 9325 9877
rect 9352 9821 9408 9877
rect 9435 9821 9491 9877
rect 9518 9821 9574 9877
rect 9601 9844 9650 9877
rect 9650 9844 9657 9877
rect 9684 9844 9716 9877
rect 9716 9844 9740 9877
rect 9601 9830 9657 9844
rect 9684 9830 9740 9844
rect 9601 9821 9650 9830
rect 9650 9821 9657 9830
rect 9684 9821 9716 9830
rect 9716 9821 9740 9830
rect 9767 9821 9823 9877
rect 7691 9733 7747 9789
rect 7775 9733 7831 9789
rect 7858 9733 7914 9789
rect 7941 9778 7988 9789
rect 7988 9778 7997 9789
rect 8024 9778 8054 9789
rect 8054 9778 8080 9789
rect 7941 9764 7997 9778
rect 8024 9764 8080 9778
rect 7941 9733 7988 9764
rect 7988 9733 7997 9764
rect 8024 9733 8054 9764
rect 8054 9733 8080 9764
rect 8107 9733 8163 9789
rect 8190 9733 8246 9789
rect 8273 9733 8329 9789
rect 8356 9733 8412 9789
rect 8439 9778 8490 9789
rect 8490 9778 8495 9789
rect 8522 9778 8542 9789
rect 8542 9778 8556 9789
rect 8556 9778 8578 9789
rect 8605 9778 8608 9789
rect 8608 9778 8661 9789
rect 8439 9764 8495 9778
rect 8522 9764 8578 9778
rect 8605 9764 8661 9778
rect 8439 9733 8490 9764
rect 8490 9733 8495 9764
rect 8522 9733 8542 9764
rect 8542 9733 8556 9764
rect 8556 9733 8578 9764
rect 8605 9733 8608 9764
rect 8608 9733 8661 9764
rect 8688 9733 8744 9789
rect 8771 9733 8827 9789
rect 8854 9733 8910 9789
rect 8937 9733 8993 9789
rect 9020 9778 9044 9789
rect 9044 9778 9076 9789
rect 9103 9778 9110 9789
rect 9110 9778 9159 9789
rect 9020 9764 9076 9778
rect 9103 9764 9159 9778
rect 9020 9733 9044 9764
rect 9044 9733 9076 9764
rect 9103 9733 9110 9764
rect 9110 9733 9159 9764
rect 9186 9733 9242 9789
rect 9269 9733 9325 9789
rect 9352 9733 9408 9789
rect 9435 9733 9491 9789
rect 9518 9733 9574 9789
rect 9601 9778 9650 9789
rect 9650 9778 9657 9789
rect 9684 9778 9716 9789
rect 9716 9778 9740 9789
rect 9601 9764 9657 9778
rect 9684 9764 9740 9778
rect 9601 9733 9650 9764
rect 9650 9733 9657 9764
rect 9684 9733 9716 9764
rect 9716 9733 9740 9764
rect 9767 9733 9823 9789
rect 7691 9645 7747 9701
rect 7775 9645 7831 9701
rect 7858 9645 7914 9701
rect 7941 9698 7997 9701
rect 8024 9698 8080 9701
rect 7941 9646 7988 9698
rect 7988 9646 7997 9698
rect 8024 9646 8054 9698
rect 8054 9646 8080 9698
rect 7941 9645 7997 9646
rect 8024 9645 8080 9646
rect 8107 9645 8163 9701
rect 8190 9645 8246 9701
rect 8273 9645 8329 9701
rect 8356 9645 8412 9701
rect 8439 9698 8495 9701
rect 8522 9698 8578 9701
rect 8605 9698 8661 9701
rect 8439 9646 8490 9698
rect 8490 9646 8495 9698
rect 8522 9646 8542 9698
rect 8542 9646 8556 9698
rect 8556 9646 8578 9698
rect 8605 9646 8608 9698
rect 8608 9646 8661 9698
rect 8439 9645 8495 9646
rect 8522 9645 8578 9646
rect 8605 9645 8661 9646
rect 8688 9645 8744 9701
rect 8771 9645 8827 9701
rect 8854 9645 8910 9701
rect 8937 9645 8993 9701
rect 9020 9698 9076 9701
rect 9103 9698 9159 9701
rect 9020 9646 9044 9698
rect 9044 9646 9076 9698
rect 9103 9646 9110 9698
rect 9110 9646 9159 9698
rect 9020 9645 9076 9646
rect 9103 9645 9159 9646
rect 9186 9645 9242 9701
rect 9269 9645 9325 9701
rect 9352 9645 9408 9701
rect 9435 9645 9491 9701
rect 9518 9645 9574 9701
rect 9601 9698 9657 9701
rect 9684 9698 9740 9701
rect 9601 9646 9650 9698
rect 9650 9646 9657 9698
rect 9684 9646 9716 9698
rect 9716 9646 9740 9698
rect 9601 9645 9657 9646
rect 9684 9645 9740 9646
rect 9767 9645 9823 9701
rect 7691 9557 7747 9613
rect 7775 9557 7831 9613
rect 7858 9557 7914 9613
rect 7941 9580 7988 9613
rect 7988 9580 7997 9613
rect 8024 9580 8054 9613
rect 8054 9580 8080 9613
rect 7941 9566 7997 9580
rect 8024 9566 8080 9580
rect 7941 9557 7988 9566
rect 7988 9557 7997 9566
rect 8024 9557 8054 9566
rect 8054 9557 8080 9566
rect 8107 9557 8163 9613
rect 8190 9557 8246 9613
rect 8273 9557 8329 9613
rect 8356 9557 8412 9613
rect 8439 9580 8490 9613
rect 8490 9580 8495 9613
rect 8522 9580 8542 9613
rect 8542 9580 8556 9613
rect 8556 9580 8578 9613
rect 8605 9580 8608 9613
rect 8608 9580 8661 9613
rect 8439 9566 8495 9580
rect 8522 9566 8578 9580
rect 8605 9566 8661 9580
rect 8439 9557 8490 9566
rect 8490 9557 8495 9566
rect 8522 9557 8542 9566
rect 8542 9557 8556 9566
rect 8556 9557 8578 9566
rect 8605 9557 8608 9566
rect 8608 9557 8661 9566
rect 8688 9557 8744 9613
rect 8771 9557 8827 9613
rect 8854 9557 8910 9613
rect 8937 9557 8993 9613
rect 9020 9580 9044 9613
rect 9044 9580 9076 9613
rect 9103 9580 9110 9613
rect 9110 9580 9159 9613
rect 9020 9566 9076 9580
rect 9103 9566 9159 9580
rect 9020 9557 9044 9566
rect 9044 9557 9076 9566
rect 9103 9557 9110 9566
rect 9110 9557 9159 9566
rect 9186 9557 9242 9613
rect 9269 9557 9325 9613
rect 9352 9557 9408 9613
rect 9435 9557 9491 9613
rect 9518 9557 9574 9613
rect 9601 9580 9650 9613
rect 9650 9580 9657 9613
rect 9684 9580 9716 9613
rect 9716 9580 9740 9613
rect 9601 9566 9657 9580
rect 9684 9566 9740 9580
rect 9601 9557 9650 9566
rect 9650 9557 9657 9566
rect 9684 9557 9716 9566
rect 9716 9557 9740 9566
rect 9767 9557 9823 9613
rect 7691 9469 7747 9525
rect 7775 9469 7831 9525
rect 7858 9469 7914 9525
rect 7941 9514 7988 9525
rect 7988 9514 7997 9525
rect 8024 9514 8054 9525
rect 8054 9514 8080 9525
rect 7941 9499 7997 9514
rect 8024 9499 8080 9514
rect 7941 9469 7988 9499
rect 7988 9469 7997 9499
rect 8024 9469 8054 9499
rect 8054 9469 8080 9499
rect 8107 9469 8163 9525
rect 8190 9469 8246 9525
rect 8273 9469 8329 9525
rect 8356 9469 8412 9525
rect 8439 9514 8490 9525
rect 8490 9514 8495 9525
rect 8522 9514 8542 9525
rect 8542 9514 8556 9525
rect 8556 9514 8578 9525
rect 8605 9514 8608 9525
rect 8608 9514 8661 9525
rect 8439 9499 8495 9514
rect 8522 9499 8578 9514
rect 8605 9499 8661 9514
rect 8439 9469 8490 9499
rect 8490 9469 8495 9499
rect 8522 9469 8542 9499
rect 8542 9469 8556 9499
rect 8556 9469 8578 9499
rect 8605 9469 8608 9499
rect 8608 9469 8661 9499
rect 8688 9469 8744 9525
rect 8771 9469 8827 9525
rect 8854 9469 8910 9525
rect 8937 9469 8993 9525
rect 9020 9514 9044 9525
rect 9044 9514 9076 9525
rect 9103 9514 9110 9525
rect 9110 9514 9159 9525
rect 9020 9499 9076 9514
rect 9103 9499 9159 9514
rect 9020 9469 9044 9499
rect 9044 9469 9076 9499
rect 9103 9469 9110 9499
rect 9110 9469 9159 9499
rect 9186 9469 9242 9525
rect 9269 9469 9325 9525
rect 9352 9469 9408 9525
rect 9435 9469 9491 9525
rect 9518 9469 9574 9525
rect 9601 9514 9650 9525
rect 9650 9514 9657 9525
rect 9684 9514 9716 9525
rect 9716 9514 9740 9525
rect 9601 9499 9657 9514
rect 9684 9499 9740 9514
rect 9601 9469 9650 9499
rect 9650 9469 9657 9499
rect 9684 9469 9716 9499
rect 9716 9469 9740 9499
rect 9767 9469 9823 9525
rect 7691 9381 7747 9437
rect 7775 9381 7831 9437
rect 7858 9381 7914 9437
rect 7941 9432 7997 9437
rect 8024 9432 8080 9437
rect 7941 9381 7988 9432
rect 7988 9381 7997 9432
rect 8024 9381 8054 9432
rect 8054 9381 8080 9432
rect 8107 9381 8163 9437
rect 8190 9381 8246 9437
rect 8273 9381 8329 9437
rect 8356 9381 8412 9437
rect 8439 9432 8495 9437
rect 8522 9432 8578 9437
rect 8605 9432 8661 9437
rect 8439 9381 8490 9432
rect 8490 9381 8495 9432
rect 8522 9381 8542 9432
rect 8542 9381 8556 9432
rect 8556 9381 8578 9432
rect 8605 9381 8608 9432
rect 8608 9381 8661 9432
rect 8688 9381 8744 9437
rect 8771 9381 8827 9437
rect 8854 9381 8910 9437
rect 8937 9381 8993 9437
rect 9020 9432 9076 9437
rect 9103 9432 9159 9437
rect 9020 9381 9044 9432
rect 9044 9381 9076 9432
rect 9103 9381 9110 9432
rect 9110 9381 9159 9432
rect 9186 9381 9242 9437
rect 9269 9381 9325 9437
rect 9352 9381 9408 9437
rect 9435 9381 9491 9437
rect 9518 9381 9574 9437
rect 9601 9432 9657 9437
rect 9684 9432 9740 9437
rect 9601 9381 9650 9432
rect 9650 9381 9657 9432
rect 9684 9381 9716 9432
rect 9716 9381 9740 9432
rect 9767 9381 9823 9437
rect 7691 7826 7747 7882
rect 7775 7826 7831 7882
rect 7858 7826 7914 7882
rect 7941 7840 7988 7882
rect 7988 7840 7997 7882
rect 8024 7840 8054 7882
rect 8054 7840 8080 7882
rect 7941 7826 7997 7840
rect 8024 7826 8080 7840
rect 8107 7826 8163 7882
rect 8190 7826 8246 7882
rect 8273 7826 8329 7882
rect 8356 7826 8412 7882
rect 8439 7840 8490 7882
rect 8490 7840 8495 7882
rect 8522 7840 8542 7882
rect 8542 7840 8556 7882
rect 8556 7840 8578 7882
rect 8605 7840 8608 7882
rect 8608 7840 8661 7882
rect 8439 7826 8495 7840
rect 8522 7826 8578 7840
rect 8605 7826 8661 7840
rect 8688 7826 8744 7882
rect 8771 7826 8827 7882
rect 8854 7826 8910 7882
rect 8937 7826 8993 7882
rect 9020 7840 9044 7882
rect 9044 7840 9076 7882
rect 9103 7840 9110 7882
rect 9110 7840 9159 7882
rect 9020 7826 9076 7840
rect 9103 7826 9159 7840
rect 9186 7826 9242 7882
rect 9269 7826 9325 7882
rect 9352 7826 9408 7882
rect 9435 7826 9491 7882
rect 9518 7826 9574 7882
rect 9601 7840 9650 7882
rect 9650 7840 9657 7882
rect 9684 7840 9716 7882
rect 9716 7840 9740 7882
rect 9601 7826 9657 7840
rect 9684 7826 9740 7840
rect 9767 7826 9823 7882
rect 7691 7738 7747 7794
rect 7775 7738 7831 7794
rect 7858 7738 7914 7794
rect 7941 7774 7988 7794
rect 7988 7774 7997 7794
rect 8024 7774 8054 7794
rect 8054 7774 8080 7794
rect 7941 7760 7997 7774
rect 8024 7760 8080 7774
rect 7941 7738 7988 7760
rect 7988 7738 7997 7760
rect 8024 7738 8054 7760
rect 8054 7738 8080 7760
rect 8107 7738 8163 7794
rect 8190 7738 8246 7794
rect 8273 7738 8329 7794
rect 8356 7738 8412 7794
rect 8439 7774 8490 7794
rect 8490 7774 8495 7794
rect 8522 7774 8542 7794
rect 8542 7774 8556 7794
rect 8556 7774 8578 7794
rect 8605 7774 8608 7794
rect 8608 7774 8661 7794
rect 8439 7760 8495 7774
rect 8522 7760 8578 7774
rect 8605 7760 8661 7774
rect 8439 7738 8490 7760
rect 8490 7738 8495 7760
rect 8522 7738 8542 7760
rect 8542 7738 8556 7760
rect 8556 7738 8578 7760
rect 8605 7738 8608 7760
rect 8608 7738 8661 7760
rect 8688 7738 8744 7794
rect 8771 7738 8827 7794
rect 8854 7738 8910 7794
rect 8937 7738 8993 7794
rect 9020 7774 9044 7794
rect 9044 7774 9076 7794
rect 9103 7774 9110 7794
rect 9110 7774 9159 7794
rect 9020 7760 9076 7774
rect 9103 7760 9159 7774
rect 9020 7738 9044 7760
rect 9044 7738 9076 7760
rect 9103 7738 9110 7760
rect 9110 7738 9159 7760
rect 9186 7738 9242 7794
rect 9269 7738 9325 7794
rect 9352 7738 9408 7794
rect 9435 7738 9491 7794
rect 9518 7738 9574 7794
rect 9601 7774 9650 7794
rect 9650 7774 9657 7794
rect 9684 7774 9716 7794
rect 9716 7774 9740 7794
rect 9601 7760 9657 7774
rect 9684 7760 9740 7774
rect 9601 7738 9650 7760
rect 9650 7738 9657 7760
rect 9684 7738 9716 7760
rect 9716 7738 9740 7760
rect 9767 7738 9823 7794
rect 7691 7650 7747 7706
rect 7775 7650 7831 7706
rect 7858 7650 7914 7706
rect 7941 7694 7997 7706
rect 8024 7694 8080 7706
rect 7941 7650 7988 7694
rect 7988 7650 7997 7694
rect 8024 7650 8054 7694
rect 8054 7650 8080 7694
rect 8107 7650 8163 7706
rect 8190 7650 8246 7706
rect 8273 7650 8329 7706
rect 8356 7650 8412 7706
rect 8439 7694 8495 7706
rect 8522 7694 8578 7706
rect 8605 7694 8661 7706
rect 8439 7650 8490 7694
rect 8490 7650 8495 7694
rect 8522 7650 8542 7694
rect 8542 7650 8556 7694
rect 8556 7650 8578 7694
rect 8605 7650 8608 7694
rect 8608 7650 8661 7694
rect 8688 7650 8744 7706
rect 8771 7650 8827 7706
rect 8854 7650 8910 7706
rect 8937 7650 8993 7706
rect 9020 7694 9076 7706
rect 9103 7694 9159 7706
rect 9020 7650 9044 7694
rect 9044 7650 9076 7694
rect 9103 7650 9110 7694
rect 9110 7650 9159 7694
rect 9186 7650 9242 7706
rect 9269 7650 9325 7706
rect 9352 7650 9408 7706
rect 9435 7650 9491 7706
rect 9518 7650 9574 7706
rect 9601 7694 9657 7706
rect 9684 7694 9740 7706
rect 9601 7650 9650 7694
rect 9650 7650 9657 7694
rect 9684 7650 9716 7694
rect 9716 7650 9740 7694
rect 9767 7650 9823 7706
rect 7691 7562 7747 7618
rect 7775 7562 7831 7618
rect 7858 7562 7914 7618
rect 7941 7576 7988 7618
rect 7988 7576 7997 7618
rect 8024 7576 8054 7618
rect 8054 7576 8080 7618
rect 7941 7562 7997 7576
rect 8024 7562 8080 7576
rect 8107 7562 8163 7618
rect 8190 7562 8246 7618
rect 8273 7562 8329 7618
rect 8356 7562 8412 7618
rect 8439 7576 8490 7618
rect 8490 7576 8495 7618
rect 8522 7576 8542 7618
rect 8542 7576 8556 7618
rect 8556 7576 8578 7618
rect 8605 7576 8608 7618
rect 8608 7576 8661 7618
rect 8439 7562 8495 7576
rect 8522 7562 8578 7576
rect 8605 7562 8661 7576
rect 8688 7562 8744 7618
rect 8771 7562 8827 7618
rect 8854 7562 8910 7618
rect 8937 7562 8993 7618
rect 9020 7576 9044 7618
rect 9044 7576 9076 7618
rect 9103 7576 9110 7618
rect 9110 7576 9159 7618
rect 9020 7562 9076 7576
rect 9103 7562 9159 7576
rect 9186 7562 9242 7618
rect 9269 7562 9325 7618
rect 9352 7562 9408 7618
rect 9435 7562 9491 7618
rect 9518 7562 9574 7618
rect 9601 7576 9650 7618
rect 9650 7576 9657 7618
rect 9684 7576 9716 7618
rect 9716 7576 9740 7618
rect 9601 7562 9657 7576
rect 9684 7562 9740 7576
rect 9767 7562 9823 7618
rect 7691 7474 7747 7530
rect 7775 7474 7831 7530
rect 7858 7474 7914 7530
rect 7941 7510 7988 7530
rect 7988 7510 7997 7530
rect 8024 7510 8054 7530
rect 8054 7510 8080 7530
rect 7941 7495 7997 7510
rect 8024 7495 8080 7510
rect 7941 7474 7988 7495
rect 7988 7474 7997 7495
rect 8024 7474 8054 7495
rect 8054 7474 8080 7495
rect 8107 7474 8163 7530
rect 8190 7474 8246 7530
rect 8273 7474 8329 7530
rect 8356 7474 8412 7530
rect 8439 7510 8490 7530
rect 8490 7510 8495 7530
rect 8522 7510 8542 7530
rect 8542 7510 8556 7530
rect 8556 7510 8578 7530
rect 8605 7510 8608 7530
rect 8608 7510 8661 7530
rect 8439 7495 8495 7510
rect 8522 7495 8578 7510
rect 8605 7495 8661 7510
rect 8439 7474 8490 7495
rect 8490 7474 8495 7495
rect 8522 7474 8542 7495
rect 8542 7474 8556 7495
rect 8556 7474 8578 7495
rect 8605 7474 8608 7495
rect 8608 7474 8661 7495
rect 8688 7474 8744 7530
rect 8771 7474 8827 7530
rect 8854 7474 8910 7530
rect 8937 7474 8993 7530
rect 9020 7510 9044 7530
rect 9044 7510 9076 7530
rect 9103 7510 9110 7530
rect 9110 7510 9159 7530
rect 9020 7495 9076 7510
rect 9103 7495 9159 7510
rect 9020 7474 9044 7495
rect 9044 7474 9076 7495
rect 9103 7474 9110 7495
rect 9110 7474 9159 7495
rect 9186 7474 9242 7530
rect 9269 7474 9325 7530
rect 9352 7474 9408 7530
rect 9435 7474 9491 7530
rect 9518 7474 9574 7530
rect 9601 7510 9650 7530
rect 9650 7510 9657 7530
rect 9684 7510 9716 7530
rect 9716 7510 9740 7530
rect 9601 7495 9657 7510
rect 9684 7495 9740 7510
rect 9601 7474 9650 7495
rect 9650 7474 9657 7495
rect 9684 7474 9716 7495
rect 9716 7474 9740 7495
rect 9767 7474 9823 7530
rect 7691 7386 7747 7442
rect 7775 7386 7831 7442
rect 7858 7386 7914 7442
rect 7941 7428 7997 7442
rect 8024 7428 8080 7442
rect 7941 7386 7988 7428
rect 7988 7386 7997 7428
rect 8024 7386 8054 7428
rect 8054 7386 8080 7428
rect 8107 7386 8163 7442
rect 8190 7386 8246 7442
rect 8273 7386 8329 7442
rect 8356 7386 8412 7442
rect 8439 7428 8495 7442
rect 8522 7428 8578 7442
rect 8605 7428 8661 7442
rect 8439 7386 8490 7428
rect 8490 7386 8495 7428
rect 8522 7386 8542 7428
rect 8542 7386 8556 7428
rect 8556 7386 8578 7428
rect 8605 7386 8608 7428
rect 8608 7386 8661 7428
rect 8688 7386 8744 7442
rect 8771 7386 8827 7442
rect 8854 7386 8910 7442
rect 8937 7386 8993 7442
rect 9020 7428 9076 7442
rect 9103 7428 9159 7442
rect 9020 7386 9044 7428
rect 9044 7386 9076 7428
rect 9103 7386 9110 7428
rect 9110 7386 9159 7428
rect 9186 7386 9242 7442
rect 9269 7386 9325 7442
rect 9352 7386 9408 7442
rect 9435 7386 9491 7442
rect 9518 7386 9574 7442
rect 9601 7428 9657 7442
rect 9684 7428 9740 7442
rect 9601 7386 9650 7428
rect 9650 7386 9657 7428
rect 9684 7386 9716 7428
rect 9716 7386 9740 7428
rect 9767 7386 9823 7442
rect 7691 5821 7747 5877
rect 7775 5821 7831 5877
rect 7858 5821 7914 5877
rect 7941 5844 7988 5877
rect 7988 5844 7997 5877
rect 8024 5844 8054 5877
rect 8054 5844 8080 5877
rect 7941 5830 7997 5844
rect 8024 5830 8080 5844
rect 7941 5821 7988 5830
rect 7988 5821 7997 5830
rect 8024 5821 8054 5830
rect 8054 5821 8080 5830
rect 8107 5821 8163 5877
rect 8190 5821 8246 5877
rect 8273 5821 8329 5877
rect 8356 5821 8412 5877
rect 8439 5844 8490 5877
rect 8490 5844 8495 5877
rect 8522 5844 8542 5877
rect 8542 5844 8556 5877
rect 8556 5844 8578 5877
rect 8605 5844 8608 5877
rect 8608 5844 8661 5877
rect 8439 5830 8495 5844
rect 8522 5830 8578 5844
rect 8605 5830 8661 5844
rect 8439 5821 8490 5830
rect 8490 5821 8495 5830
rect 8522 5821 8542 5830
rect 8542 5821 8556 5830
rect 8556 5821 8578 5830
rect 8605 5821 8608 5830
rect 8608 5821 8661 5830
rect 8688 5821 8744 5877
rect 8771 5821 8827 5877
rect 8854 5821 8910 5877
rect 8937 5821 8993 5877
rect 9020 5844 9044 5877
rect 9044 5844 9076 5877
rect 9103 5844 9110 5877
rect 9110 5844 9159 5877
rect 9020 5830 9076 5844
rect 9103 5830 9159 5844
rect 9020 5821 9044 5830
rect 9044 5821 9076 5830
rect 9103 5821 9110 5830
rect 9110 5821 9159 5830
rect 9186 5821 9242 5877
rect 9269 5821 9325 5877
rect 9352 5821 9408 5877
rect 9435 5821 9491 5877
rect 9518 5821 9574 5877
rect 9601 5844 9650 5877
rect 9650 5844 9657 5877
rect 9684 5844 9716 5877
rect 9716 5844 9740 5877
rect 9601 5830 9657 5844
rect 9684 5830 9740 5844
rect 9601 5821 9650 5830
rect 9650 5821 9657 5830
rect 9684 5821 9716 5830
rect 9716 5821 9740 5830
rect 9767 5821 9823 5877
rect 7691 5733 7747 5789
rect 7775 5733 7831 5789
rect 7858 5733 7914 5789
rect 7941 5778 7988 5789
rect 7988 5778 7997 5789
rect 8024 5778 8054 5789
rect 8054 5778 8080 5789
rect 7941 5764 7997 5778
rect 8024 5764 8080 5778
rect 7941 5733 7988 5764
rect 7988 5733 7997 5764
rect 8024 5733 8054 5764
rect 8054 5733 8080 5764
rect 8107 5733 8163 5789
rect 8190 5733 8246 5789
rect 8273 5733 8329 5789
rect 8356 5733 8412 5789
rect 8439 5778 8490 5789
rect 8490 5778 8495 5789
rect 8522 5778 8542 5789
rect 8542 5778 8556 5789
rect 8556 5778 8578 5789
rect 8605 5778 8608 5789
rect 8608 5778 8661 5789
rect 8439 5764 8495 5778
rect 8522 5764 8578 5778
rect 8605 5764 8661 5778
rect 8439 5733 8490 5764
rect 8490 5733 8495 5764
rect 8522 5733 8542 5764
rect 8542 5733 8556 5764
rect 8556 5733 8578 5764
rect 8605 5733 8608 5764
rect 8608 5733 8661 5764
rect 8688 5733 8744 5789
rect 8771 5733 8827 5789
rect 8854 5733 8910 5789
rect 8937 5733 8993 5789
rect 9020 5778 9044 5789
rect 9044 5778 9076 5789
rect 9103 5778 9110 5789
rect 9110 5778 9159 5789
rect 9020 5764 9076 5778
rect 9103 5764 9159 5778
rect 9020 5733 9044 5764
rect 9044 5733 9076 5764
rect 9103 5733 9110 5764
rect 9110 5733 9159 5764
rect 9186 5733 9242 5789
rect 9269 5733 9325 5789
rect 9352 5733 9408 5789
rect 9435 5733 9491 5789
rect 9518 5733 9574 5789
rect 9601 5778 9650 5789
rect 9650 5778 9657 5789
rect 9684 5778 9716 5789
rect 9716 5778 9740 5789
rect 9601 5764 9657 5778
rect 9684 5764 9740 5778
rect 9601 5733 9650 5764
rect 9650 5733 9657 5764
rect 9684 5733 9716 5764
rect 9716 5733 9740 5764
rect 9767 5733 9823 5789
rect 7691 5645 7747 5701
rect 7775 5645 7831 5701
rect 7858 5645 7914 5701
rect 7941 5698 7997 5701
rect 8024 5698 8080 5701
rect 7941 5646 7988 5698
rect 7988 5646 7997 5698
rect 8024 5646 8054 5698
rect 8054 5646 8080 5698
rect 7941 5645 7997 5646
rect 8024 5645 8080 5646
rect 8107 5645 8163 5701
rect 8190 5645 8246 5701
rect 8273 5645 8329 5701
rect 8356 5645 8412 5701
rect 8439 5698 8495 5701
rect 8522 5698 8578 5701
rect 8605 5698 8661 5701
rect 8439 5646 8490 5698
rect 8490 5646 8495 5698
rect 8522 5646 8542 5698
rect 8542 5646 8556 5698
rect 8556 5646 8578 5698
rect 8605 5646 8608 5698
rect 8608 5646 8661 5698
rect 8439 5645 8495 5646
rect 8522 5645 8578 5646
rect 8605 5645 8661 5646
rect 8688 5645 8744 5701
rect 8771 5645 8827 5701
rect 8854 5645 8910 5701
rect 8937 5645 8993 5701
rect 9020 5698 9076 5701
rect 9103 5698 9159 5701
rect 9020 5646 9044 5698
rect 9044 5646 9076 5698
rect 9103 5646 9110 5698
rect 9110 5646 9159 5698
rect 9020 5645 9076 5646
rect 9103 5645 9159 5646
rect 9186 5645 9242 5701
rect 9269 5645 9325 5701
rect 9352 5645 9408 5701
rect 9435 5645 9491 5701
rect 9518 5645 9574 5701
rect 9601 5698 9657 5701
rect 9684 5698 9740 5701
rect 9601 5646 9650 5698
rect 9650 5646 9657 5698
rect 9684 5646 9716 5698
rect 9716 5646 9740 5698
rect 9601 5645 9657 5646
rect 9684 5645 9740 5646
rect 9767 5645 9823 5701
rect 7691 5557 7747 5613
rect 7775 5557 7831 5613
rect 7858 5557 7914 5613
rect 7941 5580 7988 5613
rect 7988 5580 7997 5613
rect 8024 5580 8054 5613
rect 8054 5580 8080 5613
rect 7941 5566 7997 5580
rect 8024 5566 8080 5580
rect 7941 5557 7988 5566
rect 7988 5557 7997 5566
rect 8024 5557 8054 5566
rect 8054 5557 8080 5566
rect 8107 5557 8163 5613
rect 8190 5557 8246 5613
rect 8273 5557 8329 5613
rect 8356 5557 8412 5613
rect 8439 5580 8490 5613
rect 8490 5580 8495 5613
rect 8522 5580 8542 5613
rect 8542 5580 8556 5613
rect 8556 5580 8578 5613
rect 8605 5580 8608 5613
rect 8608 5580 8661 5613
rect 8439 5566 8495 5580
rect 8522 5566 8578 5580
rect 8605 5566 8661 5580
rect 8439 5557 8490 5566
rect 8490 5557 8495 5566
rect 8522 5557 8542 5566
rect 8542 5557 8556 5566
rect 8556 5557 8578 5566
rect 8605 5557 8608 5566
rect 8608 5557 8661 5566
rect 8688 5557 8744 5613
rect 8771 5557 8827 5613
rect 8854 5557 8910 5613
rect 8937 5557 8993 5613
rect 9020 5580 9044 5613
rect 9044 5580 9076 5613
rect 9103 5580 9110 5613
rect 9110 5580 9159 5613
rect 9020 5566 9076 5580
rect 9103 5566 9159 5580
rect 9020 5557 9044 5566
rect 9044 5557 9076 5566
rect 9103 5557 9110 5566
rect 9110 5557 9159 5566
rect 9186 5557 9242 5613
rect 9269 5557 9325 5613
rect 9352 5557 9408 5613
rect 9435 5557 9491 5613
rect 9518 5557 9574 5613
rect 9601 5580 9650 5613
rect 9650 5580 9657 5613
rect 9684 5580 9716 5613
rect 9716 5580 9740 5613
rect 9601 5566 9657 5580
rect 9684 5566 9740 5580
rect 9601 5557 9650 5566
rect 9650 5557 9657 5566
rect 9684 5557 9716 5566
rect 9716 5557 9740 5566
rect 9767 5557 9823 5613
rect 7691 5469 7747 5525
rect 7775 5469 7831 5525
rect 7858 5469 7914 5525
rect 7941 5514 7988 5525
rect 7988 5514 7997 5525
rect 8024 5514 8054 5525
rect 8054 5514 8080 5525
rect 7941 5499 7997 5514
rect 8024 5499 8080 5514
rect 7941 5469 7988 5499
rect 7988 5469 7997 5499
rect 8024 5469 8054 5499
rect 8054 5469 8080 5499
rect 8107 5469 8163 5525
rect 8190 5469 8246 5525
rect 8273 5469 8329 5525
rect 8356 5469 8412 5525
rect 8439 5514 8490 5525
rect 8490 5514 8495 5525
rect 8522 5514 8542 5525
rect 8542 5514 8556 5525
rect 8556 5514 8578 5525
rect 8605 5514 8608 5525
rect 8608 5514 8661 5525
rect 8439 5499 8495 5514
rect 8522 5499 8578 5514
rect 8605 5499 8661 5514
rect 8439 5469 8490 5499
rect 8490 5469 8495 5499
rect 8522 5469 8542 5499
rect 8542 5469 8556 5499
rect 8556 5469 8578 5499
rect 8605 5469 8608 5499
rect 8608 5469 8661 5499
rect 8688 5469 8744 5525
rect 8771 5469 8827 5525
rect 8854 5469 8910 5525
rect 8937 5469 8993 5525
rect 9020 5514 9044 5525
rect 9044 5514 9076 5525
rect 9103 5514 9110 5525
rect 9110 5514 9159 5525
rect 9020 5499 9076 5514
rect 9103 5499 9159 5514
rect 9020 5469 9044 5499
rect 9044 5469 9076 5499
rect 9103 5469 9110 5499
rect 9110 5469 9159 5499
rect 9186 5469 9242 5525
rect 9269 5469 9325 5525
rect 9352 5469 9408 5525
rect 9435 5469 9491 5525
rect 9518 5469 9574 5525
rect 9601 5514 9650 5525
rect 9650 5514 9657 5525
rect 9684 5514 9716 5525
rect 9716 5514 9740 5525
rect 9601 5499 9657 5514
rect 9684 5499 9740 5514
rect 9601 5469 9650 5499
rect 9650 5469 9657 5499
rect 9684 5469 9716 5499
rect 9716 5469 9740 5499
rect 9767 5469 9823 5525
rect 7691 5381 7747 5437
rect 7775 5381 7831 5437
rect 7858 5381 7914 5437
rect 7941 5432 7997 5437
rect 8024 5432 8080 5437
rect 7941 5381 7988 5432
rect 7988 5381 7997 5432
rect 8024 5381 8054 5432
rect 8054 5381 8080 5432
rect 8107 5381 8163 5437
rect 8190 5381 8246 5437
rect 8273 5381 8329 5437
rect 8356 5381 8412 5437
rect 8439 5432 8495 5437
rect 8522 5432 8578 5437
rect 8605 5432 8661 5437
rect 8439 5381 8490 5432
rect 8490 5381 8495 5432
rect 8522 5381 8542 5432
rect 8542 5381 8556 5432
rect 8556 5381 8578 5432
rect 8605 5381 8608 5432
rect 8608 5381 8661 5432
rect 8688 5381 8744 5437
rect 8771 5381 8827 5437
rect 8854 5381 8910 5437
rect 8937 5381 8993 5437
rect 9020 5432 9076 5437
rect 9103 5432 9159 5437
rect 9020 5381 9044 5432
rect 9044 5381 9076 5432
rect 9103 5381 9110 5432
rect 9110 5381 9159 5432
rect 9186 5381 9242 5437
rect 9269 5381 9325 5437
rect 9352 5381 9408 5437
rect 9435 5381 9491 5437
rect 9518 5381 9574 5437
rect 9601 5432 9657 5437
rect 9684 5432 9740 5437
rect 9601 5381 9650 5432
rect 9650 5381 9657 5432
rect 9684 5381 9716 5432
rect 9716 5381 9740 5432
rect 9767 5381 9823 5437
rect 5013 5145 5069 5201
rect 5013 5065 5069 5121
rect 5022 4811 5078 4867
rect 5022 4729 5078 4785
rect 5022 4646 5078 4702
rect 5212 4168 5261 4220
rect 5261 4168 5268 4220
rect 5347 4168 5398 4220
rect 5398 4168 5403 4220
rect 5481 4168 5482 4220
rect 5482 4168 5534 4220
rect 5534 4168 5537 4220
rect 5615 4168 5618 4220
rect 5618 4168 5670 4220
rect 5670 4168 5671 4220
rect 5749 4168 5754 4220
rect 5754 4168 5805 4220
rect 5883 4168 5890 4220
rect 5890 4168 5939 4220
rect 5212 4164 5268 4168
rect 5347 4164 5403 4168
rect 5481 4164 5537 4168
rect 5615 4164 5671 4168
rect 5749 4164 5805 4168
rect 5883 4164 5939 4168
rect 5212 4096 5268 4100
rect 5347 4096 5403 4100
rect 5481 4096 5537 4100
rect 5615 4096 5671 4100
rect 5749 4096 5805 4100
rect 5883 4096 5939 4100
rect 5212 4044 5261 4096
rect 5261 4044 5268 4096
rect 5347 4044 5398 4096
rect 5398 4044 5403 4096
rect 5481 4044 5482 4096
rect 5482 4044 5534 4096
rect 5534 4044 5537 4096
rect 5615 4044 5618 4096
rect 5618 4044 5670 4096
rect 5670 4044 5671 4096
rect 5749 4044 5754 4096
rect 5754 4044 5805 4096
rect 5883 4044 5890 4096
rect 5890 4044 5939 4096
rect 7692 4668 7748 4724
rect 7853 4668 7909 4724
rect 8014 4668 8070 4724
rect 8175 4668 8231 4724
rect 8336 4668 8392 4724
rect 8497 4668 8553 4724
rect 8658 4668 8714 4724
rect 8819 4668 8875 4724
rect 8980 4668 9036 4724
rect 9141 4668 9197 4724
rect 9302 4668 9358 4724
rect 9462 4668 9518 4724
rect 9622 4668 9678 4724
rect 9782 4668 9838 4724
rect 7692 4580 7748 4636
rect 7853 4580 7909 4636
rect 8014 4580 8070 4636
rect 8175 4580 8231 4636
rect 8336 4580 8392 4636
rect 8497 4580 8553 4636
rect 8658 4580 8714 4636
rect 8819 4580 8875 4636
rect 8980 4580 9036 4636
rect 9141 4580 9197 4636
rect 9302 4580 9358 4636
rect 9462 4580 9518 4636
rect 9622 4580 9678 4636
rect 9782 4580 9838 4636
<< metal3 >>
rect 3121 37892 5023 37903
rect 3121 37836 3513 37892
rect 3569 37836 3594 37892
rect 3650 37836 3675 37892
rect 3731 37836 3756 37892
rect 3812 37836 3837 37892
rect 3893 37836 3918 37892
rect 3121 37812 3918 37836
rect 3121 37756 3513 37812
rect 3569 37756 3594 37812
rect 3650 37756 3675 37812
rect 3731 37756 3756 37812
rect 3812 37756 3837 37812
rect 3893 37756 3918 37812
rect 3121 37732 3918 37756
rect 3121 37676 3513 37732
rect 3569 37676 3594 37732
rect 3650 37676 3675 37732
rect 3731 37676 3756 37732
rect 3812 37676 3837 37732
rect 3893 37676 3918 37732
rect 3121 37652 3918 37676
rect 3121 37596 3513 37652
rect 3569 37596 3594 37652
rect 3650 37596 3675 37652
rect 3731 37596 3756 37652
rect 3812 37596 3837 37652
rect 3893 37596 3918 37652
rect 3121 37572 3918 37596
rect 3121 37516 3513 37572
rect 3569 37516 3594 37572
rect 3650 37516 3675 37572
rect 3731 37516 3756 37572
rect 3812 37516 3837 37572
rect 3893 37516 3918 37572
rect 3121 37492 3918 37516
rect 3121 37436 3513 37492
rect 3569 37436 3594 37492
rect 3650 37436 3675 37492
rect 3731 37436 3756 37492
rect 3812 37436 3837 37492
rect 3893 37436 3918 37492
rect 3121 37412 3918 37436
rect 3121 37356 3513 37412
rect 3569 37356 3594 37412
rect 3650 37356 3675 37412
rect 3731 37356 3756 37412
rect 3812 37356 3837 37412
rect 3893 37356 3918 37412
rect 3121 37332 3918 37356
rect 3121 37276 3513 37332
rect 3569 37276 3594 37332
rect 3650 37276 3675 37332
rect 3731 37276 3756 37332
rect 3812 37276 3837 37332
rect 3893 37276 3918 37332
rect 3121 37252 3918 37276
rect 3121 37196 3513 37252
rect 3569 37196 3594 37252
rect 3650 37196 3675 37252
rect 3731 37196 3756 37252
rect 3812 37196 3837 37252
rect 3893 37196 3918 37252
rect 3121 37172 3918 37196
rect 3121 37116 3513 37172
rect 3569 37116 3594 37172
rect 3650 37116 3675 37172
rect 3731 37116 3756 37172
rect 3812 37116 3837 37172
rect 3893 37116 3918 37172
rect 3121 37092 3918 37116
rect 3121 37036 3513 37092
rect 3569 37036 3594 37092
rect 3650 37036 3675 37092
rect 3731 37036 3756 37092
rect 3812 37036 3837 37092
rect 3893 37036 3918 37092
rect 5014 37036 5023 37892
rect 3121 35896 5023 37036
rect 3121 35840 3513 35896
rect 3569 35840 3593 35896
rect 3649 35840 3673 35896
rect 3729 35840 3753 35896
rect 3809 35840 3833 35896
rect 3889 35840 3913 35896
rect 3969 35840 3993 35896
rect 4049 35840 4073 35896
rect 4129 35840 4153 35896
rect 4209 35840 4233 35896
rect 4289 35840 4314 35896
rect 4370 35840 4395 35896
rect 4451 35840 4476 35896
rect 4532 35840 4557 35896
rect 4613 35840 4638 35896
rect 4694 35840 4719 35896
rect 4775 35840 4800 35896
rect 4856 35840 4881 35896
rect 4937 35840 4962 35896
rect 5018 35840 5023 35896
rect 3121 35802 5023 35840
rect 3121 35746 3513 35802
rect 3569 35746 3593 35802
rect 3649 35746 3673 35802
rect 3729 35746 3753 35802
rect 3809 35746 3833 35802
rect 3889 35746 3913 35802
rect 3969 35746 3993 35802
rect 4049 35746 4073 35802
rect 4129 35746 4153 35802
rect 4209 35746 4233 35802
rect 4289 35746 4314 35802
rect 4370 35746 4395 35802
rect 4451 35746 4476 35802
rect 4532 35746 4557 35802
rect 4613 35746 4638 35802
rect 4694 35746 4719 35802
rect 4775 35746 4800 35802
rect 4856 35746 4881 35802
rect 4937 35746 4962 35802
rect 5018 35746 5023 35802
rect 3121 35708 5023 35746
rect 3121 35652 3513 35708
rect 3569 35652 3593 35708
rect 3649 35652 3673 35708
rect 3729 35652 3753 35708
rect 3809 35652 3833 35708
rect 3889 35652 3913 35708
rect 3969 35652 3993 35708
rect 4049 35652 4073 35708
rect 4129 35652 4153 35708
rect 4209 35652 4233 35708
rect 4289 35652 4314 35708
rect 4370 35652 4395 35708
rect 4451 35652 4476 35708
rect 4532 35652 4557 35708
rect 4613 35652 4638 35708
rect 4694 35652 4719 35708
rect 4775 35652 4800 35708
rect 4856 35652 4881 35708
rect 4937 35652 4962 35708
rect 5018 35652 5023 35708
rect 3121 35614 5023 35652
rect 3121 35558 3513 35614
rect 3569 35558 3593 35614
rect 3649 35558 3673 35614
rect 3729 35558 3753 35614
rect 3809 35558 3833 35614
rect 3889 35558 3913 35614
rect 3969 35558 3993 35614
rect 4049 35558 4073 35614
rect 4129 35558 4153 35614
rect 4209 35558 4233 35614
rect 4289 35558 4314 35614
rect 4370 35558 4395 35614
rect 4451 35558 4476 35614
rect 4532 35558 4557 35614
rect 4613 35558 4638 35614
rect 4694 35558 4719 35614
rect 4775 35558 4800 35614
rect 4856 35558 4881 35614
rect 4937 35558 4962 35614
rect 5018 35558 5023 35614
rect 3121 35520 5023 35558
rect 3121 35464 3513 35520
rect 3569 35464 3593 35520
rect 3649 35464 3673 35520
rect 3729 35464 3753 35520
rect 3809 35464 3833 35520
rect 3889 35464 3913 35520
rect 3969 35464 3993 35520
rect 4049 35464 4073 35520
rect 4129 35464 4153 35520
rect 4209 35464 4233 35520
rect 4289 35464 4314 35520
rect 4370 35464 4395 35520
rect 4451 35464 4476 35520
rect 4532 35464 4557 35520
rect 4613 35464 4638 35520
rect 4694 35464 4719 35520
rect 4775 35464 4800 35520
rect 4856 35464 4881 35520
rect 4937 35464 4962 35520
rect 5018 35464 5023 35520
rect 3121 35426 5023 35464
rect 3121 35370 3513 35426
rect 3569 35370 3593 35426
rect 3649 35370 3673 35426
rect 3729 35370 3753 35426
rect 3809 35370 3833 35426
rect 3889 35370 3913 35426
rect 3969 35370 3993 35426
rect 4049 35370 4073 35426
rect 4129 35370 4153 35426
rect 4209 35370 4233 35426
rect 4289 35370 4314 35426
rect 4370 35370 4395 35426
rect 4451 35370 4476 35426
rect 4532 35370 4557 35426
rect 4613 35370 4638 35426
rect 4694 35370 4719 35426
rect 4775 35370 4800 35426
rect 4856 35370 4881 35426
rect 4937 35370 4962 35426
rect 5018 35370 5023 35426
rect 100 34197 2580 34239
rect 100 34137 2394 34197
rect 100 34073 2220 34137
rect 2284 34073 2305 34137
rect 2369 34133 2394 34137
rect 2458 34133 2502 34197
rect 2566 34133 2580 34197
rect 2369 34089 2580 34133
rect 2369 34073 2394 34089
rect 100 34051 2394 34073
rect 100 33987 2123 34051
rect 2187 33987 2204 34051
rect 2268 33987 2284 34051
rect 2348 34025 2394 34051
rect 2458 34025 2502 34089
rect 2566 34025 2580 34089
rect 2348 33987 2580 34025
rect 100 33981 2580 33987
rect 100 33933 2394 33981
rect 100 33915 2123 33933
rect 100 33851 1998 33915
rect 2062 33869 2123 33915
rect 2187 33869 2204 33933
rect 2268 33869 2284 33933
rect 2348 33917 2394 33933
rect 2458 33917 2502 33981
rect 2566 33917 2580 33981
rect 2348 33872 2580 33917
rect 2348 33869 2394 33872
rect 2062 33851 2394 33869
rect 100 33818 2394 33851
rect 100 33754 1893 33818
rect 1957 33754 1975 33818
rect 2039 33754 2057 33818
rect 2121 33754 2139 33818
rect 2203 33754 2221 33818
rect 2285 33754 2302 33818
rect 2366 33808 2394 33818
rect 2458 33808 2502 33872
rect 2566 33808 2580 33872
rect 2366 33763 2580 33808
rect 2366 33754 2394 33763
rect 100 33699 2394 33754
rect 2458 33699 2502 33763
rect 2566 33699 2580 33763
rect 100 33683 2580 33699
rect 100 33619 1766 33683
rect 1830 33670 2580 33683
rect 1830 33619 1893 33670
rect 100 33606 1893 33619
rect 1957 33606 1975 33670
rect 2039 33606 2057 33670
rect 2121 33606 2139 33670
rect 2203 33606 2221 33670
rect 2285 33606 2302 33670
rect 2366 33606 2580 33670
rect 100 33572 2580 33606
rect 100 33508 1684 33572
rect 1748 33508 1782 33572
rect 1846 33508 1880 33572
rect 1944 33508 1978 33572
rect 2042 33508 2075 33572
rect 2139 33564 2580 33572
rect 2139 33508 2220 33564
rect 100 33500 2220 33508
rect 2284 33500 2580 33564
rect 100 33468 2580 33500
rect 100 33404 1551 33468
rect 1615 33448 2580 33468
rect 1615 33404 1684 33448
rect 100 33384 1684 33404
rect 1748 33384 1782 33448
rect 1846 33384 1880 33448
rect 1944 33384 1978 33448
rect 2042 33384 2075 33448
rect 2139 33384 2580 33448
rect 100 33366 2580 33384
rect 100 33302 1471 33366
rect 1535 33302 1553 33366
rect 1617 33302 1635 33366
rect 1699 33302 1717 33366
rect 1781 33302 1799 33366
rect 1863 33302 1880 33366
rect 1944 33349 2580 33366
rect 1944 33302 2005 33349
rect 100 33285 2005 33302
rect 2069 33285 2580 33349
rect 100 33229 2580 33285
rect 100 33165 1312 33229
rect 1376 33218 2580 33229
rect 1376 33165 1471 33218
rect 100 33154 1471 33165
rect 1535 33154 1553 33218
rect 1617 33154 1635 33218
rect 1699 33154 1717 33218
rect 1781 33154 1799 33218
rect 1863 33154 1880 33218
rect 1944 33154 2580 33218
rect 100 33138 2580 33154
rect 100 33074 1215 33138
rect 1279 33074 1297 33138
rect 1361 33074 1379 33138
rect 1443 33074 1461 33138
rect 1525 33074 1543 33138
rect 1607 33074 1624 33138
rect 1688 33110 2580 33138
rect 1688 33074 1766 33110
rect 100 33046 1766 33074
rect 1830 33046 2580 33110
rect 100 33006 2580 33046
rect 100 32942 1089 33006
rect 1153 32990 2580 33006
rect 1153 32942 1215 32990
rect 100 32926 1215 32942
rect 1279 32926 1297 32990
rect 1361 32926 1379 32990
rect 1443 32926 1461 32990
rect 1525 32926 1543 32990
rect 1607 32926 1624 32990
rect 1688 32926 2580 32990
rect 100 32908 2580 32926
rect 100 32844 967 32908
rect 1031 32844 1059 32908
rect 1123 32844 1151 32908
rect 1215 32844 1243 32908
rect 1307 32844 1335 32908
rect 1399 32844 1427 32908
rect 1491 32887 2580 32908
rect 1491 32844 1543 32887
rect 100 32828 1543 32844
rect 100 32764 967 32828
rect 1031 32764 1059 32828
rect 1123 32764 1151 32828
rect 1215 32764 1243 32828
rect 1307 32764 1335 32828
rect 1399 32764 1427 32828
rect 1491 32823 1543 32828
rect 1607 32823 2580 32887
rect 1491 32764 2580 32823
rect 100 32748 2580 32764
rect 100 32684 967 32748
rect 1031 32684 1059 32748
rect 1123 32684 1151 32748
rect 1215 32684 1243 32748
rect 1307 32684 1335 32748
rect 1399 32684 1427 32748
rect 1491 32684 2580 32748
rect 100 32668 2580 32684
rect 100 32604 967 32668
rect 1031 32604 1059 32668
rect 1123 32604 1151 32668
rect 1215 32604 1243 32668
rect 1307 32604 1335 32668
rect 1399 32604 1427 32668
rect 1491 32604 2580 32668
rect 100 32588 2580 32604
rect 100 32524 967 32588
rect 1031 32524 1059 32588
rect 1123 32524 1151 32588
rect 1215 32524 1243 32588
rect 1307 32524 1335 32588
rect 1399 32524 1427 32588
rect 1491 32524 2580 32588
rect 100 32508 2580 32524
rect 100 32444 967 32508
rect 1031 32444 1059 32508
rect 1123 32444 1151 32508
rect 1215 32444 1243 32508
rect 1307 32444 1335 32508
rect 1399 32444 1427 32508
rect 1491 32444 2580 32508
rect 100 32428 2580 32444
rect 100 32364 967 32428
rect 1031 32364 1059 32428
rect 1123 32364 1151 32428
rect 1215 32364 1243 32428
rect 1307 32364 1335 32428
rect 1399 32364 1427 32428
rect 1491 32364 2580 32428
rect 100 32348 2580 32364
rect 100 32284 967 32348
rect 1031 32284 1059 32348
rect 1123 32284 1151 32348
rect 1215 32284 1243 32348
rect 1307 32284 1335 32348
rect 1399 32284 1427 32348
rect 1491 32284 2580 32348
rect 100 32268 2580 32284
rect 100 32204 967 32268
rect 1031 32204 1059 32268
rect 1123 32204 1151 32268
rect 1215 32204 1243 32268
rect 1307 32204 1335 32268
rect 1399 32204 1427 32268
rect 1491 32204 2580 32268
rect 100 32188 2580 32204
rect 100 32124 967 32188
rect 1031 32124 1059 32188
rect 1123 32124 1151 32188
rect 1215 32124 1243 32188
rect 1307 32124 1335 32188
rect 1399 32124 1427 32188
rect 1491 32124 2580 32188
rect 100 32108 2580 32124
rect 100 32044 967 32108
rect 1031 32044 1059 32108
rect 1123 32044 1151 32108
rect 1215 32044 1243 32108
rect 1307 32044 1335 32108
rect 1399 32044 1427 32108
rect 1491 32044 2580 32108
rect 100 32028 2580 32044
rect 100 31964 967 32028
rect 1031 31964 1059 32028
rect 1123 31964 1151 32028
rect 1215 31964 1243 32028
rect 1307 31964 1335 32028
rect 1399 31964 1427 32028
rect 1491 31964 2580 32028
rect 100 31948 2580 31964
rect 100 31884 967 31948
rect 1031 31884 1059 31948
rect 1123 31884 1151 31948
rect 1215 31884 1243 31948
rect 1307 31884 1335 31948
rect 1399 31884 1427 31948
rect 1491 31884 2580 31948
rect 100 31868 2580 31884
rect 100 31804 967 31868
rect 1031 31804 1059 31868
rect 1123 31804 1151 31868
rect 1215 31804 1243 31868
rect 1307 31804 1335 31868
rect 1399 31804 1427 31868
rect 1491 31804 2580 31868
rect 100 31788 2580 31804
rect 100 31724 967 31788
rect 1031 31724 1059 31788
rect 1123 31724 1151 31788
rect 1215 31724 1243 31788
rect 1307 31724 1335 31788
rect 1399 31724 1427 31788
rect 1491 31724 2580 31788
rect 100 31708 2580 31724
rect 100 31644 967 31708
rect 1031 31644 1059 31708
rect 1123 31644 1151 31708
rect 1215 31644 1243 31708
rect 1307 31644 1335 31708
rect 1399 31644 1427 31708
rect 1491 31644 2580 31708
rect 100 31628 2580 31644
rect 100 31564 967 31628
rect 1031 31564 1059 31628
rect 1123 31564 1151 31628
rect 1215 31564 1243 31628
rect 1307 31564 1335 31628
rect 1399 31564 1427 31628
rect 1491 31564 2580 31628
rect 100 31548 2580 31564
rect 100 31484 967 31548
rect 1031 31484 1059 31548
rect 1123 31484 1151 31548
rect 1215 31484 1243 31548
rect 1307 31484 1335 31548
rect 1399 31484 1427 31548
rect 1491 31484 2580 31548
rect 100 31468 2580 31484
rect 100 31404 967 31468
rect 1031 31404 1059 31468
rect 1123 31404 1151 31468
rect 1215 31404 1243 31468
rect 1307 31404 1335 31468
rect 1399 31404 1427 31468
rect 1491 31404 2580 31468
rect 100 31388 2580 31404
rect 100 31324 967 31388
rect 1031 31324 1059 31388
rect 1123 31324 1151 31388
rect 1215 31324 1243 31388
rect 1307 31324 1335 31388
rect 1399 31324 1427 31388
rect 1491 31324 2580 31388
rect 100 31308 2580 31324
rect 100 31244 967 31308
rect 1031 31244 1059 31308
rect 1123 31244 1151 31308
rect 1215 31244 1243 31308
rect 1307 31244 1335 31308
rect 1399 31244 1427 31308
rect 1491 31244 2580 31308
rect 100 31228 2580 31244
rect 100 31164 967 31228
rect 1031 31164 1059 31228
rect 1123 31164 1151 31228
rect 1215 31164 1243 31228
rect 1307 31164 1335 31228
rect 1399 31164 1427 31228
rect 1491 31164 2580 31228
rect 100 31148 2580 31164
rect 100 31084 967 31148
rect 1031 31084 1059 31148
rect 1123 31084 1151 31148
rect 1215 31084 1243 31148
rect 1307 31084 1335 31148
rect 1399 31084 1427 31148
rect 1491 31084 2580 31148
rect 100 31068 2580 31084
rect 100 31004 967 31068
rect 1031 31004 1059 31068
rect 1123 31004 1151 31068
rect 1215 31004 1243 31068
rect 1307 31004 1335 31068
rect 1399 31004 1427 31068
rect 1491 31004 2580 31068
rect 100 30988 2580 31004
rect 100 30924 967 30988
rect 1031 30924 1059 30988
rect 1123 30924 1151 30988
rect 1215 30924 1243 30988
rect 1307 30924 1335 30988
rect 1399 30924 1427 30988
rect 1491 30924 2580 30988
rect 100 30908 2580 30924
rect 100 30844 967 30908
rect 1031 30844 1059 30908
rect 1123 30844 1151 30908
rect 1215 30844 1243 30908
rect 1307 30844 1335 30908
rect 1399 30844 1427 30908
rect 1491 30844 2580 30908
rect 100 30828 2580 30844
rect 100 30764 967 30828
rect 1031 30764 1059 30828
rect 1123 30764 1151 30828
rect 1215 30764 1243 30828
rect 1307 30764 1335 30828
rect 1399 30764 1427 30828
rect 1491 30764 2580 30828
rect 100 30748 2580 30764
rect 100 30684 967 30748
rect 1031 30684 1059 30748
rect 1123 30684 1151 30748
rect 1215 30684 1243 30748
rect 1307 30684 1335 30748
rect 1399 30684 1427 30748
rect 1491 30684 2580 30748
rect 100 30668 2580 30684
rect 100 30604 967 30668
rect 1031 30604 1059 30668
rect 1123 30604 1151 30668
rect 1215 30604 1243 30668
rect 1307 30604 1335 30668
rect 1399 30604 1427 30668
rect 1491 30604 2580 30668
rect 100 30588 2580 30604
rect 100 30524 967 30588
rect 1031 30524 1059 30588
rect 1123 30524 1151 30588
rect 1215 30524 1243 30588
rect 1307 30524 1335 30588
rect 1399 30524 1427 30588
rect 1491 30524 2580 30588
rect 100 30508 2580 30524
rect 100 30444 967 30508
rect 1031 30444 1059 30508
rect 1123 30444 1151 30508
rect 1215 30444 1243 30508
rect 1307 30444 1335 30508
rect 1399 30444 1427 30508
rect 1491 30444 2580 30508
rect 100 30428 2580 30444
rect 100 30364 967 30428
rect 1031 30364 1059 30428
rect 1123 30364 1151 30428
rect 1215 30364 1243 30428
rect 1307 30364 1335 30428
rect 1399 30364 1427 30428
rect 1491 30364 2580 30428
rect 100 30348 2580 30364
rect 100 30284 967 30348
rect 1031 30284 1059 30348
rect 1123 30284 1151 30348
rect 1215 30284 1243 30348
rect 1307 30284 1335 30348
rect 1399 30284 1427 30348
rect 1491 30284 2580 30348
rect 100 30268 2580 30284
rect 100 30204 967 30268
rect 1031 30204 1059 30268
rect 1123 30204 1151 30268
rect 1215 30204 1243 30268
rect 1307 30204 1335 30268
rect 1399 30204 1427 30268
rect 1491 30204 2580 30268
rect 100 30188 2580 30204
rect 100 30124 967 30188
rect 1031 30124 1059 30188
rect 1123 30124 1151 30188
rect 1215 30124 1243 30188
rect 1307 30124 1335 30188
rect 1399 30124 1427 30188
rect 1491 30124 2580 30188
rect 100 30108 2580 30124
rect 100 30044 967 30108
rect 1031 30044 1059 30108
rect 1123 30044 1151 30108
rect 1215 30044 1243 30108
rect 1307 30044 1335 30108
rect 1399 30044 1427 30108
rect 1491 30044 2580 30108
rect 100 30028 2580 30044
rect 100 29964 967 30028
rect 1031 29964 1059 30028
rect 1123 29964 1151 30028
rect 1215 29964 1243 30028
rect 1307 29964 1335 30028
rect 1399 29964 1427 30028
rect 1491 29964 2580 30028
rect 100 29948 2580 29964
rect 100 29884 967 29948
rect 1031 29884 1059 29948
rect 1123 29884 1151 29948
rect 1215 29884 1243 29948
rect 1307 29884 1335 29948
rect 1399 29884 1427 29948
rect 1491 29884 2580 29948
rect 100 29868 2580 29884
rect 100 29804 967 29868
rect 1031 29804 1059 29868
rect 1123 29804 1151 29868
rect 1215 29804 1243 29868
rect 1307 29804 1335 29868
rect 1399 29804 1427 29868
rect 1491 29804 2580 29868
rect 100 29788 2580 29804
rect 100 29724 967 29788
rect 1031 29724 1059 29788
rect 1123 29724 1151 29788
rect 1215 29724 1243 29788
rect 1307 29724 1335 29788
rect 1399 29724 1427 29788
rect 1491 29724 2580 29788
rect 100 29708 2580 29724
rect 100 29644 967 29708
rect 1031 29644 1059 29708
rect 1123 29644 1151 29708
rect 1215 29644 1243 29708
rect 1307 29644 1335 29708
rect 1399 29644 1427 29708
rect 1491 29644 2580 29708
rect 100 29628 2580 29644
rect 100 29564 967 29628
rect 1031 29564 1059 29628
rect 1123 29564 1151 29628
rect 1215 29564 1243 29628
rect 1307 29564 1335 29628
rect 1399 29564 1427 29628
rect 1491 29564 2580 29628
rect 100 29548 2580 29564
rect 100 29484 967 29548
rect 1031 29484 1059 29548
rect 1123 29484 1151 29548
rect 1215 29484 1243 29548
rect 1307 29484 1335 29548
rect 1399 29484 1427 29548
rect 1491 29484 2580 29548
rect 100 29468 2580 29484
rect 100 29404 967 29468
rect 1031 29404 1059 29468
rect 1123 29404 1151 29468
rect 1215 29404 1243 29468
rect 1307 29404 1335 29468
rect 1399 29404 1427 29468
rect 1491 29404 2580 29468
rect 100 29388 2580 29404
rect 100 29324 967 29388
rect 1031 29324 1059 29388
rect 1123 29324 1151 29388
rect 1215 29324 1243 29388
rect 1307 29324 1335 29388
rect 1399 29324 1427 29388
rect 1491 29324 2580 29388
rect 100 29308 2580 29324
rect 100 29244 967 29308
rect 1031 29244 1059 29308
rect 1123 29244 1151 29308
rect 1215 29244 1243 29308
rect 1307 29244 1335 29308
rect 1399 29244 1427 29308
rect 1491 29244 2580 29308
rect 100 29228 2580 29244
rect 100 29164 967 29228
rect 1031 29164 1059 29228
rect 1123 29164 1151 29228
rect 1215 29164 1243 29228
rect 1307 29164 1335 29228
rect 1399 29164 1427 29228
rect 1491 29164 2580 29228
rect 100 29148 2580 29164
rect 100 29084 967 29148
rect 1031 29084 1059 29148
rect 1123 29084 1151 29148
rect 1215 29084 1243 29148
rect 1307 29084 1335 29148
rect 1399 29084 1427 29148
rect 1491 29084 2580 29148
rect 100 29068 2580 29084
rect 100 29004 967 29068
rect 1031 29004 1059 29068
rect 1123 29004 1151 29068
rect 1215 29004 1243 29068
rect 1307 29004 1335 29068
rect 1399 29004 1427 29068
rect 1491 29004 2580 29068
rect 100 28988 2580 29004
rect 100 28924 967 28988
rect 1031 28924 1059 28988
rect 1123 28924 1151 28988
rect 1215 28924 1243 28988
rect 1307 28924 1335 28988
rect 1399 28924 1427 28988
rect 1491 28924 2580 28988
rect 100 28908 2580 28924
rect 100 28844 967 28908
rect 1031 28844 1059 28908
rect 1123 28844 1151 28908
rect 1215 28844 1243 28908
rect 1307 28844 1335 28908
rect 1399 28844 1427 28908
rect 1491 28844 2580 28908
rect 100 28828 2580 28844
rect 100 28764 967 28828
rect 1031 28764 1059 28828
rect 1123 28764 1151 28828
rect 1215 28764 1243 28828
rect 1307 28764 1335 28828
rect 1399 28764 1427 28828
rect 1491 28764 2580 28828
rect 100 28748 2580 28764
rect 100 28684 967 28748
rect 1031 28684 1059 28748
rect 1123 28684 1151 28748
rect 1215 28684 1243 28748
rect 1307 28684 1335 28748
rect 1399 28684 1427 28748
rect 1491 28684 2580 28748
rect 100 28668 2580 28684
rect 100 28604 967 28668
rect 1031 28604 1059 28668
rect 1123 28604 1151 28668
rect 1215 28604 1243 28668
rect 1307 28604 1335 28668
rect 1399 28604 1427 28668
rect 1491 28604 2580 28668
rect 100 28588 2580 28604
rect 100 28524 967 28588
rect 1031 28524 1059 28588
rect 1123 28524 1151 28588
rect 1215 28524 1243 28588
rect 1307 28524 1335 28588
rect 1399 28524 1427 28588
rect 1491 28524 2580 28588
rect 100 28508 2580 28524
rect 100 28444 967 28508
rect 1031 28444 1059 28508
rect 1123 28444 1151 28508
rect 1215 28444 1243 28508
rect 1307 28444 1335 28508
rect 1399 28444 1427 28508
rect 1491 28444 2580 28508
rect 100 28428 2580 28444
rect 100 28364 967 28428
rect 1031 28364 1059 28428
rect 1123 28364 1151 28428
rect 1215 28364 1243 28428
rect 1307 28364 1335 28428
rect 1399 28364 1427 28428
rect 1491 28364 2580 28428
rect 100 28348 2580 28364
rect 100 28284 967 28348
rect 1031 28284 1059 28348
rect 1123 28284 1151 28348
rect 1215 28284 1243 28348
rect 1307 28284 1335 28348
rect 1399 28284 1427 28348
rect 1491 28284 2580 28348
rect 100 28268 2580 28284
rect 100 28204 967 28268
rect 1031 28204 1059 28268
rect 1123 28204 1151 28268
rect 1215 28204 1243 28268
rect 1307 28204 1335 28268
rect 1399 28204 1427 28268
rect 1491 28204 2580 28268
rect 100 28188 2580 28204
rect 100 28124 967 28188
rect 1031 28124 1059 28188
rect 1123 28124 1151 28188
rect 1215 28124 1243 28188
rect 1307 28124 1335 28188
rect 1399 28124 1427 28188
rect 1491 28124 2580 28188
rect 100 28108 2580 28124
rect 100 28044 967 28108
rect 1031 28044 1059 28108
rect 1123 28044 1151 28108
rect 1215 28044 1243 28108
rect 1307 28044 1335 28108
rect 1399 28044 1427 28108
rect 1491 28044 2580 28108
rect 100 28028 2580 28044
rect 100 27964 967 28028
rect 1031 27964 1059 28028
rect 1123 27964 1151 28028
rect 1215 27964 1243 28028
rect 1307 27964 1335 28028
rect 1399 27964 1427 28028
rect 1491 27964 2580 28028
rect 100 27948 2580 27964
rect 100 27884 967 27948
rect 1031 27884 1059 27948
rect 1123 27884 1151 27948
rect 1215 27884 1243 27948
rect 1307 27884 1335 27948
rect 1399 27884 1427 27948
rect 1491 27884 2580 27948
rect 100 27868 2580 27884
rect 100 27804 967 27868
rect 1031 27804 1059 27868
rect 1123 27804 1151 27868
rect 1215 27804 1243 27868
rect 1307 27804 1335 27868
rect 1399 27804 1427 27868
rect 1491 27804 2580 27868
rect 100 27788 2580 27804
rect 100 27724 967 27788
rect 1031 27724 1059 27788
rect 1123 27724 1151 27788
rect 1215 27724 1243 27788
rect 1307 27724 1335 27788
rect 1399 27724 1427 27788
rect 1491 27724 2580 27788
rect 100 27708 2580 27724
rect 100 27644 967 27708
rect 1031 27644 1059 27708
rect 1123 27644 1151 27708
rect 1215 27644 1243 27708
rect 1307 27644 1335 27708
rect 1399 27644 1427 27708
rect 1491 27644 2580 27708
rect 100 27628 2580 27644
rect 100 27564 967 27628
rect 1031 27564 1059 27628
rect 1123 27564 1151 27628
rect 1215 27564 1243 27628
rect 1307 27564 1335 27628
rect 1399 27564 1427 27628
rect 1491 27564 2580 27628
rect 100 27548 2580 27564
rect 100 27484 967 27548
rect 1031 27484 1059 27548
rect 1123 27484 1151 27548
rect 1215 27484 1243 27548
rect 1307 27484 1335 27548
rect 1399 27484 1427 27548
rect 1491 27484 2580 27548
rect 100 27468 2580 27484
rect 100 27404 967 27468
rect 1031 27404 1059 27468
rect 1123 27404 1151 27468
rect 1215 27404 1243 27468
rect 1307 27404 1335 27468
rect 1399 27404 1427 27468
rect 1491 27404 2580 27468
rect 100 27388 2580 27404
rect 100 27324 967 27388
rect 1031 27324 1059 27388
rect 1123 27324 1151 27388
rect 1215 27324 1243 27388
rect 1307 27324 1335 27388
rect 1399 27324 1427 27388
rect 1491 27324 2580 27388
rect 100 27308 2580 27324
rect 100 27244 967 27308
rect 1031 27244 1059 27308
rect 1123 27244 1151 27308
rect 1215 27244 1243 27308
rect 1307 27244 1335 27308
rect 1399 27244 1427 27308
rect 1491 27244 2580 27308
rect 100 27228 2580 27244
rect 100 27164 967 27228
rect 1031 27164 1059 27228
rect 1123 27164 1151 27228
rect 1215 27164 1243 27228
rect 1307 27164 1335 27228
rect 1399 27164 1427 27228
rect 1491 27164 2580 27228
rect 100 27148 2580 27164
rect 100 27084 967 27148
rect 1031 27084 1059 27148
rect 1123 27084 1151 27148
rect 1215 27084 1243 27148
rect 1307 27084 1335 27148
rect 1399 27084 1427 27148
rect 1491 27084 2580 27148
rect 100 27068 2580 27084
rect 100 27004 967 27068
rect 1031 27004 1059 27068
rect 1123 27004 1151 27068
rect 1215 27004 1243 27068
rect 1307 27004 1335 27068
rect 1399 27004 1427 27068
rect 1491 27004 2580 27068
rect 100 26988 2580 27004
rect 100 26924 967 26988
rect 1031 26924 1059 26988
rect 1123 26924 1151 26988
rect 1215 26924 1243 26988
rect 1307 26924 1335 26988
rect 1399 26924 1427 26988
rect 1491 26924 2580 26988
rect 100 26908 2580 26924
rect 100 26844 967 26908
rect 1031 26844 1059 26908
rect 1123 26844 1151 26908
rect 1215 26844 1243 26908
rect 1307 26844 1335 26908
rect 1399 26844 1427 26908
rect 1491 26844 2580 26908
rect 100 26828 2580 26844
rect 100 26764 967 26828
rect 1031 26764 1059 26828
rect 1123 26764 1151 26828
rect 1215 26764 1243 26828
rect 1307 26764 1335 26828
rect 1399 26764 1427 26828
rect 1491 26764 2580 26828
rect 100 26748 2580 26764
rect 100 26684 967 26748
rect 1031 26684 1059 26748
rect 1123 26684 1151 26748
rect 1215 26684 1243 26748
rect 1307 26684 1335 26748
rect 1399 26684 1427 26748
rect 1491 26684 2580 26748
rect 100 26668 2580 26684
rect 100 26604 967 26668
rect 1031 26604 1059 26668
rect 1123 26604 1151 26668
rect 1215 26604 1243 26668
rect 1307 26604 1335 26668
rect 1399 26604 1427 26668
rect 1491 26604 2580 26668
rect 100 26588 2580 26604
rect 100 26524 967 26588
rect 1031 26524 1059 26588
rect 1123 26524 1151 26588
rect 1215 26524 1243 26588
rect 1307 26524 1335 26588
rect 1399 26524 1427 26588
rect 1491 26524 2580 26588
rect 100 26508 2580 26524
rect 100 26444 967 26508
rect 1031 26444 1059 26508
rect 1123 26444 1151 26508
rect 1215 26444 1243 26508
rect 1307 26444 1335 26508
rect 1399 26444 1427 26508
rect 1491 26444 2580 26508
rect 100 26428 2580 26444
rect 100 26364 967 26428
rect 1031 26364 1059 26428
rect 1123 26364 1151 26428
rect 1215 26364 1243 26428
rect 1307 26364 1335 26428
rect 1399 26364 1427 26428
rect 1491 26364 2580 26428
rect 100 26348 2580 26364
rect 100 26284 967 26348
rect 1031 26284 1059 26348
rect 1123 26284 1151 26348
rect 1215 26284 1243 26348
rect 1307 26284 1335 26348
rect 1399 26284 1427 26348
rect 1491 26284 2580 26348
rect 100 26268 2580 26284
rect 100 26204 967 26268
rect 1031 26204 1059 26268
rect 1123 26204 1151 26268
rect 1215 26204 1243 26268
rect 1307 26204 1335 26268
rect 1399 26204 1427 26268
rect 1491 26204 2580 26268
rect 100 26188 2580 26204
rect 100 26124 967 26188
rect 1031 26124 1059 26188
rect 1123 26124 1151 26188
rect 1215 26124 1243 26188
rect 1307 26124 1335 26188
rect 1399 26124 1427 26188
rect 1491 26124 2580 26188
rect 100 26108 2580 26124
rect 100 26044 967 26108
rect 1031 26044 1059 26108
rect 1123 26044 1151 26108
rect 1215 26044 1243 26108
rect 1307 26044 1335 26108
rect 1399 26044 1427 26108
rect 1491 26044 2580 26108
rect 100 26028 2580 26044
rect 100 25964 967 26028
rect 1031 25964 1059 26028
rect 1123 25964 1151 26028
rect 1215 25964 1243 26028
rect 1307 25964 1335 26028
rect 1399 25964 1427 26028
rect 1491 25964 2580 26028
rect 100 25948 2580 25964
rect 100 25884 967 25948
rect 1031 25884 1059 25948
rect 1123 25884 1151 25948
rect 1215 25884 1243 25948
rect 1307 25884 1335 25948
rect 1399 25884 1427 25948
rect 1491 25884 2580 25948
rect 100 25868 2580 25884
rect 100 25804 967 25868
rect 1031 25804 1059 25868
rect 1123 25804 1151 25868
rect 1215 25804 1243 25868
rect 1307 25804 1335 25868
rect 1399 25804 1427 25868
rect 1491 25804 2580 25868
rect 100 25788 2580 25804
rect 100 25724 967 25788
rect 1031 25724 1059 25788
rect 1123 25724 1151 25788
rect 1215 25724 1243 25788
rect 1307 25724 1335 25788
rect 1399 25724 1427 25788
rect 1491 25724 2580 25788
rect 100 25708 2580 25724
rect 100 25644 967 25708
rect 1031 25644 1059 25708
rect 1123 25644 1151 25708
rect 1215 25644 1243 25708
rect 1307 25644 1335 25708
rect 1399 25644 1427 25708
rect 1491 25644 2580 25708
rect 100 25628 2580 25644
rect 100 25564 967 25628
rect 1031 25564 1059 25628
rect 1123 25564 1151 25628
rect 1215 25564 1243 25628
rect 1307 25564 1335 25628
rect 1399 25564 1427 25628
rect 1491 25564 2580 25628
rect 100 25547 2580 25564
rect 100 25483 967 25547
rect 1031 25483 1059 25547
rect 1123 25483 1151 25547
rect 1215 25483 1243 25547
rect 1307 25483 1335 25547
rect 1399 25483 1427 25547
rect 1491 25483 2580 25547
rect 100 25466 2580 25483
rect 100 25402 967 25466
rect 1031 25402 1059 25466
rect 1123 25402 1151 25466
rect 1215 25402 1243 25466
rect 1307 25402 1335 25466
rect 1399 25402 1427 25466
rect 1491 25402 2580 25466
rect 100 25385 2580 25402
rect 100 25321 967 25385
rect 1031 25321 1059 25385
rect 1123 25321 1151 25385
rect 1215 25321 1243 25385
rect 1307 25321 1335 25385
rect 1399 25321 1427 25385
rect 1491 25321 2580 25385
rect 100 25304 2580 25321
rect 100 25240 967 25304
rect 1031 25240 1059 25304
rect 1123 25240 1151 25304
rect 1215 25240 1243 25304
rect 1307 25240 1335 25304
rect 1399 25240 1427 25304
rect 1491 25240 2580 25304
rect 100 25223 2580 25240
rect 100 25159 967 25223
rect 1031 25159 1059 25223
rect 1123 25159 1151 25223
rect 1215 25159 1243 25223
rect 1307 25159 1335 25223
rect 1399 25159 1427 25223
rect 1491 25159 2580 25223
rect 100 25142 2580 25159
rect 100 25078 967 25142
rect 1031 25078 1059 25142
rect 1123 25078 1151 25142
rect 1215 25078 1243 25142
rect 1307 25078 1335 25142
rect 1399 25078 1427 25142
rect 1491 25078 2580 25142
rect 100 25061 2580 25078
rect 100 24997 967 25061
rect 1031 24997 1059 25061
rect 1123 24997 1151 25061
rect 1215 24997 1243 25061
rect 1307 24997 1335 25061
rect 1399 24997 1427 25061
rect 1491 24997 2580 25061
rect 100 24980 2580 24997
rect 100 24916 967 24980
rect 1031 24916 1059 24980
rect 1123 24916 1151 24980
rect 1215 24916 1243 24980
rect 1307 24916 1335 24980
rect 1399 24916 1427 24980
rect 1491 24916 2580 24980
rect 100 24899 2580 24916
rect 100 24835 967 24899
rect 1031 24835 1059 24899
rect 1123 24835 1151 24899
rect 1215 24835 1243 24899
rect 1307 24835 1335 24899
rect 1399 24835 1427 24899
rect 1491 24835 2580 24899
rect 100 24818 2580 24835
rect 100 24754 967 24818
rect 1031 24754 1059 24818
rect 1123 24754 1151 24818
rect 1215 24754 1243 24818
rect 1307 24754 1335 24818
rect 1399 24754 1427 24818
rect 1491 24754 2580 24818
rect 100 24737 2580 24754
rect 100 24673 967 24737
rect 1031 24673 1059 24737
rect 1123 24673 1151 24737
rect 1215 24673 1243 24737
rect 1307 24673 1335 24737
rect 1399 24673 1427 24737
rect 1491 24673 2580 24737
rect 100 24656 2580 24673
rect 100 24592 967 24656
rect 1031 24592 1059 24656
rect 1123 24592 1151 24656
rect 1215 24592 1243 24656
rect 1307 24592 1335 24656
rect 1399 24592 1427 24656
rect 1491 24592 2580 24656
rect 100 24575 2580 24592
rect 100 24511 967 24575
rect 1031 24511 1059 24575
rect 1123 24511 1151 24575
rect 1215 24511 1243 24575
rect 1307 24511 1335 24575
rect 1399 24511 1427 24575
rect 1491 24511 2580 24575
rect 100 24494 2580 24511
rect 100 24430 967 24494
rect 1031 24430 1059 24494
rect 1123 24430 1151 24494
rect 1215 24430 1243 24494
rect 1307 24430 1335 24494
rect 1399 24430 1427 24494
rect 1491 24430 2580 24494
rect 100 24413 2580 24430
rect 100 24349 967 24413
rect 1031 24349 1059 24413
rect 1123 24349 1151 24413
rect 1215 24349 1243 24413
rect 1307 24349 1335 24413
rect 1399 24349 1427 24413
rect 1491 24349 2580 24413
rect 100 24332 2580 24349
rect 100 24268 967 24332
rect 1031 24268 1059 24332
rect 1123 24268 1151 24332
rect 1215 24268 1243 24332
rect 1307 24268 1335 24332
rect 1399 24268 1427 24332
rect 1491 24268 2580 24332
rect 100 24251 2580 24268
rect 100 24187 967 24251
rect 1031 24187 1059 24251
rect 1123 24187 1151 24251
rect 1215 24187 1243 24251
rect 1307 24187 1335 24251
rect 1399 24187 1427 24251
rect 1491 24187 2580 24251
rect 100 24170 2580 24187
rect 100 24106 967 24170
rect 1031 24106 1059 24170
rect 1123 24106 1151 24170
rect 1215 24106 1243 24170
rect 1307 24106 1335 24170
rect 1399 24106 1427 24170
rect 1491 24106 2580 24170
rect 100 24089 2580 24106
rect 100 24025 967 24089
rect 1031 24025 1059 24089
rect 1123 24025 1151 24089
rect 1215 24025 1243 24089
rect 1307 24025 1335 24089
rect 1399 24025 1427 24089
rect 1491 24025 2580 24089
rect 100 24008 2580 24025
rect 100 23944 967 24008
rect 1031 23944 1059 24008
rect 1123 23944 1151 24008
rect 1215 23944 1243 24008
rect 1307 23944 1335 24008
rect 1399 23944 1427 24008
rect 1491 23944 2580 24008
rect 100 23927 2580 23944
rect 100 23863 967 23927
rect 1031 23863 1059 23927
rect 1123 23863 1151 23927
rect 1215 23863 1243 23927
rect 1307 23863 1335 23927
rect 1399 23863 1427 23927
rect 1491 23863 2580 23927
rect 100 23846 2580 23863
rect 100 23782 967 23846
rect 1031 23782 1059 23846
rect 1123 23782 1151 23846
rect 1215 23782 1243 23846
rect 1307 23782 1335 23846
rect 1399 23782 1427 23846
rect 1491 23782 2580 23846
rect 100 23765 2580 23782
rect 100 23701 967 23765
rect 1031 23701 1059 23765
rect 1123 23701 1151 23765
rect 1215 23701 1243 23765
rect 1307 23701 1335 23765
rect 1399 23701 1427 23765
rect 1491 23701 2580 23765
rect 100 23684 2580 23701
rect 100 23620 967 23684
rect 1031 23620 1059 23684
rect 1123 23620 1151 23684
rect 1215 23620 1243 23684
rect 1307 23620 1335 23684
rect 1399 23620 1427 23684
rect 1491 23620 2580 23684
rect 100 23603 2580 23620
rect 100 23539 967 23603
rect 1031 23539 1059 23603
rect 1123 23539 1151 23603
rect 1215 23539 1243 23603
rect 1307 23539 1335 23603
rect 1399 23539 1427 23603
rect 1491 23539 2580 23603
rect 100 23522 2580 23539
rect 100 23458 967 23522
rect 1031 23458 1059 23522
rect 1123 23458 1151 23522
rect 1215 23458 1243 23522
rect 1307 23458 1335 23522
rect 1399 23458 1427 23522
rect 1491 23458 2580 23522
rect 100 23441 2580 23458
rect 100 23377 967 23441
rect 1031 23377 1059 23441
rect 1123 23377 1151 23441
rect 1215 23377 1243 23441
rect 1307 23377 1335 23441
rect 1399 23377 1427 23441
rect 1491 23377 2580 23441
rect 100 23360 2580 23377
rect 100 23296 967 23360
rect 1031 23296 1059 23360
rect 1123 23296 1151 23360
rect 1215 23296 1243 23360
rect 1307 23296 1335 23360
rect 1399 23296 1427 23360
rect 1491 23296 2580 23360
rect 100 23279 2580 23296
rect 100 23215 967 23279
rect 1031 23215 1059 23279
rect 1123 23215 1151 23279
rect 1215 23215 1243 23279
rect 1307 23215 1335 23279
rect 1399 23215 1427 23279
rect 1491 23215 2580 23279
rect 100 23198 2580 23215
rect 100 23134 967 23198
rect 1031 23134 1059 23198
rect 1123 23134 1151 23198
rect 1215 23134 1243 23198
rect 1307 23134 1335 23198
rect 1399 23134 1427 23198
rect 1491 23134 2580 23198
rect 100 23117 2580 23134
rect 100 23053 967 23117
rect 1031 23053 1059 23117
rect 1123 23053 1151 23117
rect 1215 23053 1243 23117
rect 1307 23053 1335 23117
rect 1399 23053 1427 23117
rect 1491 23053 2580 23117
rect 100 23036 2580 23053
rect 100 22972 967 23036
rect 1031 22972 1059 23036
rect 1123 22972 1151 23036
rect 1215 22972 1243 23036
rect 1307 22972 1335 23036
rect 1399 22972 1427 23036
rect 1491 22972 2580 23036
rect 100 22955 2580 22972
rect 100 22891 967 22955
rect 1031 22891 1059 22955
rect 1123 22891 1151 22955
rect 1215 22891 1243 22955
rect 1307 22891 1335 22955
rect 1399 22891 1427 22955
rect 1491 22891 2580 22955
rect 100 22874 2580 22891
rect 100 22810 967 22874
rect 1031 22810 1059 22874
rect 1123 22810 1151 22874
rect 1215 22810 1243 22874
rect 1307 22810 1335 22874
rect 1399 22810 1427 22874
rect 1491 22810 2580 22874
rect 100 22793 2580 22810
rect 100 22729 967 22793
rect 1031 22729 1059 22793
rect 1123 22729 1151 22793
rect 1215 22729 1243 22793
rect 1307 22729 1335 22793
rect 1399 22729 1427 22793
rect 1491 22729 2580 22793
rect 100 22712 2580 22729
rect 100 22648 967 22712
rect 1031 22648 1059 22712
rect 1123 22648 1151 22712
rect 1215 22648 1243 22712
rect 1307 22648 1335 22712
rect 1399 22648 1427 22712
rect 1491 22648 2580 22712
rect 100 22631 2580 22648
rect 100 22567 967 22631
rect 1031 22567 1059 22631
rect 1123 22567 1151 22631
rect 1215 22567 1243 22631
rect 1307 22567 1335 22631
rect 1399 22567 1427 22631
rect 1491 22567 2580 22631
rect 100 22550 2580 22567
rect 100 22486 967 22550
rect 1031 22486 1059 22550
rect 1123 22486 1151 22550
rect 1215 22486 1243 22550
rect 1307 22486 1335 22550
rect 1399 22486 1427 22550
rect 1491 22486 2580 22550
rect 100 22469 2580 22486
rect 100 22405 967 22469
rect 1031 22405 1059 22469
rect 1123 22405 1151 22469
rect 1215 22405 1243 22469
rect 1307 22405 1335 22469
rect 1399 22405 1427 22469
rect 1491 22405 2580 22469
rect 100 22388 2580 22405
rect 100 22324 967 22388
rect 1031 22324 1059 22388
rect 1123 22324 1151 22388
rect 1215 22324 1243 22388
rect 1307 22324 1335 22388
rect 1399 22324 1427 22388
rect 1491 22324 2580 22388
rect 100 22307 2580 22324
rect 100 22243 967 22307
rect 1031 22243 1059 22307
rect 1123 22243 1151 22307
rect 1215 22243 1243 22307
rect 1307 22243 1335 22307
rect 1399 22243 1427 22307
rect 1491 22243 2580 22307
rect 100 22226 2580 22243
rect 100 22162 967 22226
rect 1031 22162 1059 22226
rect 1123 22162 1151 22226
rect 1215 22162 1243 22226
rect 1307 22162 1335 22226
rect 1399 22162 1427 22226
rect 1491 22162 2580 22226
rect 100 22145 2580 22162
rect 100 22081 967 22145
rect 1031 22081 1059 22145
rect 1123 22081 1151 22145
rect 1215 22081 1243 22145
rect 1307 22081 1335 22145
rect 1399 22081 1427 22145
rect 1491 22081 2580 22145
rect 100 22064 2580 22081
rect 100 22000 967 22064
rect 1031 22000 1059 22064
rect 1123 22000 1151 22064
rect 1215 22000 1243 22064
rect 1307 22000 1335 22064
rect 1399 22000 1427 22064
rect 1491 22000 2580 22064
rect 100 21983 2580 22000
rect 100 21919 967 21983
rect 1031 21919 1059 21983
rect 1123 21919 1151 21983
rect 1215 21919 1243 21983
rect 1307 21919 1335 21983
rect 1399 21919 1427 21983
rect 1491 21919 2580 21983
rect 100 21902 2580 21919
rect 100 21838 967 21902
rect 1031 21838 1059 21902
rect 1123 21838 1151 21902
rect 1215 21838 1243 21902
rect 1307 21838 1335 21902
rect 1399 21838 1427 21902
rect 1491 21838 2580 21902
rect 100 21821 2580 21838
rect 100 21757 967 21821
rect 1031 21757 1059 21821
rect 1123 21757 1151 21821
rect 1215 21757 1243 21821
rect 1307 21757 1335 21821
rect 1399 21757 1427 21821
rect 1491 21757 2580 21821
rect 100 21740 2580 21757
rect 100 21676 967 21740
rect 1031 21676 1059 21740
rect 1123 21676 1151 21740
rect 1215 21676 1243 21740
rect 1307 21676 1335 21740
rect 1399 21676 1427 21740
rect 1491 21676 2580 21740
rect 100 21659 2580 21676
rect 100 21595 967 21659
rect 1031 21595 1059 21659
rect 1123 21595 1151 21659
rect 1215 21595 1243 21659
rect 1307 21595 1335 21659
rect 1399 21595 1427 21659
rect 1491 21595 2580 21659
rect 100 21578 2580 21595
rect 100 21514 967 21578
rect 1031 21514 1059 21578
rect 1123 21514 1151 21578
rect 1215 21514 1243 21578
rect 1307 21514 1335 21578
rect 1399 21514 1427 21578
rect 1491 21514 2580 21578
rect 100 21497 2580 21514
rect 100 21433 967 21497
rect 1031 21433 1059 21497
rect 1123 21433 1151 21497
rect 1215 21433 1243 21497
rect 1307 21433 1335 21497
rect 1399 21433 1427 21497
rect 1491 21433 2580 21497
rect 100 21416 2580 21433
rect 100 21352 967 21416
rect 1031 21352 1059 21416
rect 1123 21352 1151 21416
rect 1215 21352 1243 21416
rect 1307 21352 1335 21416
rect 1399 21352 1427 21416
rect 1491 21352 2580 21416
rect 100 21335 2580 21352
rect 100 21271 967 21335
rect 1031 21271 1059 21335
rect 1123 21271 1151 21335
rect 1215 21271 1243 21335
rect 1307 21271 1335 21335
rect 1399 21271 1427 21335
rect 1491 21271 2580 21335
rect 100 21254 2580 21271
rect 100 21190 967 21254
rect 1031 21190 1059 21254
rect 1123 21190 1151 21254
rect 1215 21190 1243 21254
rect 1307 21190 1335 21254
rect 1399 21190 1427 21254
rect 1491 21190 2580 21254
rect 100 21173 2580 21190
rect 100 21109 967 21173
rect 1031 21109 1059 21173
rect 1123 21109 1151 21173
rect 1215 21109 1243 21173
rect 1307 21109 1335 21173
rect 1399 21109 1427 21173
rect 1491 21109 2580 21173
rect 100 21092 2580 21109
rect 100 21028 967 21092
rect 1031 21028 1059 21092
rect 1123 21028 1151 21092
rect 1215 21028 1243 21092
rect 1307 21028 1335 21092
rect 1399 21028 1427 21092
rect 1491 21028 2580 21092
rect 100 21011 2580 21028
rect 100 20947 967 21011
rect 1031 20947 1059 21011
rect 1123 20947 1151 21011
rect 1215 20947 1243 21011
rect 1307 20947 1335 21011
rect 1399 20947 1427 21011
rect 1491 20947 2580 21011
rect 100 20930 2580 20947
rect 100 20866 967 20930
rect 1031 20866 1059 20930
rect 1123 20866 1151 20930
rect 1215 20866 1243 20930
rect 1307 20866 1335 20930
rect 1399 20866 1427 20930
rect 1491 20866 2580 20930
rect 100 20849 2580 20866
rect 100 20785 967 20849
rect 1031 20785 1059 20849
rect 1123 20785 1151 20849
rect 1215 20785 1243 20849
rect 1307 20785 1335 20849
rect 1399 20785 1427 20849
rect 1491 20785 2580 20849
rect 100 20768 2580 20785
rect 100 20704 967 20768
rect 1031 20704 1059 20768
rect 1123 20704 1151 20768
rect 1215 20704 1243 20768
rect 1307 20704 1335 20768
rect 1399 20704 1427 20768
rect 1491 20704 2580 20768
rect 100 20687 2580 20704
rect 100 20623 967 20687
rect 1031 20623 1059 20687
rect 1123 20623 1151 20687
rect 1215 20623 1243 20687
rect 1307 20623 1335 20687
rect 1399 20623 1427 20687
rect 1491 20623 2580 20687
rect 100 20606 2580 20623
rect 100 20542 967 20606
rect 1031 20542 1059 20606
rect 1123 20542 1151 20606
rect 1215 20542 1243 20606
rect 1307 20542 1335 20606
rect 1399 20542 1427 20606
rect 1491 20542 2580 20606
rect 100 20534 2580 20542
rect 100 20525 1543 20534
rect 100 20461 967 20525
rect 1031 20461 1059 20525
rect 1123 20461 1151 20525
rect 1215 20461 1243 20525
rect 1307 20461 1335 20525
rect 1399 20461 1427 20525
rect 1491 20470 1543 20525
rect 1607 20470 2580 20534
rect 1491 20461 2580 20470
rect 100 20431 2580 20461
rect 100 20415 1215 20431
rect 100 20351 1089 20415
rect 1153 20367 1215 20415
rect 1279 20367 1297 20431
rect 1361 20367 1379 20431
rect 1443 20367 1461 20431
rect 1525 20367 1543 20431
rect 1607 20367 1624 20431
rect 1688 20367 2580 20431
rect 1153 20351 2580 20367
rect 100 20311 2580 20351
rect 100 20283 1766 20311
rect 100 20219 1215 20283
rect 1279 20219 1297 20283
rect 1361 20219 1379 20283
rect 1443 20219 1461 20283
rect 1525 20219 1543 20283
rect 1607 20219 1624 20283
rect 1688 20247 1766 20283
rect 1830 20247 2580 20311
rect 1688 20219 2580 20247
rect 100 20203 2580 20219
rect 100 20192 1471 20203
rect 100 20128 1312 20192
rect 1376 20139 1471 20192
rect 1535 20139 1553 20203
rect 1617 20139 1635 20203
rect 1699 20139 1717 20203
rect 1781 20139 1799 20203
rect 1863 20139 1880 20203
rect 1944 20139 2580 20203
rect 1376 20128 2580 20139
rect 100 20072 2580 20128
rect 100 20055 2005 20072
rect 100 19991 1471 20055
rect 1535 19991 1553 20055
rect 1617 19991 1635 20055
rect 1699 19991 1717 20055
rect 1781 19991 1799 20055
rect 1863 19991 1880 20055
rect 1944 20008 2005 20055
rect 2069 20008 2580 20072
rect 1944 19991 2580 20008
rect 100 19975 2580 19991
rect 100 19953 1669 19975
rect 100 19889 1551 19953
rect 1615 19911 1669 19953
rect 1733 19911 1751 19975
rect 1815 19911 1833 19975
rect 1897 19911 1915 19975
rect 1979 19911 1997 19975
rect 2061 19911 2078 19975
rect 2142 19911 2580 19975
rect 1615 19889 2580 19911
rect 100 19857 2580 19889
rect 100 19827 2220 19857
rect 100 19763 1669 19827
rect 1733 19763 1751 19827
rect 1815 19763 1833 19827
rect 1897 19763 1915 19827
rect 1979 19763 1997 19827
rect 2061 19763 2078 19827
rect 2142 19793 2220 19827
rect 2284 19793 2580 19857
rect 2142 19763 2580 19793
rect 100 19742 2580 19763
rect 100 19738 1893 19742
rect 100 19674 1766 19738
rect 1830 19678 1893 19738
rect 1957 19678 1975 19742
rect 2039 19678 2057 19742
rect 2121 19678 2139 19742
rect 2203 19678 2221 19742
rect 2285 19678 2302 19742
rect 2366 19678 2580 19742
rect 1830 19674 2580 19678
rect 100 19658 2580 19674
rect 100 19594 2394 19658
rect 2458 19594 2502 19658
rect 2566 19594 2580 19658
rect 100 19530 1893 19594
rect 1957 19530 1975 19594
rect 2039 19530 2057 19594
rect 2121 19530 2139 19594
rect 2203 19530 2221 19594
rect 2285 19530 2302 19594
rect 2366 19549 2580 19594
rect 2366 19530 2394 19549
rect 100 19508 2394 19530
rect 100 19499 2120 19508
rect 100 19435 1998 19499
rect 2062 19444 2120 19499
rect 2184 19444 2211 19508
rect 2275 19444 2302 19508
rect 2366 19485 2394 19508
rect 2458 19485 2502 19549
rect 2566 19485 2580 19549
rect 2366 19444 2580 19485
rect 2062 19440 2580 19444
rect 2062 19435 2394 19440
rect 100 19376 2394 19435
rect 2458 19376 2502 19440
rect 2566 19376 2580 19440
rect 100 19360 2580 19376
rect 100 19296 2120 19360
rect 2184 19296 2211 19360
rect 2275 19296 2302 19360
rect 2366 19332 2580 19360
rect 2366 19296 2394 19332
rect 100 19275 2394 19296
rect 100 19211 2220 19275
rect 2284 19211 2305 19275
rect 2369 19268 2394 19275
rect 2458 19268 2502 19332
rect 2566 19268 2580 19332
rect 2369 19224 2580 19268
rect 2369 19211 2394 19224
rect 100 19160 2394 19211
rect 2458 19160 2502 19224
rect 2566 19160 2580 19224
rect 100 18472 2580 19160
rect 3121 34122 5023 35370
rect 3121 33896 4786 34122
rect 3121 33840 3513 33896
rect 3569 33840 3594 33896
rect 3650 33840 3675 33896
rect 3731 33840 3757 33896
rect 3813 33840 3839 33896
rect 3895 33840 3921 33896
rect 3977 33840 4003 33896
rect 4059 33840 4085 33896
rect 4141 33840 4167 33896
rect 4223 33840 4249 33896
rect 4305 33886 4786 33896
rect 4305 33880 4556 33886
rect 4305 33840 4354 33880
rect 3121 33824 4354 33840
rect 4410 33824 4446 33880
rect 4502 33830 4556 33880
rect 4612 33885 4786 33886
tri 4786 33885 5023 34122 nw
rect 5207 37892 7385 37903
rect 5207 37836 5216 37892
rect 5272 37836 5297 37892
rect 5353 37836 5378 37892
rect 5434 37836 5459 37892
rect 5515 37836 5540 37892
rect 5596 37836 5621 37892
rect 5677 37836 5702 37892
rect 5758 37836 5783 37892
rect 5839 37836 5864 37892
rect 5920 37836 5945 37892
rect 6001 37836 6026 37892
rect 6082 37836 6107 37892
rect 6163 37836 6188 37892
rect 6244 37836 6269 37892
rect 6325 37836 6350 37892
rect 6406 37836 6431 37892
rect 6487 37836 6512 37892
rect 6568 37836 6593 37892
rect 6649 37836 6674 37892
rect 6730 37836 6755 37892
rect 6811 37836 6836 37892
rect 6892 37836 6917 37892
rect 6973 37836 6998 37892
rect 7054 37836 7079 37892
rect 7135 37836 7160 37892
rect 5207 37812 7160 37836
rect 5207 37756 5216 37812
rect 5272 37756 5297 37812
rect 5353 37756 5378 37812
rect 5434 37756 5459 37812
rect 5515 37756 5540 37812
rect 5596 37756 5621 37812
rect 5677 37756 5702 37812
rect 5758 37756 5783 37812
rect 5839 37756 5864 37812
rect 5920 37756 5945 37812
rect 6001 37756 6026 37812
rect 6082 37756 6107 37812
rect 6163 37756 6188 37812
rect 6244 37756 6269 37812
rect 6325 37756 6350 37812
rect 6406 37756 6431 37812
rect 6487 37756 6512 37812
rect 6568 37756 6593 37812
rect 6649 37756 6674 37812
rect 6730 37756 6755 37812
rect 6811 37756 6836 37812
rect 6892 37756 6917 37812
rect 6973 37756 6998 37812
rect 7054 37756 7079 37812
rect 7135 37756 7160 37812
rect 5207 37732 7160 37756
rect 5207 37676 5216 37732
rect 5272 37676 5297 37732
rect 5353 37676 5378 37732
rect 5434 37676 5459 37732
rect 5515 37676 5540 37732
rect 5596 37676 5621 37732
rect 5677 37676 5702 37732
rect 5758 37676 5783 37732
rect 5839 37676 5864 37732
rect 5920 37676 5945 37732
rect 6001 37676 6026 37732
rect 6082 37676 6107 37732
rect 6163 37676 6188 37732
rect 6244 37676 6269 37732
rect 6325 37676 6350 37732
rect 6406 37676 6431 37732
rect 6487 37676 6512 37732
rect 6568 37676 6593 37732
rect 6649 37676 6674 37732
rect 6730 37676 6755 37732
rect 6811 37676 6836 37732
rect 6892 37676 6917 37732
rect 6973 37676 6998 37732
rect 7054 37676 7079 37732
rect 7135 37676 7160 37732
rect 5207 37652 7160 37676
rect 5207 37596 5216 37652
rect 5272 37596 5297 37652
rect 5353 37596 5378 37652
rect 5434 37596 5459 37652
rect 5515 37596 5540 37652
rect 5596 37596 5621 37652
rect 5677 37596 5702 37652
rect 5758 37596 5783 37652
rect 5839 37596 5864 37652
rect 5920 37596 5945 37652
rect 6001 37596 6026 37652
rect 6082 37596 6107 37652
rect 6163 37596 6188 37652
rect 6244 37596 6269 37652
rect 6325 37596 6350 37652
rect 6406 37596 6431 37652
rect 6487 37596 6512 37652
rect 6568 37596 6593 37652
rect 6649 37596 6674 37652
rect 6730 37596 6755 37652
rect 6811 37596 6836 37652
rect 6892 37596 6917 37652
rect 6973 37596 6998 37652
rect 7054 37596 7079 37652
rect 7135 37596 7160 37652
rect 5207 37572 7160 37596
rect 5207 37516 5216 37572
rect 5272 37516 5297 37572
rect 5353 37516 5378 37572
rect 5434 37516 5459 37572
rect 5515 37516 5540 37572
rect 5596 37516 5621 37572
rect 5677 37516 5702 37572
rect 5758 37516 5783 37572
rect 5839 37516 5864 37572
rect 5920 37516 5945 37572
rect 6001 37516 6026 37572
rect 6082 37516 6107 37572
rect 6163 37516 6188 37572
rect 6244 37516 6269 37572
rect 6325 37516 6350 37572
rect 6406 37516 6431 37572
rect 6487 37516 6512 37572
rect 6568 37516 6593 37572
rect 6649 37516 6674 37572
rect 6730 37516 6755 37572
rect 6811 37516 6836 37572
rect 6892 37516 6917 37572
rect 6973 37516 6998 37572
rect 7054 37516 7079 37572
rect 7135 37516 7160 37572
rect 5207 37492 7160 37516
rect 5207 37436 5216 37492
rect 5272 37436 5297 37492
rect 5353 37436 5378 37492
rect 5434 37436 5459 37492
rect 5515 37436 5540 37492
rect 5596 37436 5621 37492
rect 5677 37436 5702 37492
rect 5758 37436 5783 37492
rect 5839 37436 5864 37492
rect 5920 37436 5945 37492
rect 6001 37436 6026 37492
rect 6082 37436 6107 37492
rect 6163 37436 6188 37492
rect 6244 37436 6269 37492
rect 6325 37436 6350 37492
rect 6406 37436 6431 37492
rect 6487 37436 6512 37492
rect 6568 37436 6593 37492
rect 6649 37436 6674 37492
rect 6730 37436 6755 37492
rect 6811 37436 6836 37492
rect 6892 37436 6917 37492
rect 6973 37436 6998 37492
rect 7054 37436 7079 37492
rect 7135 37436 7160 37492
rect 5207 37412 7160 37436
rect 5207 37356 5216 37412
rect 5272 37356 5297 37412
rect 5353 37356 5378 37412
rect 5434 37356 5459 37412
rect 5515 37356 5540 37412
rect 5596 37356 5621 37412
rect 5677 37356 5702 37412
rect 5758 37356 5783 37412
rect 5839 37356 5864 37412
rect 5920 37356 5945 37412
rect 6001 37356 6026 37412
rect 6082 37356 6107 37412
rect 6163 37356 6188 37412
rect 6244 37356 6269 37412
rect 6325 37356 6350 37412
rect 6406 37356 6431 37412
rect 6487 37356 6512 37412
rect 6568 37356 6593 37412
rect 6649 37356 6674 37412
rect 6730 37356 6755 37412
rect 6811 37356 6836 37412
rect 6892 37356 6917 37412
rect 6973 37356 6998 37412
rect 7054 37356 7079 37412
rect 7135 37356 7160 37412
rect 5207 37332 7160 37356
rect 5207 37276 5216 37332
rect 5272 37276 5297 37332
rect 5353 37276 5378 37332
rect 5434 37276 5459 37332
rect 5515 37276 5540 37332
rect 5596 37276 5621 37332
rect 5677 37276 5702 37332
rect 5758 37276 5783 37332
rect 5839 37276 5864 37332
rect 5920 37276 5945 37332
rect 6001 37276 6026 37332
rect 6082 37276 6107 37332
rect 6163 37276 6188 37332
rect 6244 37276 6269 37332
rect 6325 37276 6350 37332
rect 6406 37276 6431 37332
rect 6487 37276 6512 37332
rect 6568 37276 6593 37332
rect 6649 37276 6674 37332
rect 6730 37276 6755 37332
rect 6811 37276 6836 37332
rect 6892 37276 6917 37332
rect 6973 37276 6998 37332
rect 7054 37276 7079 37332
rect 7135 37276 7160 37332
rect 5207 37252 7160 37276
rect 5207 37196 5216 37252
rect 5272 37196 5297 37252
rect 5353 37196 5378 37252
rect 5434 37196 5459 37252
rect 5515 37196 5540 37252
rect 5596 37196 5621 37252
rect 5677 37196 5702 37252
rect 5758 37196 5783 37252
rect 5839 37196 5864 37252
rect 5920 37196 5945 37252
rect 6001 37196 6026 37252
rect 6082 37196 6107 37252
rect 6163 37196 6188 37252
rect 6244 37196 6269 37252
rect 6325 37196 6350 37252
rect 6406 37196 6431 37252
rect 6487 37196 6512 37252
rect 6568 37196 6593 37252
rect 6649 37196 6674 37252
rect 6730 37196 6755 37252
rect 6811 37196 6836 37252
rect 6892 37196 6917 37252
rect 6973 37196 6998 37252
rect 7054 37196 7079 37252
rect 7135 37196 7160 37252
rect 5207 37172 7160 37196
rect 5207 37116 5216 37172
rect 5272 37116 5297 37172
rect 5353 37116 5378 37172
rect 5434 37116 5459 37172
rect 5515 37116 5540 37172
rect 5596 37116 5621 37172
rect 5677 37116 5702 37172
rect 5758 37116 5783 37172
rect 5839 37116 5864 37172
rect 5920 37116 5945 37172
rect 6001 37116 6026 37172
rect 6082 37116 6107 37172
rect 6163 37116 6188 37172
rect 6244 37116 6269 37172
rect 6325 37116 6350 37172
rect 6406 37116 6431 37172
rect 6487 37116 6512 37172
rect 6568 37116 6593 37172
rect 6649 37116 6674 37172
rect 6730 37116 6755 37172
rect 6811 37116 6836 37172
rect 6892 37116 6917 37172
rect 6973 37116 6998 37172
rect 7054 37116 7079 37172
rect 7135 37116 7160 37172
rect 5207 37092 7160 37116
rect 5207 37036 5216 37092
rect 5272 37036 5297 37092
rect 5353 37036 5378 37092
rect 5434 37036 5459 37092
rect 5515 37036 5540 37092
rect 5596 37036 5621 37092
rect 5677 37036 5702 37092
rect 5758 37036 5783 37092
rect 5839 37036 5864 37092
rect 5920 37036 5945 37092
rect 6001 37036 6026 37092
rect 6082 37036 6107 37092
rect 6163 37036 6188 37092
rect 6244 37036 6269 37092
rect 6325 37036 6350 37092
rect 6406 37036 6431 37092
rect 6487 37036 6512 37092
rect 6568 37036 6593 37092
rect 6649 37036 6674 37092
rect 6730 37036 6755 37092
rect 6811 37036 6836 37092
rect 6892 37036 6917 37092
rect 6973 37036 6998 37092
rect 7054 37036 7079 37092
rect 7135 37036 7160 37092
rect 7376 37036 7385 37892
rect 5207 35877 7385 37036
rect 5207 35821 5215 35877
rect 5271 35821 5296 35877
rect 5352 35821 5377 35877
rect 5433 35821 5458 35877
rect 5514 35821 5539 35877
rect 5595 35821 5620 35877
rect 5676 35821 5701 35877
rect 5757 35821 5782 35877
rect 5838 35821 5863 35877
rect 5919 35821 5944 35877
rect 6000 35821 6025 35877
rect 6081 35821 6106 35877
rect 6162 35821 6187 35877
rect 6243 35821 6268 35877
rect 6324 35821 6349 35877
rect 6405 35821 6430 35877
rect 6486 35821 6511 35877
rect 6567 35821 6592 35877
rect 6648 35821 6673 35877
rect 6729 35821 6754 35877
rect 6810 35821 6835 35877
rect 6891 35821 6916 35877
rect 6972 35821 6997 35877
rect 7053 35821 7078 35877
rect 7134 35821 7159 35877
rect 7215 35821 7240 35877
rect 7296 35821 7320 35877
rect 7376 35821 7385 35877
rect 5207 35789 7385 35821
rect 5207 35733 5215 35789
rect 5271 35733 5296 35789
rect 5352 35733 5377 35789
rect 5433 35733 5458 35789
rect 5514 35733 5539 35789
rect 5595 35733 5620 35789
rect 5676 35733 5701 35789
rect 5757 35733 5782 35789
rect 5838 35733 5863 35789
rect 5919 35733 5944 35789
rect 6000 35733 6025 35789
rect 6081 35733 6106 35789
rect 6162 35733 6187 35789
rect 6243 35733 6268 35789
rect 6324 35733 6349 35789
rect 6405 35733 6430 35789
rect 6486 35733 6511 35789
rect 6567 35733 6592 35789
rect 6648 35733 6673 35789
rect 6729 35733 6754 35789
rect 6810 35733 6835 35789
rect 6891 35733 6916 35789
rect 6972 35733 6997 35789
rect 7053 35733 7078 35789
rect 7134 35733 7159 35789
rect 7215 35733 7240 35789
rect 7296 35733 7320 35789
rect 7376 35733 7385 35789
rect 5207 35701 7385 35733
rect 5207 35645 5215 35701
rect 5271 35645 5296 35701
rect 5352 35645 5377 35701
rect 5433 35645 5458 35701
rect 5514 35645 5539 35701
rect 5595 35645 5620 35701
rect 5676 35645 5701 35701
rect 5757 35645 5782 35701
rect 5838 35645 5863 35701
rect 5919 35645 5944 35701
rect 6000 35645 6025 35701
rect 6081 35645 6106 35701
rect 6162 35645 6187 35701
rect 6243 35645 6268 35701
rect 6324 35645 6349 35701
rect 6405 35645 6430 35701
rect 6486 35645 6511 35701
rect 6567 35645 6592 35701
rect 6648 35645 6673 35701
rect 6729 35645 6754 35701
rect 6810 35645 6835 35701
rect 6891 35645 6916 35701
rect 6972 35645 6997 35701
rect 7053 35645 7078 35701
rect 7134 35645 7159 35701
rect 7215 35645 7240 35701
rect 7296 35645 7320 35701
rect 7376 35645 7385 35701
rect 5207 35613 7385 35645
rect 5207 35557 5215 35613
rect 5271 35557 5296 35613
rect 5352 35557 5377 35613
rect 5433 35557 5458 35613
rect 5514 35557 5539 35613
rect 5595 35557 5620 35613
rect 5676 35557 5701 35613
rect 5757 35557 5782 35613
rect 5838 35557 5863 35613
rect 5919 35557 5944 35613
rect 6000 35557 6025 35613
rect 6081 35557 6106 35613
rect 6162 35557 6187 35613
rect 6243 35557 6268 35613
rect 6324 35557 6349 35613
rect 6405 35557 6430 35613
rect 6486 35557 6511 35613
rect 6567 35557 6592 35613
rect 6648 35557 6673 35613
rect 6729 35557 6754 35613
rect 6810 35557 6835 35613
rect 6891 35557 6916 35613
rect 6972 35557 6997 35613
rect 7053 35557 7078 35613
rect 7134 35557 7159 35613
rect 7215 35557 7240 35613
rect 7296 35557 7320 35613
rect 7376 35557 7385 35613
rect 5207 35525 7385 35557
rect 5207 35469 5215 35525
rect 5271 35469 5296 35525
rect 5352 35469 5377 35525
rect 5433 35469 5458 35525
rect 5514 35469 5539 35525
rect 5595 35469 5620 35525
rect 5676 35469 5701 35525
rect 5757 35469 5782 35525
rect 5838 35469 5863 35525
rect 5919 35469 5944 35525
rect 6000 35469 6025 35525
rect 6081 35469 6106 35525
rect 6162 35469 6187 35525
rect 6243 35469 6268 35525
rect 6324 35469 6349 35525
rect 6405 35469 6430 35525
rect 6486 35469 6511 35525
rect 6567 35469 6592 35525
rect 6648 35469 6673 35525
rect 6729 35469 6754 35525
rect 6810 35469 6835 35525
rect 6891 35469 6916 35525
rect 6972 35469 6997 35525
rect 7053 35469 7078 35525
rect 7134 35469 7159 35525
rect 7215 35469 7240 35525
rect 7296 35469 7320 35525
rect 7376 35469 7385 35525
rect 5207 35437 7385 35469
rect 5207 35381 5215 35437
rect 5271 35381 5296 35437
rect 5352 35381 5377 35437
rect 5433 35381 5458 35437
rect 5514 35381 5539 35437
rect 5595 35381 5620 35437
rect 5676 35381 5701 35437
rect 5757 35381 5782 35437
rect 5838 35381 5863 35437
rect 5919 35381 5944 35437
rect 6000 35381 6025 35437
rect 6081 35381 6106 35437
rect 6162 35381 6187 35437
rect 6243 35381 6268 35437
rect 6324 35381 6349 35437
rect 6405 35381 6430 35437
rect 6486 35381 6511 35437
rect 6567 35381 6592 35437
rect 6648 35381 6673 35437
rect 6729 35381 6754 35437
rect 6810 35381 6835 35437
rect 6891 35381 6916 35437
rect 6972 35381 6997 35437
rect 7053 35381 7078 35437
rect 7134 35381 7159 35437
rect 7215 35381 7240 35437
rect 7296 35381 7320 35437
rect 7376 35381 7385 35437
rect 4612 33881 4782 33885
tri 4782 33881 4786 33885 nw
rect 4612 33878 4779 33881
tri 4779 33878 4782 33881 nw
rect 5207 33878 7385 35381
rect 4612 33830 4723 33878
rect 4502 33824 4723 33830
rect 3121 33822 4723 33824
tri 4723 33822 4779 33878 nw
rect 5207 33822 5216 33878
rect 5272 33822 5299 33878
rect 5355 33822 5382 33878
rect 5438 33822 5465 33878
rect 5521 33822 5548 33878
rect 5604 33822 5631 33878
rect 5687 33822 5714 33878
rect 5770 33822 5797 33878
rect 5853 33822 5880 33878
rect 5936 33822 5963 33878
rect 6019 33822 6046 33878
rect 6102 33822 6129 33878
rect 6185 33822 6211 33878
rect 6267 33822 6293 33878
rect 6349 33822 6375 33878
rect 6431 33822 6457 33878
rect 6513 33822 6539 33878
rect 6595 33822 6621 33878
rect 6677 33822 6703 33878
rect 6759 33822 6785 33878
rect 6841 33822 6867 33878
rect 6923 33822 6949 33878
rect 7005 33822 7031 33878
rect 7087 33822 7113 33878
rect 7169 33822 7195 33878
rect 7251 33822 7385 33878
rect 3121 33804 4703 33822
rect 3121 33802 4556 33804
rect 3121 33746 3513 33802
rect 3569 33746 3594 33802
rect 3650 33746 3675 33802
rect 3731 33746 3757 33802
rect 3813 33746 3839 33802
rect 3895 33746 3921 33802
rect 3977 33746 4003 33802
rect 4059 33746 4085 33802
rect 4141 33746 4167 33802
rect 4223 33746 4249 33802
rect 4305 33780 4556 33802
rect 4305 33746 4354 33780
rect 3121 33724 4354 33746
rect 4410 33724 4446 33780
rect 4502 33748 4556 33780
rect 4612 33802 4703 33804
tri 4703 33802 4723 33822 nw
rect 4612 33790 4691 33802
tri 4691 33790 4703 33802 nw
rect 5207 33790 7385 33822
rect 7589 37892 9767 37903
rect 7589 37836 7598 37892
rect 7654 37836 7679 37892
rect 7735 37836 7760 37892
rect 7816 37836 7841 37892
rect 7897 37836 7922 37892
rect 7978 37836 8003 37892
rect 8059 37836 8084 37892
rect 8140 37836 8165 37892
rect 8221 37836 8246 37892
rect 8302 37836 8327 37892
rect 8383 37836 8408 37892
rect 8464 37836 8489 37892
rect 8545 37836 8570 37892
rect 8626 37836 8651 37892
rect 8707 37836 8732 37892
rect 8788 37836 8813 37892
rect 8869 37836 8894 37892
rect 8950 37836 8975 37892
rect 9031 37836 9056 37892
rect 9112 37836 9137 37892
rect 9193 37836 9218 37892
rect 9274 37836 9299 37892
rect 9355 37836 9380 37892
rect 9436 37836 9461 37892
rect 9517 37836 9542 37892
rect 7589 37812 9542 37836
rect 7589 37756 7598 37812
rect 7654 37756 7679 37812
rect 7735 37756 7760 37812
rect 7816 37756 7841 37812
rect 7897 37756 7922 37812
rect 7978 37756 8003 37812
rect 8059 37756 8084 37812
rect 8140 37756 8165 37812
rect 8221 37756 8246 37812
rect 8302 37756 8327 37812
rect 8383 37756 8408 37812
rect 8464 37756 8489 37812
rect 8545 37756 8570 37812
rect 8626 37756 8651 37812
rect 8707 37756 8732 37812
rect 8788 37756 8813 37812
rect 8869 37756 8894 37812
rect 8950 37756 8975 37812
rect 9031 37756 9056 37812
rect 9112 37756 9137 37812
rect 9193 37756 9218 37812
rect 9274 37756 9299 37812
rect 9355 37756 9380 37812
rect 9436 37756 9461 37812
rect 9517 37756 9542 37812
rect 7589 37732 9542 37756
rect 7589 37676 7598 37732
rect 7654 37676 7679 37732
rect 7735 37676 7760 37732
rect 7816 37676 7841 37732
rect 7897 37676 7922 37732
rect 7978 37676 8003 37732
rect 8059 37676 8084 37732
rect 8140 37676 8165 37732
rect 8221 37676 8246 37732
rect 8302 37676 8327 37732
rect 8383 37676 8408 37732
rect 8464 37676 8489 37732
rect 8545 37676 8570 37732
rect 8626 37676 8651 37732
rect 8707 37676 8732 37732
rect 8788 37676 8813 37732
rect 8869 37676 8894 37732
rect 8950 37676 8975 37732
rect 9031 37676 9056 37732
rect 9112 37676 9137 37732
rect 9193 37676 9218 37732
rect 9274 37676 9299 37732
rect 9355 37676 9380 37732
rect 9436 37676 9461 37732
rect 9517 37676 9542 37732
rect 7589 37652 9542 37676
rect 7589 37596 7598 37652
rect 7654 37596 7679 37652
rect 7735 37596 7760 37652
rect 7816 37596 7841 37652
rect 7897 37596 7922 37652
rect 7978 37596 8003 37652
rect 8059 37596 8084 37652
rect 8140 37596 8165 37652
rect 8221 37596 8246 37652
rect 8302 37596 8327 37652
rect 8383 37596 8408 37652
rect 8464 37596 8489 37652
rect 8545 37596 8570 37652
rect 8626 37596 8651 37652
rect 8707 37596 8732 37652
rect 8788 37596 8813 37652
rect 8869 37596 8894 37652
rect 8950 37596 8975 37652
rect 9031 37596 9056 37652
rect 9112 37596 9137 37652
rect 9193 37596 9218 37652
rect 9274 37596 9299 37652
rect 9355 37596 9380 37652
rect 9436 37596 9461 37652
rect 9517 37596 9542 37652
rect 7589 37572 9542 37596
rect 7589 37516 7598 37572
rect 7654 37516 7679 37572
rect 7735 37516 7760 37572
rect 7816 37516 7841 37572
rect 7897 37516 7922 37572
rect 7978 37516 8003 37572
rect 8059 37516 8084 37572
rect 8140 37516 8165 37572
rect 8221 37516 8246 37572
rect 8302 37516 8327 37572
rect 8383 37516 8408 37572
rect 8464 37516 8489 37572
rect 8545 37516 8570 37572
rect 8626 37516 8651 37572
rect 8707 37516 8732 37572
rect 8788 37516 8813 37572
rect 8869 37516 8894 37572
rect 8950 37516 8975 37572
rect 9031 37516 9056 37572
rect 9112 37516 9137 37572
rect 9193 37516 9218 37572
rect 9274 37516 9299 37572
rect 9355 37516 9380 37572
rect 9436 37516 9461 37572
rect 9517 37516 9542 37572
rect 7589 37492 9542 37516
rect 7589 37436 7598 37492
rect 7654 37436 7679 37492
rect 7735 37436 7760 37492
rect 7816 37436 7841 37492
rect 7897 37436 7922 37492
rect 7978 37436 8003 37492
rect 8059 37436 8084 37492
rect 8140 37436 8165 37492
rect 8221 37436 8246 37492
rect 8302 37436 8327 37492
rect 8383 37436 8408 37492
rect 8464 37436 8489 37492
rect 8545 37436 8570 37492
rect 8626 37436 8651 37492
rect 8707 37436 8732 37492
rect 8788 37436 8813 37492
rect 8869 37436 8894 37492
rect 8950 37436 8975 37492
rect 9031 37436 9056 37492
rect 9112 37436 9137 37492
rect 9193 37436 9218 37492
rect 9274 37436 9299 37492
rect 9355 37436 9380 37492
rect 9436 37436 9461 37492
rect 9517 37436 9542 37492
rect 7589 37412 9542 37436
rect 7589 37356 7598 37412
rect 7654 37356 7679 37412
rect 7735 37356 7760 37412
rect 7816 37356 7841 37412
rect 7897 37356 7922 37412
rect 7978 37356 8003 37412
rect 8059 37356 8084 37412
rect 8140 37356 8165 37412
rect 8221 37356 8246 37412
rect 8302 37356 8327 37412
rect 8383 37356 8408 37412
rect 8464 37356 8489 37412
rect 8545 37356 8570 37412
rect 8626 37356 8651 37412
rect 8707 37356 8732 37412
rect 8788 37356 8813 37412
rect 8869 37356 8894 37412
rect 8950 37356 8975 37412
rect 9031 37356 9056 37412
rect 9112 37356 9137 37412
rect 9193 37356 9218 37412
rect 9274 37356 9299 37412
rect 9355 37356 9380 37412
rect 9436 37356 9461 37412
rect 9517 37356 9542 37412
rect 7589 37332 9542 37356
rect 7589 37276 7598 37332
rect 7654 37276 7679 37332
rect 7735 37276 7760 37332
rect 7816 37276 7841 37332
rect 7897 37276 7922 37332
rect 7978 37276 8003 37332
rect 8059 37276 8084 37332
rect 8140 37276 8165 37332
rect 8221 37276 8246 37332
rect 8302 37276 8327 37332
rect 8383 37276 8408 37332
rect 8464 37276 8489 37332
rect 8545 37276 8570 37332
rect 8626 37276 8651 37332
rect 8707 37276 8732 37332
rect 8788 37276 8813 37332
rect 8869 37276 8894 37332
rect 8950 37276 8975 37332
rect 9031 37276 9056 37332
rect 9112 37276 9137 37332
rect 9193 37276 9218 37332
rect 9274 37276 9299 37332
rect 9355 37276 9380 37332
rect 9436 37276 9461 37332
rect 9517 37276 9542 37332
rect 7589 37252 9542 37276
rect 7589 37196 7598 37252
rect 7654 37196 7679 37252
rect 7735 37196 7760 37252
rect 7816 37196 7841 37252
rect 7897 37196 7922 37252
rect 7978 37196 8003 37252
rect 8059 37196 8084 37252
rect 8140 37196 8165 37252
rect 8221 37196 8246 37252
rect 8302 37196 8327 37252
rect 8383 37196 8408 37252
rect 8464 37196 8489 37252
rect 8545 37196 8570 37252
rect 8626 37196 8651 37252
rect 8707 37196 8732 37252
rect 8788 37196 8813 37252
rect 8869 37196 8894 37252
rect 8950 37196 8975 37252
rect 9031 37196 9056 37252
rect 9112 37196 9137 37252
rect 9193 37196 9218 37252
rect 9274 37196 9299 37252
rect 9355 37196 9380 37252
rect 9436 37196 9461 37252
rect 9517 37196 9542 37252
rect 7589 37172 9542 37196
rect 7589 37116 7598 37172
rect 7654 37116 7679 37172
rect 7735 37116 7760 37172
rect 7816 37116 7841 37172
rect 7897 37116 7922 37172
rect 7978 37116 8003 37172
rect 8059 37116 8084 37172
rect 8140 37116 8165 37172
rect 8221 37116 8246 37172
rect 8302 37116 8327 37172
rect 8383 37116 8408 37172
rect 8464 37116 8489 37172
rect 8545 37116 8570 37172
rect 8626 37116 8651 37172
rect 8707 37116 8732 37172
rect 8788 37116 8813 37172
rect 8869 37116 8894 37172
rect 8950 37116 8975 37172
rect 9031 37116 9056 37172
rect 9112 37116 9137 37172
rect 9193 37116 9218 37172
rect 9274 37116 9299 37172
rect 9355 37116 9380 37172
rect 9436 37116 9461 37172
rect 9517 37116 9542 37172
rect 7589 37092 9542 37116
rect 7589 37036 7598 37092
rect 7654 37036 7679 37092
rect 7735 37036 7760 37092
rect 7816 37036 7841 37092
rect 7897 37036 7922 37092
rect 7978 37036 8003 37092
rect 8059 37036 8084 37092
rect 8140 37036 8165 37092
rect 8221 37036 8246 37092
rect 8302 37036 8327 37092
rect 8383 37036 8408 37092
rect 8464 37036 8489 37092
rect 8545 37036 8570 37092
rect 8626 37036 8651 37092
rect 8707 37036 8732 37092
rect 8788 37036 8813 37092
rect 8869 37036 8894 37092
rect 8950 37036 8975 37092
rect 9031 37036 9056 37092
rect 9112 37036 9137 37092
rect 9193 37036 9218 37092
rect 9274 37036 9299 37092
rect 9355 37036 9380 37092
rect 9436 37036 9461 37092
rect 9517 37036 9542 37092
rect 9758 37036 9767 37892
rect 7589 35877 9767 37036
rect 7589 35821 7598 35877
rect 7654 35821 7678 35877
rect 7734 35821 7759 35877
rect 7815 35821 7840 35877
rect 7896 35821 7921 35877
rect 7977 35821 8002 35877
rect 8058 35821 8083 35877
rect 8139 35821 8164 35877
rect 8220 35821 8245 35877
rect 8301 35821 8326 35877
rect 8382 35821 8407 35877
rect 8463 35821 8488 35877
rect 8544 35821 8569 35877
rect 8625 35821 8650 35877
rect 8706 35821 8731 35877
rect 8787 35821 8812 35877
rect 8868 35821 8893 35877
rect 8949 35821 8974 35877
rect 9030 35821 9055 35877
rect 9111 35821 9136 35877
rect 9192 35821 9217 35877
rect 9273 35821 9298 35877
rect 9354 35821 9379 35877
rect 9435 35821 9460 35877
rect 9516 35821 9541 35877
rect 9597 35821 9622 35877
rect 9678 35821 9703 35877
rect 9759 35821 9767 35877
rect 7589 35789 9767 35821
rect 7589 35733 7598 35789
rect 7654 35733 7678 35789
rect 7734 35733 7759 35789
rect 7815 35733 7840 35789
rect 7896 35733 7921 35789
rect 7977 35733 8002 35789
rect 8058 35733 8083 35789
rect 8139 35733 8164 35789
rect 8220 35733 8245 35789
rect 8301 35733 8326 35789
rect 8382 35733 8407 35789
rect 8463 35733 8488 35789
rect 8544 35733 8569 35789
rect 8625 35733 8650 35789
rect 8706 35733 8731 35789
rect 8787 35733 8812 35789
rect 8868 35733 8893 35789
rect 8949 35733 8974 35789
rect 9030 35733 9055 35789
rect 9111 35733 9136 35789
rect 9192 35733 9217 35789
rect 9273 35733 9298 35789
rect 9354 35733 9379 35789
rect 9435 35733 9460 35789
rect 9516 35733 9541 35789
rect 9597 35733 9622 35789
rect 9678 35733 9703 35789
rect 9759 35733 9767 35789
rect 7589 35701 9767 35733
rect 7589 35645 7598 35701
rect 7654 35645 7678 35701
rect 7734 35645 7759 35701
rect 7815 35645 7840 35701
rect 7896 35645 7921 35701
rect 7977 35645 8002 35701
rect 8058 35645 8083 35701
rect 8139 35645 8164 35701
rect 8220 35645 8245 35701
rect 8301 35645 8326 35701
rect 8382 35645 8407 35701
rect 8463 35645 8488 35701
rect 8544 35645 8569 35701
rect 8625 35645 8650 35701
rect 8706 35645 8731 35701
rect 8787 35645 8812 35701
rect 8868 35645 8893 35701
rect 8949 35645 8974 35701
rect 9030 35645 9055 35701
rect 9111 35645 9136 35701
rect 9192 35645 9217 35701
rect 9273 35645 9298 35701
rect 9354 35645 9379 35701
rect 9435 35645 9460 35701
rect 9516 35645 9541 35701
rect 9597 35645 9622 35701
rect 9678 35645 9703 35701
rect 9759 35645 9767 35701
rect 7589 35613 9767 35645
rect 7589 35557 7598 35613
rect 7654 35557 7678 35613
rect 7734 35557 7759 35613
rect 7815 35557 7840 35613
rect 7896 35557 7921 35613
rect 7977 35557 8002 35613
rect 8058 35557 8083 35613
rect 8139 35557 8164 35613
rect 8220 35557 8245 35613
rect 8301 35557 8326 35613
rect 8382 35557 8407 35613
rect 8463 35557 8488 35613
rect 8544 35557 8569 35613
rect 8625 35557 8650 35613
rect 8706 35557 8731 35613
rect 8787 35557 8812 35613
rect 8868 35557 8893 35613
rect 8949 35557 8974 35613
rect 9030 35557 9055 35613
rect 9111 35557 9136 35613
rect 9192 35557 9217 35613
rect 9273 35557 9298 35613
rect 9354 35557 9379 35613
rect 9435 35557 9460 35613
rect 9516 35557 9541 35613
rect 9597 35557 9622 35613
rect 9678 35557 9703 35613
rect 9759 35557 9767 35613
rect 7589 35525 9767 35557
rect 7589 35469 7598 35525
rect 7654 35469 7678 35525
rect 7734 35469 7759 35525
rect 7815 35469 7840 35525
rect 7896 35469 7921 35525
rect 7977 35469 8002 35525
rect 8058 35469 8083 35525
rect 8139 35469 8164 35525
rect 8220 35469 8245 35525
rect 8301 35469 8326 35525
rect 8382 35469 8407 35525
rect 8463 35469 8488 35525
rect 8544 35469 8569 35525
rect 8625 35469 8650 35525
rect 8706 35469 8731 35525
rect 8787 35469 8812 35525
rect 8868 35469 8893 35525
rect 8949 35469 8974 35525
rect 9030 35469 9055 35525
rect 9111 35469 9136 35525
rect 9192 35469 9217 35525
rect 9273 35469 9298 35525
rect 9354 35469 9379 35525
rect 9435 35469 9460 35525
rect 9516 35469 9541 35525
rect 9597 35469 9622 35525
rect 9678 35469 9703 35525
rect 9759 35469 9767 35525
rect 7589 35437 9767 35469
rect 7589 35381 7598 35437
rect 7654 35381 7678 35437
rect 7734 35381 7759 35437
rect 7815 35381 7840 35437
rect 7896 35381 7921 35437
rect 7977 35381 8002 35437
rect 8058 35381 8083 35437
rect 8139 35381 8164 35437
rect 8220 35381 8245 35437
rect 8301 35381 8326 35437
rect 8382 35381 8407 35437
rect 8463 35381 8488 35437
rect 8544 35381 8569 35437
rect 8625 35381 8650 35437
rect 8706 35381 8731 35437
rect 8787 35381 8812 35437
rect 8868 35381 8893 35437
rect 8949 35381 8974 35437
rect 9030 35381 9055 35437
rect 9111 35381 9136 35437
rect 9192 35381 9217 35437
rect 9273 35381 9298 35437
rect 9354 35381 9379 35437
rect 9435 35381 9460 35437
rect 9516 35381 9541 35437
rect 9597 35381 9622 35437
rect 9678 35381 9703 35437
rect 9759 35381 9767 35437
rect 7589 33881 9767 35381
rect 7589 33858 7838 33881
rect 7589 33805 7636 33858
tri 7589 33802 7592 33805 ne
rect 7592 33802 7636 33805
rect 7692 33802 7716 33858
rect 7772 33825 7838 33858
rect 7894 33825 7922 33881
rect 7978 33878 9767 33881
rect 7978 33825 8041 33878
rect 7772 33822 8041 33825
rect 8097 33822 8124 33878
rect 8180 33822 8207 33878
rect 8263 33822 8290 33878
rect 8346 33822 8373 33878
rect 8429 33822 8456 33878
rect 8512 33822 8539 33878
rect 8595 33822 8622 33878
rect 8678 33822 8705 33878
rect 8761 33822 8788 33878
rect 8844 33822 8871 33878
rect 8927 33822 8954 33878
rect 9010 33822 9037 33878
rect 9093 33822 9120 33878
rect 9176 33822 9203 33878
rect 9259 33822 9286 33878
rect 9342 33822 9369 33878
rect 9425 33822 9452 33878
rect 9508 33822 9535 33878
rect 9591 33822 9618 33878
rect 9674 33822 9702 33878
rect 9758 33822 9767 33878
rect 7772 33802 9767 33822
tri 7592 33790 7604 33802 ne
rect 7604 33790 9767 33802
rect 4612 33748 4644 33790
rect 4502 33743 4644 33748
tri 4644 33743 4691 33790 nw
rect 4502 33734 4635 33743
tri 4635 33734 4644 33743 nw
rect 5207 33734 5216 33790
rect 5272 33734 5299 33790
rect 5355 33734 5382 33790
rect 5438 33734 5465 33790
rect 5521 33734 5548 33790
rect 5604 33734 5631 33790
rect 5687 33734 5714 33790
rect 5770 33734 5797 33790
rect 5853 33734 5880 33790
rect 5936 33734 5963 33790
rect 6019 33734 6046 33790
rect 6102 33734 6129 33790
rect 6185 33734 6211 33790
rect 6267 33734 6293 33790
rect 6349 33734 6375 33790
rect 6431 33734 6457 33790
rect 6513 33734 6539 33790
rect 6595 33734 6621 33790
rect 6677 33734 6703 33790
rect 6759 33734 6785 33790
rect 6841 33734 6867 33790
rect 6923 33734 6949 33790
rect 7005 33734 7031 33790
rect 7087 33734 7113 33790
rect 7169 33734 7195 33790
rect 7251 33734 7385 33790
tri 7604 33776 7618 33790 ne
rect 7618 33776 8041 33790
tri 7618 33766 7628 33776 ne
rect 7628 33766 8041 33776
tri 7628 33756 7638 33766 ne
rect 7638 33756 7838 33766
tri 7638 33751 7643 33756 ne
rect 7643 33751 7838 33756
rect 4502 33724 4603 33734
rect 3121 33708 4603 33724
rect 3121 33652 3513 33708
rect 3569 33652 3594 33708
rect 3650 33652 3675 33708
rect 3731 33652 3757 33708
rect 3813 33652 3839 33708
rect 3895 33652 3921 33708
rect 3977 33652 4003 33708
rect 4059 33652 4085 33708
rect 4141 33652 4167 33708
rect 4223 33652 4249 33708
rect 4305 33702 4603 33708
tri 4603 33702 4635 33734 nw
rect 5207 33702 7385 33734
rect 4305 33679 4547 33702
rect 4305 33652 4354 33679
rect 3121 33623 4354 33652
rect 4410 33623 4446 33679
rect 4502 33646 4547 33679
tri 4547 33646 4603 33702 nw
rect 5207 33646 5216 33702
rect 5272 33646 5299 33702
rect 5355 33646 5382 33702
rect 5438 33646 5465 33702
rect 5521 33646 5548 33702
rect 5604 33646 5631 33702
rect 5687 33646 5714 33702
rect 5770 33646 5797 33702
rect 5853 33646 5880 33702
rect 5936 33646 5963 33702
rect 6019 33646 6046 33702
rect 6102 33646 6129 33702
rect 6185 33646 6211 33702
rect 6267 33646 6293 33702
rect 6349 33646 6375 33702
rect 6431 33646 6457 33702
rect 6513 33646 6539 33702
rect 6595 33646 6621 33702
rect 6677 33646 6703 33702
rect 6759 33646 6785 33702
rect 6841 33646 6867 33702
rect 6923 33646 6949 33702
rect 7005 33646 7031 33702
rect 7087 33646 7113 33702
rect 7169 33646 7195 33702
rect 7251 33646 7385 33702
tri 7643 33695 7699 33751 ne
rect 7699 33695 7723 33751
rect 7779 33710 7838 33751
rect 7894 33710 7922 33766
rect 7978 33734 8041 33766
rect 8097 33734 8124 33790
rect 8180 33734 8207 33790
rect 8263 33734 8290 33790
rect 8346 33734 8373 33790
rect 8429 33734 8456 33790
rect 8512 33734 8539 33790
rect 8595 33734 8622 33790
rect 8678 33734 8705 33790
rect 8761 33734 8788 33790
rect 8844 33734 8871 33790
rect 8927 33734 8954 33790
rect 9010 33734 9037 33790
rect 9093 33734 9120 33790
rect 9176 33734 9203 33790
rect 9259 33734 9286 33790
rect 9342 33734 9369 33790
rect 9425 33734 9452 33790
rect 9508 33734 9535 33790
rect 9591 33734 9618 33790
rect 9674 33734 9702 33790
rect 9758 33734 9767 33790
rect 9974 37892 12066 37903
rect 9974 37836 9983 37892
rect 10039 37836 10064 37892
rect 10120 37836 10145 37892
rect 10201 37836 10226 37892
rect 10282 37836 10307 37892
rect 10363 37836 10388 37892
rect 10444 37836 10469 37892
rect 10525 37836 10550 37892
rect 10606 37836 10631 37892
rect 10687 37836 10712 37892
rect 10768 37836 10793 37892
rect 10849 37836 10874 37892
rect 10930 37836 10955 37892
rect 11011 37836 11036 37892
rect 11092 37836 11117 37892
rect 11173 37836 11198 37892
rect 11254 37836 11279 37892
rect 11335 37836 11360 37892
rect 11416 37836 11441 37892
rect 9974 37812 11441 37836
rect 9974 37756 9983 37812
rect 10039 37756 10064 37812
rect 10120 37756 10145 37812
rect 10201 37756 10226 37812
rect 10282 37756 10307 37812
rect 10363 37756 10388 37812
rect 10444 37756 10469 37812
rect 10525 37756 10550 37812
rect 10606 37756 10631 37812
rect 10687 37756 10712 37812
rect 10768 37756 10793 37812
rect 10849 37756 10874 37812
rect 10930 37756 10955 37812
rect 11011 37756 11036 37812
rect 11092 37756 11117 37812
rect 11173 37756 11198 37812
rect 11254 37756 11279 37812
rect 11335 37756 11360 37812
rect 11416 37756 11441 37812
rect 9974 37732 11441 37756
rect 9974 37676 9983 37732
rect 10039 37676 10064 37732
rect 10120 37676 10145 37732
rect 10201 37676 10226 37732
rect 10282 37676 10307 37732
rect 10363 37676 10388 37732
rect 10444 37676 10469 37732
rect 10525 37676 10550 37732
rect 10606 37676 10631 37732
rect 10687 37676 10712 37732
rect 10768 37676 10793 37732
rect 10849 37676 10874 37732
rect 10930 37676 10955 37732
rect 11011 37676 11036 37732
rect 11092 37676 11117 37732
rect 11173 37676 11198 37732
rect 11254 37676 11279 37732
rect 11335 37676 11360 37732
rect 11416 37676 11441 37732
rect 9974 37652 11441 37676
rect 9974 37596 9983 37652
rect 10039 37596 10064 37652
rect 10120 37596 10145 37652
rect 10201 37596 10226 37652
rect 10282 37596 10307 37652
rect 10363 37596 10388 37652
rect 10444 37596 10469 37652
rect 10525 37596 10550 37652
rect 10606 37596 10631 37652
rect 10687 37596 10712 37652
rect 10768 37596 10793 37652
rect 10849 37596 10874 37652
rect 10930 37596 10955 37652
rect 11011 37596 11036 37652
rect 11092 37596 11117 37652
rect 11173 37596 11198 37652
rect 11254 37596 11279 37652
rect 11335 37596 11360 37652
rect 11416 37596 11441 37652
rect 9974 37572 11441 37596
rect 9974 37516 9983 37572
rect 10039 37516 10064 37572
rect 10120 37516 10145 37572
rect 10201 37516 10226 37572
rect 10282 37516 10307 37572
rect 10363 37516 10388 37572
rect 10444 37516 10469 37572
rect 10525 37516 10550 37572
rect 10606 37516 10631 37572
rect 10687 37516 10712 37572
rect 10768 37516 10793 37572
rect 10849 37516 10874 37572
rect 10930 37516 10955 37572
rect 11011 37516 11036 37572
rect 11092 37516 11117 37572
rect 11173 37516 11198 37572
rect 11254 37516 11279 37572
rect 11335 37516 11360 37572
rect 11416 37516 11441 37572
rect 9974 37492 11441 37516
rect 9974 37436 9983 37492
rect 10039 37436 10064 37492
rect 10120 37436 10145 37492
rect 10201 37436 10226 37492
rect 10282 37436 10307 37492
rect 10363 37436 10388 37492
rect 10444 37436 10469 37492
rect 10525 37436 10550 37492
rect 10606 37436 10631 37492
rect 10687 37436 10712 37492
rect 10768 37436 10793 37492
rect 10849 37436 10874 37492
rect 10930 37436 10955 37492
rect 11011 37436 11036 37492
rect 11092 37436 11117 37492
rect 11173 37436 11198 37492
rect 11254 37436 11279 37492
rect 11335 37436 11360 37492
rect 11416 37436 11441 37492
rect 9974 37412 11441 37436
rect 9974 37356 9983 37412
rect 10039 37356 10064 37412
rect 10120 37356 10145 37412
rect 10201 37356 10226 37412
rect 10282 37356 10307 37412
rect 10363 37356 10388 37412
rect 10444 37356 10469 37412
rect 10525 37356 10550 37412
rect 10606 37356 10631 37412
rect 10687 37356 10712 37412
rect 10768 37356 10793 37412
rect 10849 37356 10874 37412
rect 10930 37356 10955 37412
rect 11011 37356 11036 37412
rect 11092 37356 11117 37412
rect 11173 37356 11198 37412
rect 11254 37356 11279 37412
rect 11335 37356 11360 37412
rect 11416 37356 11441 37412
rect 9974 37332 11441 37356
rect 9974 37276 9983 37332
rect 10039 37276 10064 37332
rect 10120 37276 10145 37332
rect 10201 37276 10226 37332
rect 10282 37276 10307 37332
rect 10363 37276 10388 37332
rect 10444 37276 10469 37332
rect 10525 37276 10550 37332
rect 10606 37276 10631 37332
rect 10687 37276 10712 37332
rect 10768 37276 10793 37332
rect 10849 37276 10874 37332
rect 10930 37276 10955 37332
rect 11011 37276 11036 37332
rect 11092 37276 11117 37332
rect 11173 37276 11198 37332
rect 11254 37276 11279 37332
rect 11335 37276 11360 37332
rect 11416 37276 11441 37332
rect 9974 37252 11441 37276
rect 9974 37196 9983 37252
rect 10039 37196 10064 37252
rect 10120 37196 10145 37252
rect 10201 37196 10226 37252
rect 10282 37196 10307 37252
rect 10363 37196 10388 37252
rect 10444 37196 10469 37252
rect 10525 37196 10550 37252
rect 10606 37196 10631 37252
rect 10687 37196 10712 37252
rect 10768 37196 10793 37252
rect 10849 37196 10874 37252
rect 10930 37196 10955 37252
rect 11011 37196 11036 37252
rect 11092 37196 11117 37252
rect 11173 37196 11198 37252
rect 11254 37196 11279 37252
rect 11335 37196 11360 37252
rect 11416 37196 11441 37252
rect 9974 37172 11441 37196
rect 9974 37116 9983 37172
rect 10039 37116 10064 37172
rect 10120 37116 10145 37172
rect 10201 37116 10226 37172
rect 10282 37116 10307 37172
rect 10363 37116 10388 37172
rect 10444 37116 10469 37172
rect 10525 37116 10550 37172
rect 10606 37116 10631 37172
rect 10687 37116 10712 37172
rect 10768 37116 10793 37172
rect 10849 37116 10874 37172
rect 10930 37116 10955 37172
rect 11011 37116 11036 37172
rect 11092 37116 11117 37172
rect 11173 37116 11198 37172
rect 11254 37116 11279 37172
rect 11335 37116 11360 37172
rect 11416 37116 11441 37172
rect 9974 37092 11441 37116
rect 9974 37036 9983 37092
rect 10039 37036 10064 37092
rect 10120 37036 10145 37092
rect 10201 37036 10226 37092
rect 10282 37036 10307 37092
rect 10363 37036 10388 37092
rect 10444 37036 10469 37092
rect 10525 37036 10550 37092
rect 10606 37036 10631 37092
rect 10687 37036 10712 37092
rect 10768 37036 10793 37092
rect 10849 37036 10874 37092
rect 10930 37036 10955 37092
rect 11011 37036 11036 37092
rect 11092 37036 11117 37092
rect 11173 37036 11198 37092
rect 11254 37036 11279 37092
rect 11335 37036 11360 37092
rect 11416 37036 11441 37092
rect 12057 37036 12066 37892
rect 9974 35877 12066 37036
rect 9974 35821 9983 35877
rect 10039 35821 10063 35877
rect 10119 35821 10143 35877
rect 10199 35821 10223 35877
rect 10279 35821 10303 35877
rect 10359 35821 10383 35877
rect 10439 35821 10463 35877
rect 10519 35821 10544 35877
rect 10600 35821 10625 35877
rect 10681 35821 10706 35877
rect 10762 35821 10787 35877
rect 10843 35821 10868 35877
rect 10924 35821 10949 35877
rect 11005 35821 11030 35877
rect 11086 35821 11111 35877
rect 11167 35821 11192 35877
rect 11248 35821 11273 35877
rect 11329 35821 11354 35877
rect 11410 35821 11435 35877
rect 11491 35821 11516 35877
rect 11572 35821 11597 35877
rect 11653 35821 11678 35877
rect 11734 35821 11759 35877
rect 11815 35821 11840 35877
rect 11896 35821 11921 35877
rect 11977 35821 12002 35877
rect 12058 35821 12066 35877
rect 9974 35789 12066 35821
rect 9974 35733 9983 35789
rect 10039 35733 10063 35789
rect 10119 35733 10143 35789
rect 10199 35733 10223 35789
rect 10279 35733 10303 35789
rect 10359 35733 10383 35789
rect 10439 35733 10463 35789
rect 10519 35733 10544 35789
rect 10600 35733 10625 35789
rect 10681 35733 10706 35789
rect 10762 35733 10787 35789
rect 10843 35733 10868 35789
rect 10924 35733 10949 35789
rect 11005 35733 11030 35789
rect 11086 35733 11111 35789
rect 11167 35733 11192 35789
rect 11248 35733 11273 35789
rect 11329 35733 11354 35789
rect 11410 35733 11435 35789
rect 11491 35733 11516 35789
rect 11572 35733 11597 35789
rect 11653 35733 11678 35789
rect 11734 35733 11759 35789
rect 11815 35733 11840 35789
rect 11896 35733 11921 35789
rect 11977 35733 12002 35789
rect 12058 35733 12066 35789
rect 9974 35701 12066 35733
rect 9974 35645 9983 35701
rect 10039 35645 10063 35701
rect 10119 35645 10143 35701
rect 10199 35645 10223 35701
rect 10279 35645 10303 35701
rect 10359 35645 10383 35701
rect 10439 35645 10463 35701
rect 10519 35645 10544 35701
rect 10600 35645 10625 35701
rect 10681 35645 10706 35701
rect 10762 35645 10787 35701
rect 10843 35645 10868 35701
rect 10924 35645 10949 35701
rect 11005 35645 11030 35701
rect 11086 35645 11111 35701
rect 11167 35645 11192 35701
rect 11248 35645 11273 35701
rect 11329 35645 11354 35701
rect 11410 35645 11435 35701
rect 11491 35645 11516 35701
rect 11572 35645 11597 35701
rect 11653 35645 11678 35701
rect 11734 35645 11759 35701
rect 11815 35645 11840 35701
rect 11896 35645 11921 35701
rect 11977 35645 12002 35701
rect 12058 35645 12066 35701
rect 9974 35613 12066 35645
rect 9974 35557 9983 35613
rect 10039 35557 10063 35613
rect 10119 35557 10143 35613
rect 10199 35557 10223 35613
rect 10279 35557 10303 35613
rect 10359 35557 10383 35613
rect 10439 35557 10463 35613
rect 10519 35557 10544 35613
rect 10600 35557 10625 35613
rect 10681 35557 10706 35613
rect 10762 35557 10787 35613
rect 10843 35557 10868 35613
rect 10924 35557 10949 35613
rect 11005 35557 11030 35613
rect 11086 35557 11111 35613
rect 11167 35557 11192 35613
rect 11248 35557 11273 35613
rect 11329 35557 11354 35613
rect 11410 35557 11435 35613
rect 11491 35557 11516 35613
rect 11572 35557 11597 35613
rect 11653 35557 11678 35613
rect 11734 35557 11759 35613
rect 11815 35557 11840 35613
rect 11896 35557 11921 35613
rect 11977 35557 12002 35613
rect 12058 35557 12066 35613
rect 9974 35525 12066 35557
rect 9974 35469 9983 35525
rect 10039 35469 10063 35525
rect 10119 35469 10143 35525
rect 10199 35469 10223 35525
rect 10279 35469 10303 35525
rect 10359 35469 10383 35525
rect 10439 35469 10463 35525
rect 10519 35469 10544 35525
rect 10600 35469 10625 35525
rect 10681 35469 10706 35525
rect 10762 35469 10787 35525
rect 10843 35469 10868 35525
rect 10924 35469 10949 35525
rect 11005 35469 11030 35525
rect 11086 35469 11111 35525
rect 11167 35469 11192 35525
rect 11248 35469 11273 35525
rect 11329 35469 11354 35525
rect 11410 35469 11435 35525
rect 11491 35469 11516 35525
rect 11572 35469 11597 35525
rect 11653 35469 11678 35525
rect 11734 35469 11759 35525
rect 11815 35469 11840 35525
rect 11896 35469 11921 35525
rect 11977 35469 12002 35525
rect 12058 35469 12066 35525
rect 9974 35437 12066 35469
rect 9974 35381 9983 35437
rect 10039 35381 10063 35437
rect 10119 35381 10143 35437
rect 10199 35381 10223 35437
rect 10279 35381 10303 35437
rect 10359 35381 10383 35437
rect 10439 35381 10463 35437
rect 10519 35381 10544 35437
rect 10600 35381 10625 35437
rect 10681 35381 10706 35437
rect 10762 35381 10787 35437
rect 10843 35381 10868 35437
rect 10924 35381 10949 35437
rect 11005 35381 11030 35437
rect 11086 35381 11111 35437
rect 11167 35381 11192 35437
rect 11248 35381 11273 35437
rect 11329 35381 11354 35437
rect 11410 35381 11435 35437
rect 11491 35381 11516 35437
rect 11572 35381 11597 35437
rect 11653 35381 11678 35437
rect 11734 35381 11759 35437
rect 11815 35381 11840 35437
rect 11896 35381 11921 35437
rect 11977 35381 12002 35437
rect 12058 35381 12066 35437
rect 9974 33881 12066 35381
rect 9974 33858 10202 33881
rect 9974 33802 10000 33858
rect 10056 33802 10080 33858
rect 10136 33825 10202 33858
rect 10258 33825 10286 33881
rect 10342 33878 12066 33881
rect 10342 33825 10397 33878
rect 10136 33822 10397 33825
rect 10453 33822 10477 33878
rect 10533 33822 10557 33878
rect 10613 33822 10637 33878
rect 10693 33822 10717 33878
rect 10773 33822 10797 33878
rect 10853 33822 10877 33878
rect 10933 33822 10957 33878
rect 11013 33822 11037 33878
rect 11093 33822 11117 33878
rect 11173 33822 11197 33878
rect 11253 33822 11277 33878
rect 11333 33822 11357 33878
rect 11413 33822 11437 33878
rect 11493 33822 11517 33878
rect 11573 33822 11597 33878
rect 11653 33822 11677 33878
rect 11733 33822 11758 33878
rect 11814 33822 11839 33878
rect 11895 33822 11920 33878
rect 11976 33822 12001 33878
rect 12057 33822 12066 33878
rect 10136 33802 12066 33822
rect 9974 33790 12066 33802
rect 9974 33784 10397 33790
tri 9974 33776 9982 33784 ne
rect 9982 33776 10397 33784
tri 9982 33766 9992 33776 ne
rect 9992 33766 10397 33776
tri 9992 33756 10002 33766 ne
rect 10002 33756 10202 33766
tri 10002 33751 10007 33756 ne
rect 10007 33751 10202 33756
rect 7978 33710 9767 33734
rect 7779 33702 9767 33710
rect 7779 33695 8041 33702
tri 7699 33690 7704 33695 ne
rect 7704 33690 8041 33695
tri 7704 33650 7744 33690 ne
rect 7744 33650 8041 33690
rect 4502 33623 4519 33646
rect 3121 33618 4519 33623
tri 4519 33618 4547 33646 nw
rect 3121 33614 4515 33618
tri 4515 33614 4519 33618 nw
rect 5207 33614 7385 33646
rect 3121 33558 3513 33614
rect 3569 33558 3594 33614
rect 3650 33558 3675 33614
rect 3731 33558 3757 33614
rect 3813 33558 3839 33614
rect 3895 33558 3921 33614
rect 3977 33558 4003 33614
rect 4059 33558 4085 33614
rect 4141 33558 4167 33614
rect 4223 33558 4249 33614
rect 4305 33558 4459 33614
tri 4459 33558 4515 33614 nw
rect 5207 33558 5216 33614
rect 5272 33558 5299 33614
rect 5355 33558 5382 33614
rect 5438 33558 5465 33614
rect 5521 33558 5548 33614
rect 5604 33558 5631 33614
rect 5687 33558 5714 33614
rect 5770 33558 5797 33614
rect 5853 33558 5880 33614
rect 5936 33558 5963 33614
rect 6019 33558 6046 33614
rect 6102 33558 6129 33614
rect 6185 33558 6211 33614
rect 6267 33558 6293 33614
rect 6349 33558 6375 33614
rect 6431 33558 6457 33614
rect 6513 33558 6539 33614
rect 6595 33558 6621 33614
rect 6677 33558 6703 33614
rect 6759 33558 6785 33614
rect 6841 33558 6867 33614
rect 6923 33558 6949 33614
rect 7005 33558 7031 33614
rect 7087 33558 7113 33614
rect 7169 33558 7195 33614
rect 7251 33558 7385 33614
tri 7744 33594 7800 33650 ne
rect 7800 33594 7838 33650
rect 7894 33594 7922 33650
rect 7978 33646 8041 33650
rect 8097 33646 8124 33702
rect 8180 33646 8207 33702
rect 8263 33646 8290 33702
rect 8346 33646 8373 33702
rect 8429 33646 8456 33702
rect 8512 33646 8539 33702
rect 8595 33646 8622 33702
rect 8678 33646 8705 33702
rect 8761 33646 8788 33702
rect 8844 33646 8871 33702
rect 8927 33646 8954 33702
rect 9010 33646 9037 33702
rect 9093 33646 9120 33702
rect 9176 33646 9203 33702
rect 9259 33646 9286 33702
rect 9342 33646 9369 33702
rect 9425 33646 9452 33702
rect 9508 33646 9535 33702
rect 9591 33646 9618 33702
rect 9674 33646 9702 33702
rect 9758 33646 9767 33702
tri 10007 33695 10063 33751 ne
rect 10063 33695 10087 33751
rect 10143 33710 10202 33751
rect 10258 33710 10286 33766
rect 10342 33734 10397 33766
rect 10453 33734 10477 33790
rect 10533 33734 10557 33790
rect 10613 33734 10637 33790
rect 10693 33734 10717 33790
rect 10773 33734 10797 33790
rect 10853 33734 10877 33790
rect 10933 33734 10957 33790
rect 11013 33734 11037 33790
rect 11093 33734 11117 33790
rect 11173 33734 11197 33790
rect 11253 33734 11277 33790
rect 11333 33734 11357 33790
rect 11413 33734 11437 33790
rect 11493 33734 11517 33790
rect 11573 33734 11597 33790
rect 11653 33734 11677 33790
rect 11733 33734 11758 33790
rect 11814 33734 11839 33790
rect 11895 33734 11920 33790
rect 11976 33734 12001 33790
rect 12057 33734 12066 33790
rect 10342 33710 12066 33734
rect 10143 33702 12066 33710
rect 10143 33695 10397 33702
tri 10063 33690 10068 33695 ne
rect 10068 33690 10397 33695
tri 10068 33650 10108 33690 ne
rect 10108 33650 10397 33690
rect 7978 33614 9767 33646
rect 7978 33594 8041 33614
tri 7800 33589 7805 33594 ne
rect 7805 33589 8041 33594
tri 7805 33558 7836 33589 ne
rect 7836 33558 8041 33589
rect 8097 33558 8124 33614
rect 8180 33558 8207 33614
rect 8263 33558 8290 33614
rect 8346 33558 8373 33614
rect 8429 33558 8456 33614
rect 8512 33558 8539 33614
rect 8595 33558 8622 33614
rect 8678 33558 8705 33614
rect 8761 33558 8788 33614
rect 8844 33558 8871 33614
rect 8927 33558 8954 33614
rect 9010 33558 9037 33614
rect 9093 33558 9120 33614
rect 9176 33558 9203 33614
rect 9259 33558 9286 33614
rect 9342 33558 9369 33614
rect 9425 33558 9452 33614
rect 9508 33558 9535 33614
rect 9591 33558 9618 33614
rect 9674 33558 9702 33614
rect 9758 33558 9767 33614
tri 10108 33594 10164 33650 ne
rect 10164 33594 10202 33650
rect 10258 33594 10286 33650
rect 10342 33646 10397 33650
rect 10453 33646 10477 33702
rect 10533 33646 10557 33702
rect 10613 33646 10637 33702
rect 10693 33646 10717 33702
rect 10773 33646 10797 33702
rect 10853 33646 10877 33702
rect 10933 33646 10957 33702
rect 11013 33646 11037 33702
rect 11093 33646 11117 33702
rect 11173 33646 11197 33702
rect 11253 33646 11277 33702
rect 11333 33646 11357 33702
rect 11413 33646 11437 33702
rect 11493 33646 11517 33702
rect 11573 33646 11597 33702
rect 11653 33646 11677 33702
rect 11733 33646 11758 33702
rect 11814 33646 11839 33702
rect 11895 33646 11920 33702
rect 11976 33646 12001 33702
rect 12057 33646 12066 33702
rect 10342 33614 12066 33646
rect 10342 33594 10397 33614
tri 10164 33589 10169 33594 ne
rect 10169 33589 10397 33594
tri 10169 33558 10200 33589 ne
rect 10200 33558 10397 33589
rect 10453 33558 10477 33614
rect 10533 33558 10557 33614
rect 10613 33558 10637 33614
rect 10693 33558 10717 33614
rect 10773 33558 10797 33614
rect 10853 33558 10877 33614
rect 10933 33558 10957 33614
rect 11013 33558 11037 33614
rect 11093 33558 11117 33614
rect 11173 33558 11197 33614
rect 11253 33558 11277 33614
rect 11333 33558 11357 33614
rect 11413 33558 11437 33614
rect 11493 33558 11517 33614
rect 11573 33558 11597 33614
rect 11653 33558 11677 33614
rect 11733 33558 11758 33614
rect 11814 33558 11839 33614
rect 11895 33558 11920 33614
rect 11976 33558 12001 33614
rect 12057 33558 12066 33614
rect 3121 33535 4436 33558
tri 4436 33535 4459 33558 nw
rect 3121 33526 4427 33535
tri 4427 33526 4436 33535 nw
rect 5207 33526 7385 33558
tri 7836 33540 7854 33558 ne
rect 7854 33540 9767 33558
tri 10200 33540 10218 33558 ne
rect 10218 33540 12066 33558
tri 7854 33535 7859 33540 ne
rect 7859 33535 9767 33540
tri 10218 33535 10223 33540 ne
rect 10223 33535 12066 33540
rect 3121 33520 4371 33526
rect 3121 33464 3513 33520
rect 3569 33464 3594 33520
rect 3650 33464 3675 33520
rect 3731 33464 3757 33520
rect 3813 33464 3839 33520
rect 3895 33464 3921 33520
rect 3977 33464 4003 33520
rect 4059 33464 4085 33520
rect 4141 33464 4167 33520
rect 4223 33464 4249 33520
rect 4305 33470 4371 33520
tri 4371 33470 4427 33526 nw
rect 5207 33470 5216 33526
rect 5272 33470 5299 33526
rect 5355 33470 5382 33526
rect 5438 33470 5465 33526
rect 5521 33470 5548 33526
rect 5604 33470 5631 33526
rect 5687 33470 5714 33526
rect 5770 33470 5797 33526
rect 5853 33470 5880 33526
rect 5936 33470 5963 33526
rect 6019 33470 6046 33526
rect 6102 33470 6129 33526
rect 6185 33470 6211 33526
rect 6267 33470 6293 33526
rect 6349 33470 6375 33526
rect 6431 33470 6457 33526
rect 6513 33470 6539 33526
rect 6595 33470 6621 33526
rect 6677 33470 6703 33526
rect 6759 33470 6785 33526
rect 6841 33470 6867 33526
rect 6923 33470 6949 33526
rect 7005 33470 7031 33526
rect 7087 33470 7113 33526
rect 7169 33470 7195 33526
rect 7251 33492 7385 33526
rect 7251 33479 7372 33492
tri 7372 33479 7385 33492 nw
tri 7859 33479 7915 33535 ne
rect 7915 33479 7943 33535
rect 7999 33526 9767 33535
rect 7999 33479 8041 33526
rect 7251 33470 7363 33479
tri 7363 33470 7372 33479 nw
tri 7915 33474 7920 33479 ne
rect 7920 33474 8041 33479
tri 7920 33470 7924 33474 ne
rect 7924 33470 8041 33474
rect 8097 33470 8124 33526
rect 8180 33470 8207 33526
rect 8263 33470 8290 33526
rect 8346 33470 8373 33526
rect 8429 33470 8456 33526
rect 8512 33470 8539 33526
rect 8595 33470 8622 33526
rect 8678 33470 8705 33526
rect 8761 33470 8788 33526
rect 8844 33470 8871 33526
rect 8927 33470 8954 33526
rect 9010 33470 9037 33526
rect 9093 33470 9120 33526
rect 9176 33470 9203 33526
rect 9259 33470 9286 33526
rect 9342 33470 9369 33526
rect 9425 33470 9452 33526
rect 9508 33470 9535 33526
rect 9591 33470 9618 33526
rect 9674 33470 9702 33526
rect 9758 33470 9767 33526
tri 10223 33479 10279 33535 ne
rect 10279 33479 10307 33535
rect 10363 33526 12066 33535
rect 10363 33479 10397 33526
tri 10279 33474 10284 33479 ne
rect 10284 33474 10397 33479
tri 10284 33470 10288 33474 ne
rect 10288 33470 10397 33474
rect 10453 33470 10477 33526
rect 10533 33470 10557 33526
rect 10613 33470 10637 33526
rect 10693 33470 10717 33526
rect 10773 33470 10797 33526
rect 10853 33470 10877 33526
rect 10933 33470 10957 33526
rect 11013 33470 11037 33526
rect 11093 33470 11117 33526
rect 11173 33470 11197 33526
rect 11253 33470 11277 33526
rect 11333 33470 11357 33526
rect 11413 33470 11437 33526
rect 11493 33470 11517 33526
rect 11573 33470 11597 33526
rect 11653 33470 11677 33526
rect 11733 33470 11758 33526
rect 11814 33470 11839 33526
rect 11895 33470 11920 33526
rect 11976 33470 12001 33526
rect 12057 33470 12066 33526
rect 4305 33464 4339 33470
rect 3121 33438 4339 33464
tri 4339 33438 4371 33470 nw
rect 5207 33438 7331 33470
tri 7331 33438 7363 33470 nw
tri 7924 33438 7956 33470 ne
rect 7956 33438 9767 33470
tri 10288 33438 10320 33470 ne
rect 10320 33438 12066 33470
rect 3121 33426 4321 33438
rect 3121 33370 3513 33426
rect 3569 33370 3594 33426
rect 3650 33370 3675 33426
rect 3731 33370 3757 33426
rect 3813 33370 3839 33426
rect 3895 33370 3921 33426
rect 3977 33370 4003 33426
rect 4059 33370 4085 33426
rect 4141 33370 4167 33426
rect 4223 33370 4249 33426
rect 4305 33370 4321 33426
tri 4321 33420 4339 33438 nw
rect 3121 31896 4321 33370
rect 3121 31840 3513 31896
rect 3569 31840 3596 31896
rect 3652 31840 3679 31896
rect 3735 31840 3762 31896
rect 3818 31840 3845 31896
rect 3901 31840 3928 31896
rect 3984 31840 4011 31896
rect 4067 31840 4094 31896
rect 4150 31840 4177 31896
rect 4233 31840 4260 31896
rect 4316 31840 4321 31896
rect 3121 31802 4321 31840
rect 3121 31746 3513 31802
rect 3569 31746 3596 31802
rect 3652 31746 3679 31802
rect 3735 31746 3762 31802
rect 3818 31746 3845 31802
rect 3901 31746 3928 31802
rect 3984 31746 4011 31802
rect 4067 31746 4094 31802
rect 4150 31746 4177 31802
rect 4233 31746 4260 31802
rect 4316 31746 4321 31802
rect 3121 31708 4321 31746
rect 3121 31652 3513 31708
rect 3569 31652 3596 31708
rect 3652 31652 3679 31708
rect 3735 31652 3762 31708
rect 3818 31652 3845 31708
rect 3901 31652 3928 31708
rect 3984 31652 4011 31708
rect 4067 31652 4094 31708
rect 4150 31652 4177 31708
rect 4233 31652 4260 31708
rect 4316 31652 4321 31708
rect 3121 31614 4321 31652
rect 3121 31558 3513 31614
rect 3569 31558 3596 31614
rect 3652 31558 3679 31614
rect 3735 31558 3762 31614
rect 3818 31558 3845 31614
rect 3901 31558 3928 31614
rect 3984 31558 4011 31614
rect 4067 31558 4094 31614
rect 4150 31558 4177 31614
rect 4233 31558 4260 31614
rect 4316 31558 4321 31614
rect 3121 31520 4321 31558
rect 3121 31464 3513 31520
rect 3569 31464 3596 31520
rect 3652 31464 3679 31520
rect 3735 31464 3762 31520
rect 3818 31464 3845 31520
rect 3901 31464 3928 31520
rect 3984 31464 4011 31520
rect 4067 31464 4094 31520
rect 4150 31464 4177 31520
rect 4233 31464 4260 31520
rect 4316 31464 4321 31520
rect 3121 31426 4321 31464
rect 3121 31370 3513 31426
rect 3569 31370 3596 31426
rect 3652 31370 3679 31426
rect 3735 31370 3762 31426
rect 3818 31370 3845 31426
rect 3901 31370 3928 31426
rect 3984 31370 4011 31426
rect 4067 31370 4094 31426
rect 4150 31370 4177 31426
rect 4233 31370 4260 31426
rect 4316 31370 4321 31426
rect 3121 29896 4321 31370
rect 3121 29840 3513 29896
rect 3569 29840 3596 29896
rect 3652 29840 3679 29896
rect 3735 29840 3762 29896
rect 3818 29840 3845 29896
rect 3901 29840 3928 29896
rect 3984 29840 4011 29896
rect 4067 29840 4094 29896
rect 4150 29840 4177 29896
rect 4233 29840 4260 29896
rect 4316 29840 4321 29896
rect 3121 29802 4321 29840
rect 3121 29746 3513 29802
rect 3569 29746 3596 29802
rect 3652 29746 3679 29802
rect 3735 29746 3762 29802
rect 3818 29746 3845 29802
rect 3901 29746 3928 29802
rect 3984 29746 4011 29802
rect 4067 29746 4094 29802
rect 4150 29746 4177 29802
rect 4233 29746 4260 29802
rect 4316 29746 4321 29802
rect 3121 29708 4321 29746
rect 3121 29652 3513 29708
rect 3569 29652 3596 29708
rect 3652 29652 3679 29708
rect 3735 29652 3762 29708
rect 3818 29652 3845 29708
rect 3901 29652 3928 29708
rect 3984 29652 4011 29708
rect 4067 29652 4094 29708
rect 4150 29652 4177 29708
rect 4233 29652 4260 29708
rect 4316 29652 4321 29708
rect 3121 29614 4321 29652
rect 3121 29558 3513 29614
rect 3569 29558 3596 29614
rect 3652 29558 3679 29614
rect 3735 29558 3762 29614
rect 3818 29558 3845 29614
rect 3901 29558 3928 29614
rect 3984 29558 4011 29614
rect 4067 29558 4094 29614
rect 4150 29558 4177 29614
rect 4233 29558 4260 29614
rect 4316 29558 4321 29614
rect 3121 29520 4321 29558
rect 3121 29464 3513 29520
rect 3569 29464 3596 29520
rect 3652 29464 3679 29520
rect 3735 29464 3762 29520
rect 3818 29464 3845 29520
rect 3901 29464 3928 29520
rect 3984 29464 4011 29520
rect 4067 29464 4094 29520
rect 4150 29464 4177 29520
rect 4233 29464 4260 29520
rect 4316 29464 4321 29520
rect 3121 29426 4321 29464
rect 3121 29370 3513 29426
rect 3569 29370 3596 29426
rect 3652 29370 3679 29426
rect 3735 29370 3762 29426
rect 3818 29370 3845 29426
rect 3901 29370 3928 29426
rect 3984 29370 4011 29426
rect 4067 29370 4094 29426
rect 4150 29370 4177 29426
rect 4233 29370 4260 29426
rect 4316 29370 4321 29426
rect 3121 27896 4321 29370
rect 3121 27840 3452 27896
rect 3508 27840 3532 27896
rect 3588 27840 3612 27896
rect 3668 27840 3693 27896
rect 3749 27840 3774 27896
rect 3830 27840 3855 27896
rect 3911 27840 3936 27896
rect 3992 27840 4017 27896
rect 4073 27840 4098 27896
rect 4154 27840 4179 27896
rect 4235 27840 4260 27896
rect 4316 27840 4321 27896
rect 3121 27802 4321 27840
rect 3121 27746 3452 27802
rect 3508 27746 3532 27802
rect 3588 27746 3612 27802
rect 3668 27746 3693 27802
rect 3749 27746 3774 27802
rect 3830 27746 3855 27802
rect 3911 27746 3936 27802
rect 3992 27746 4017 27802
rect 4073 27746 4098 27802
rect 4154 27746 4179 27802
rect 4235 27746 4260 27802
rect 4316 27746 4321 27802
rect 3121 27708 4321 27746
rect 3121 27652 3452 27708
rect 3508 27652 3532 27708
rect 3588 27652 3612 27708
rect 3668 27652 3693 27708
rect 3749 27652 3774 27708
rect 3830 27652 3855 27708
rect 3911 27652 3936 27708
rect 3992 27652 4017 27708
rect 4073 27652 4098 27708
rect 4154 27652 4179 27708
rect 4235 27652 4260 27708
rect 4316 27652 4321 27708
rect 3121 27614 4321 27652
rect 3121 27558 3452 27614
rect 3508 27558 3532 27614
rect 3588 27558 3612 27614
rect 3668 27558 3693 27614
rect 3749 27558 3774 27614
rect 3830 27558 3855 27614
rect 3911 27558 3936 27614
rect 3992 27558 4017 27614
rect 4073 27558 4098 27614
rect 4154 27558 4179 27614
rect 4235 27558 4260 27614
rect 4316 27558 4321 27614
rect 3121 27520 4321 27558
rect 3121 27464 3452 27520
rect 3508 27464 3532 27520
rect 3588 27464 3612 27520
rect 3668 27464 3693 27520
rect 3749 27464 3774 27520
rect 3830 27464 3855 27520
rect 3911 27464 3936 27520
rect 3992 27464 4017 27520
rect 4073 27464 4098 27520
rect 4154 27464 4179 27520
rect 4235 27464 4260 27520
rect 4316 27464 4321 27520
rect 3121 27426 4321 27464
rect 3121 27370 3452 27426
rect 3508 27370 3532 27426
rect 3588 27370 3612 27426
rect 3668 27370 3693 27426
rect 3749 27370 3774 27426
rect 3830 27370 3855 27426
rect 3911 27370 3936 27426
rect 3992 27370 4017 27426
rect 4073 27370 4098 27426
rect 4154 27370 4179 27426
rect 4235 27370 4260 27426
rect 4316 27370 4321 27426
rect 3121 25882 4321 27370
rect 3121 25826 3443 25882
rect 3499 25826 3525 25882
rect 3581 25826 3607 25882
rect 3663 25826 3689 25882
rect 3745 25826 3771 25882
rect 3827 25826 3853 25882
rect 3909 25826 3935 25882
rect 3991 25826 4017 25882
rect 4073 25826 4098 25882
rect 4154 25826 4179 25882
rect 4235 25826 4260 25882
rect 4316 25826 4321 25882
rect 3121 25794 4321 25826
rect 3121 25738 3443 25794
rect 3499 25738 3525 25794
rect 3581 25738 3607 25794
rect 3663 25738 3689 25794
rect 3745 25738 3771 25794
rect 3827 25738 3853 25794
rect 3909 25738 3935 25794
rect 3991 25738 4017 25794
rect 4073 25738 4098 25794
rect 4154 25738 4179 25794
rect 4235 25738 4260 25794
rect 4316 25738 4321 25794
rect 3121 25706 4321 25738
rect 3121 25650 3443 25706
rect 3499 25650 3525 25706
rect 3581 25650 3607 25706
rect 3663 25650 3689 25706
rect 3745 25650 3771 25706
rect 3827 25650 3853 25706
rect 3909 25650 3935 25706
rect 3991 25650 4017 25706
rect 4073 25650 4098 25706
rect 4154 25650 4179 25706
rect 4235 25650 4260 25706
rect 4316 25650 4321 25706
rect 3121 25618 4321 25650
rect 3121 25562 3443 25618
rect 3499 25562 3525 25618
rect 3581 25562 3607 25618
rect 3663 25562 3689 25618
rect 3745 25562 3771 25618
rect 3827 25562 3853 25618
rect 3909 25562 3935 25618
rect 3991 25562 4017 25618
rect 4073 25562 4098 25618
rect 4154 25562 4179 25618
rect 4235 25562 4260 25618
rect 4316 25562 4321 25618
rect 3121 25530 4321 25562
rect 3121 25474 3443 25530
rect 3499 25474 3525 25530
rect 3581 25474 3607 25530
rect 3663 25474 3689 25530
rect 3745 25474 3771 25530
rect 3827 25474 3853 25530
rect 3909 25474 3935 25530
rect 3991 25474 4017 25530
rect 4073 25474 4098 25530
rect 4154 25474 4179 25530
rect 4235 25474 4260 25530
rect 4316 25474 4321 25530
rect 3121 25442 4321 25474
rect 3121 25386 3443 25442
rect 3499 25386 3525 25442
rect 3581 25386 3607 25442
rect 3663 25386 3689 25442
rect 3745 25386 3771 25442
rect 3827 25386 3853 25442
rect 3909 25386 3935 25442
rect 3991 25386 4017 25442
rect 4073 25386 4098 25442
rect 4154 25386 4179 25442
rect 4235 25386 4260 25442
rect 4316 25386 4321 25442
rect 3121 19083 4321 25386
rect 5207 33382 5216 33438
rect 5272 33382 5299 33438
rect 5355 33382 5382 33438
rect 5438 33382 5465 33438
rect 5521 33382 5548 33438
rect 5604 33382 5631 33438
rect 5687 33382 5714 33438
rect 5770 33382 5797 33438
rect 5853 33382 5880 33438
rect 5936 33382 5963 33438
rect 6019 33382 6046 33438
rect 6102 33382 6129 33438
rect 6185 33382 6211 33438
rect 6267 33382 6293 33438
rect 6349 33382 6375 33438
rect 6431 33382 6457 33438
rect 6513 33382 6539 33438
rect 6595 33382 6621 33438
rect 6677 33382 6703 33438
rect 6759 33382 6785 33438
rect 6841 33382 6867 33438
rect 6923 33382 6949 33438
rect 7005 33382 7031 33438
rect 7087 33382 7113 33438
rect 7169 33382 7195 33438
rect 7251 33382 7275 33438
tri 7275 33382 7331 33438 nw
tri 7956 33382 8012 33438 ne
rect 8012 33382 8041 33438
rect 8097 33382 8124 33438
rect 8180 33382 8207 33438
rect 8263 33382 8290 33438
rect 8346 33382 8373 33438
rect 8429 33382 8456 33438
rect 8512 33382 8539 33438
rect 8595 33382 8622 33438
rect 8678 33382 8705 33438
rect 8761 33382 8788 33438
rect 8844 33382 8871 33438
rect 8927 33382 8954 33438
rect 9010 33382 9037 33438
rect 9093 33382 9120 33438
rect 9176 33382 9203 33438
rect 9259 33382 9286 33438
rect 9342 33382 9369 33438
rect 9425 33382 9452 33438
rect 9508 33382 9535 33438
rect 9591 33382 9618 33438
rect 9674 33382 9702 33438
rect 9758 33382 9767 33438
tri 10320 33382 10376 33438 ne
rect 10376 33382 10397 33438
rect 10453 33382 10477 33438
rect 10533 33382 10557 33438
rect 10613 33382 10637 33438
rect 10693 33382 10717 33438
rect 10773 33382 10797 33438
rect 10853 33382 10877 33438
rect 10933 33382 10957 33438
rect 11013 33382 11037 33438
rect 11093 33382 11117 33438
rect 11173 33382 11197 33438
rect 11253 33382 11277 33438
rect 11333 33382 11357 33438
rect 11413 33382 11437 33438
rect 11493 33382 11517 33438
rect 11573 33382 11597 33438
rect 11653 33382 11677 33438
rect 11733 33382 11758 33438
rect 11814 33382 11839 33438
rect 11895 33382 11920 33438
rect 11976 33382 12001 33438
rect 12057 33382 12066 33438
rect 5207 33373 7266 33382
tri 7266 33373 7275 33382 nw
tri 8012 33373 8021 33382 ne
rect 8021 33373 9767 33382
tri 10376 33373 10385 33382 ne
rect 10385 33373 12066 33382
rect 5207 32875 6768 33373
tri 6768 32875 7266 33373 nw
tri 8021 32892 8502 33373 ne
rect 8502 32892 9767 33373
tri 10385 32892 10866 33373 ne
tri 8502 32875 8519 32892 ne
rect 8519 32875 9767 32892
rect 5207 31883 6407 32875
tri 6407 32514 6768 32875 nw
tri 8519 32827 8567 32875 ne
rect 5207 31827 5215 31883
rect 5271 31827 5296 31883
rect 5352 31827 5377 31883
rect 5433 31827 5458 31883
rect 5514 31827 5539 31883
rect 5595 31827 5620 31883
rect 5676 31827 5701 31883
rect 5757 31827 5782 31883
rect 5838 31827 5863 31883
rect 5919 31827 5944 31883
rect 6000 31827 6025 31883
rect 6081 31827 6106 31883
rect 6162 31827 6186 31883
rect 6242 31827 6266 31883
rect 6322 31827 6346 31883
rect 6402 31827 6407 31883
rect 5207 31795 6407 31827
rect 5207 31739 5215 31795
rect 5271 31739 5296 31795
rect 5352 31739 5377 31795
rect 5433 31739 5458 31795
rect 5514 31739 5539 31795
rect 5595 31739 5620 31795
rect 5676 31739 5701 31795
rect 5757 31739 5782 31795
rect 5838 31739 5863 31795
rect 5919 31739 5944 31795
rect 6000 31739 6025 31795
rect 6081 31739 6106 31795
rect 6162 31739 6186 31795
rect 6242 31739 6266 31795
rect 6322 31739 6346 31795
rect 6402 31739 6407 31795
rect 5207 31707 6407 31739
rect 5207 31651 5215 31707
rect 5271 31651 5296 31707
rect 5352 31651 5377 31707
rect 5433 31651 5458 31707
rect 5514 31651 5539 31707
rect 5595 31651 5620 31707
rect 5676 31651 5701 31707
rect 5757 31651 5782 31707
rect 5838 31651 5863 31707
rect 5919 31651 5944 31707
rect 6000 31651 6025 31707
rect 6081 31651 6106 31707
rect 6162 31651 6186 31707
rect 6242 31651 6266 31707
rect 6322 31651 6346 31707
rect 6402 31651 6407 31707
rect 5207 31619 6407 31651
rect 5207 31563 5215 31619
rect 5271 31563 5296 31619
rect 5352 31563 5377 31619
rect 5433 31563 5458 31619
rect 5514 31563 5539 31619
rect 5595 31563 5620 31619
rect 5676 31563 5701 31619
rect 5757 31563 5782 31619
rect 5838 31563 5863 31619
rect 5919 31563 5944 31619
rect 6000 31563 6025 31619
rect 6081 31563 6106 31619
rect 6162 31563 6186 31619
rect 6242 31563 6266 31619
rect 6322 31563 6346 31619
rect 6402 31563 6407 31619
rect 5207 31531 6407 31563
rect 5207 31475 5215 31531
rect 5271 31475 5296 31531
rect 5352 31475 5377 31531
rect 5433 31475 5458 31531
rect 5514 31475 5539 31531
rect 5595 31475 5620 31531
rect 5676 31475 5701 31531
rect 5757 31475 5782 31531
rect 5838 31475 5863 31531
rect 5919 31475 5944 31531
rect 6000 31475 6025 31531
rect 6081 31475 6106 31531
rect 6162 31475 6186 31531
rect 6242 31475 6266 31531
rect 6322 31475 6346 31531
rect 6402 31475 6407 31531
rect 5207 31443 6407 31475
rect 5207 31387 5215 31443
rect 5271 31387 5296 31443
rect 5352 31387 5377 31443
rect 5433 31387 5458 31443
rect 5514 31387 5539 31443
rect 5595 31387 5620 31443
rect 5676 31387 5701 31443
rect 5757 31387 5782 31443
rect 5838 31387 5863 31443
rect 5919 31387 5944 31443
rect 6000 31387 6025 31443
rect 6081 31387 6106 31443
rect 6162 31387 6186 31443
rect 6242 31387 6266 31443
rect 6322 31387 6346 31443
rect 6402 31387 6407 31443
rect 5207 29883 6407 31387
rect 5207 29827 5215 29883
rect 5271 29827 5296 29883
rect 5352 29827 5377 29883
rect 5433 29827 5458 29883
rect 5514 29827 5539 29883
rect 5595 29827 5620 29883
rect 5676 29827 5701 29883
rect 5757 29827 5782 29883
rect 5838 29827 5863 29883
rect 5919 29827 5944 29883
rect 6000 29827 6025 29883
rect 6081 29827 6106 29883
rect 6162 29827 6186 29883
rect 6242 29827 6266 29883
rect 6322 29827 6346 29883
rect 6402 29827 6407 29883
rect 5207 29795 6407 29827
rect 5207 29739 5215 29795
rect 5271 29739 5296 29795
rect 5352 29739 5377 29795
rect 5433 29739 5458 29795
rect 5514 29739 5539 29795
rect 5595 29739 5620 29795
rect 5676 29739 5701 29795
rect 5757 29739 5782 29795
rect 5838 29739 5863 29795
rect 5919 29739 5944 29795
rect 6000 29739 6025 29795
rect 6081 29739 6106 29795
rect 6162 29739 6186 29795
rect 6242 29739 6266 29795
rect 6322 29739 6346 29795
rect 6402 29739 6407 29795
rect 5207 29707 6407 29739
rect 5207 29651 5215 29707
rect 5271 29651 5296 29707
rect 5352 29651 5377 29707
rect 5433 29651 5458 29707
rect 5514 29651 5539 29707
rect 5595 29651 5620 29707
rect 5676 29651 5701 29707
rect 5757 29651 5782 29707
rect 5838 29651 5863 29707
rect 5919 29651 5944 29707
rect 6000 29651 6025 29707
rect 6081 29651 6106 29707
rect 6162 29651 6186 29707
rect 6242 29651 6266 29707
rect 6322 29651 6346 29707
rect 6402 29651 6407 29707
rect 5207 29619 6407 29651
rect 5207 29563 5215 29619
rect 5271 29563 5296 29619
rect 5352 29563 5377 29619
rect 5433 29563 5458 29619
rect 5514 29563 5539 29619
rect 5595 29563 5620 29619
rect 5676 29563 5701 29619
rect 5757 29563 5782 29619
rect 5838 29563 5863 29619
rect 5919 29563 5944 29619
rect 6000 29563 6025 29619
rect 6081 29563 6106 29619
rect 6162 29563 6186 29619
rect 6242 29563 6266 29619
rect 6322 29563 6346 29619
rect 6402 29563 6407 29619
rect 5207 29531 6407 29563
rect 5207 29475 5215 29531
rect 5271 29475 5296 29531
rect 5352 29475 5377 29531
rect 5433 29475 5458 29531
rect 5514 29475 5539 29531
rect 5595 29475 5620 29531
rect 5676 29475 5701 29531
rect 5757 29475 5782 29531
rect 5838 29475 5863 29531
rect 5919 29475 5944 29531
rect 6000 29475 6025 29531
rect 6081 29475 6106 29531
rect 6162 29475 6186 29531
rect 6242 29475 6266 29531
rect 6322 29475 6346 29531
rect 6402 29475 6407 29531
rect 5207 29443 6407 29475
rect 5207 29387 5215 29443
rect 5271 29387 5296 29443
rect 5352 29387 5377 29443
rect 5433 29387 5458 29443
rect 5514 29387 5539 29443
rect 5595 29387 5620 29443
rect 5676 29387 5701 29443
rect 5757 29387 5782 29443
rect 5838 29387 5863 29443
rect 5919 29387 5944 29443
rect 6000 29387 6025 29443
rect 6081 29387 6106 29443
rect 6162 29387 6186 29443
rect 6242 29387 6266 29443
rect 6322 29387 6346 29443
rect 6402 29387 6407 29443
rect 5207 27883 6407 29387
rect 5207 27827 5215 27883
rect 5271 27827 5296 27883
rect 5352 27827 5377 27883
rect 5433 27827 5458 27883
rect 5514 27827 5539 27883
rect 5595 27827 5620 27883
rect 5676 27827 5701 27883
rect 5757 27827 5782 27883
rect 5838 27827 5863 27883
rect 5919 27827 5944 27883
rect 6000 27827 6025 27883
rect 6081 27827 6106 27883
rect 6162 27827 6186 27883
rect 6242 27827 6266 27883
rect 6322 27827 6346 27883
rect 6402 27827 6407 27883
rect 5207 27795 6407 27827
rect 5207 27739 5215 27795
rect 5271 27739 5296 27795
rect 5352 27739 5377 27795
rect 5433 27739 5458 27795
rect 5514 27739 5539 27795
rect 5595 27739 5620 27795
rect 5676 27739 5701 27795
rect 5757 27739 5782 27795
rect 5838 27739 5863 27795
rect 5919 27739 5944 27795
rect 6000 27739 6025 27795
rect 6081 27739 6106 27795
rect 6162 27739 6186 27795
rect 6242 27739 6266 27795
rect 6322 27739 6346 27795
rect 6402 27739 6407 27795
rect 5207 27707 6407 27739
rect 5207 27651 5215 27707
rect 5271 27651 5296 27707
rect 5352 27651 5377 27707
rect 5433 27651 5458 27707
rect 5514 27651 5539 27707
rect 5595 27651 5620 27707
rect 5676 27651 5701 27707
rect 5757 27651 5782 27707
rect 5838 27651 5863 27707
rect 5919 27651 5944 27707
rect 6000 27651 6025 27707
rect 6081 27651 6106 27707
rect 6162 27651 6186 27707
rect 6242 27651 6266 27707
rect 6322 27651 6346 27707
rect 6402 27651 6407 27707
rect 5207 27619 6407 27651
rect 5207 27563 5215 27619
rect 5271 27563 5296 27619
rect 5352 27563 5377 27619
rect 5433 27563 5458 27619
rect 5514 27563 5539 27619
rect 5595 27563 5620 27619
rect 5676 27563 5701 27619
rect 5757 27563 5782 27619
rect 5838 27563 5863 27619
rect 5919 27563 5944 27619
rect 6000 27563 6025 27619
rect 6081 27563 6106 27619
rect 6162 27563 6186 27619
rect 6242 27563 6266 27619
rect 6322 27563 6346 27619
rect 6402 27563 6407 27619
rect 5207 27531 6407 27563
rect 5207 27475 5215 27531
rect 5271 27475 5296 27531
rect 5352 27475 5377 27531
rect 5433 27475 5458 27531
rect 5514 27475 5539 27531
rect 5595 27475 5620 27531
rect 5676 27475 5701 27531
rect 5757 27475 5782 27531
rect 5838 27475 5863 27531
rect 5919 27475 5944 27531
rect 6000 27475 6025 27531
rect 6081 27475 6106 27531
rect 6162 27475 6186 27531
rect 6242 27475 6266 27531
rect 6322 27475 6346 27531
rect 6402 27475 6407 27531
rect 5207 27443 6407 27475
rect 5207 27387 5215 27443
rect 5271 27387 5296 27443
rect 5352 27387 5377 27443
rect 5433 27387 5458 27443
rect 5514 27387 5539 27443
rect 5595 27387 5620 27443
rect 5676 27387 5701 27443
rect 5757 27387 5782 27443
rect 5838 27387 5863 27443
rect 5919 27387 5944 27443
rect 6000 27387 6025 27443
rect 6081 27387 6106 27443
rect 6162 27387 6186 27443
rect 6242 27387 6266 27443
rect 6322 27387 6346 27443
rect 6402 27387 6407 27443
rect 5207 25882 6407 27387
rect 5207 25826 5215 25882
rect 5271 25826 5296 25882
rect 5352 25826 5377 25882
rect 5433 25826 5458 25882
rect 5514 25826 5539 25882
rect 5595 25826 5620 25882
rect 5676 25826 5701 25882
rect 5757 25826 5782 25882
rect 5838 25826 5863 25882
rect 5919 25826 5944 25882
rect 6000 25826 6025 25882
rect 6081 25826 6106 25882
rect 6162 25826 6186 25882
rect 6242 25826 6266 25882
rect 6322 25826 6346 25882
rect 6402 25826 6407 25882
rect 5207 25794 6407 25826
rect 5207 25738 5215 25794
rect 5271 25738 5296 25794
rect 5352 25738 5377 25794
rect 5433 25738 5458 25794
rect 5514 25738 5539 25794
rect 5595 25738 5620 25794
rect 5676 25738 5701 25794
rect 5757 25738 5782 25794
rect 5838 25738 5863 25794
rect 5919 25738 5944 25794
rect 6000 25738 6025 25794
rect 6081 25738 6106 25794
rect 6162 25738 6186 25794
rect 6242 25738 6266 25794
rect 6322 25738 6346 25794
rect 6402 25738 6407 25794
rect 5207 25706 6407 25738
rect 5207 25650 5215 25706
rect 5271 25650 5296 25706
rect 5352 25650 5377 25706
rect 5433 25650 5458 25706
rect 5514 25650 5539 25706
rect 5595 25650 5620 25706
rect 5676 25650 5701 25706
rect 5757 25650 5782 25706
rect 5838 25650 5863 25706
rect 5919 25650 5944 25706
rect 6000 25650 6025 25706
rect 6081 25650 6106 25706
rect 6162 25650 6186 25706
rect 6242 25650 6266 25706
rect 6322 25650 6346 25706
rect 6402 25650 6407 25706
rect 5207 25618 6407 25650
rect 5207 25562 5215 25618
rect 5271 25562 5296 25618
rect 5352 25562 5377 25618
rect 5433 25562 5458 25618
rect 5514 25562 5539 25618
rect 5595 25562 5620 25618
rect 5676 25562 5701 25618
rect 5757 25562 5782 25618
rect 5838 25562 5863 25618
rect 5919 25562 5944 25618
rect 6000 25562 6025 25618
rect 6081 25562 6106 25618
rect 6162 25562 6186 25618
rect 6242 25562 6266 25618
rect 6322 25562 6346 25618
rect 6402 25562 6407 25618
rect 5207 25530 6407 25562
rect 5207 25474 5215 25530
rect 5271 25474 5296 25530
rect 5352 25474 5377 25530
rect 5433 25474 5458 25530
rect 5514 25474 5539 25530
rect 5595 25474 5620 25530
rect 5676 25474 5701 25530
rect 5757 25474 5782 25530
rect 5838 25474 5863 25530
rect 5919 25474 5944 25530
rect 6000 25474 6025 25530
rect 6081 25474 6106 25530
rect 6162 25474 6186 25530
rect 6242 25474 6266 25530
rect 6322 25474 6346 25530
rect 6402 25474 6407 25530
rect 5207 25442 6407 25474
rect 5207 25386 5215 25442
rect 5271 25386 5296 25442
rect 5352 25386 5377 25442
rect 5433 25386 5458 25442
rect 5514 25386 5539 25442
rect 5595 25386 5620 25442
rect 5676 25386 5701 25442
rect 5757 25386 5782 25442
rect 5838 25386 5863 25442
rect 5919 25386 5944 25442
rect 6000 25386 6025 25442
rect 6081 25386 6106 25442
rect 6162 25386 6186 25442
rect 6242 25386 6266 25442
rect 6322 25386 6346 25442
rect 6402 25386 6407 25442
tri 4321 19083 4596 19358 sw
rect 3121 18900 4596 19083
tri 4596 18900 4779 19083 sw
rect 5207 18900 6407 25386
rect 8567 31883 9767 32875
rect 8567 31827 8572 31883
rect 8628 31827 8652 31883
rect 8708 31827 8732 31883
rect 8788 31827 8812 31883
rect 8868 31827 8893 31883
rect 8949 31827 8974 31883
rect 9030 31827 9055 31883
rect 9111 31827 9136 31883
rect 9192 31827 9217 31883
rect 9273 31827 9298 31883
rect 9354 31827 9379 31883
rect 9435 31827 9460 31883
rect 9516 31827 9541 31883
rect 9597 31827 9622 31883
rect 9678 31827 9703 31883
rect 9759 31827 9767 31883
rect 8567 31795 9767 31827
rect 8567 31739 8572 31795
rect 8628 31739 8652 31795
rect 8708 31739 8732 31795
rect 8788 31739 8812 31795
rect 8868 31739 8893 31795
rect 8949 31739 8974 31795
rect 9030 31739 9055 31795
rect 9111 31739 9136 31795
rect 9192 31739 9217 31795
rect 9273 31739 9298 31795
rect 9354 31739 9379 31795
rect 9435 31739 9460 31795
rect 9516 31739 9541 31795
rect 9597 31739 9622 31795
rect 9678 31739 9703 31795
rect 9759 31739 9767 31795
rect 8567 31707 9767 31739
rect 8567 31651 8572 31707
rect 8628 31651 8652 31707
rect 8708 31651 8732 31707
rect 8788 31651 8812 31707
rect 8868 31651 8893 31707
rect 8949 31651 8974 31707
rect 9030 31651 9055 31707
rect 9111 31651 9136 31707
rect 9192 31651 9217 31707
rect 9273 31651 9298 31707
rect 9354 31651 9379 31707
rect 9435 31651 9460 31707
rect 9516 31651 9541 31707
rect 9597 31651 9622 31707
rect 9678 31651 9703 31707
rect 9759 31651 9767 31707
rect 8567 31619 9767 31651
rect 8567 31563 8572 31619
rect 8628 31563 8652 31619
rect 8708 31563 8732 31619
rect 8788 31563 8812 31619
rect 8868 31563 8893 31619
rect 8949 31563 8974 31619
rect 9030 31563 9055 31619
rect 9111 31563 9136 31619
rect 9192 31563 9217 31619
rect 9273 31563 9298 31619
rect 9354 31563 9379 31619
rect 9435 31563 9460 31619
rect 9516 31563 9541 31619
rect 9597 31563 9622 31619
rect 9678 31563 9703 31619
rect 9759 31563 9767 31619
rect 8567 31531 9767 31563
rect 8567 31475 8572 31531
rect 8628 31475 8652 31531
rect 8708 31475 8732 31531
rect 8788 31475 8812 31531
rect 8868 31475 8893 31531
rect 8949 31475 8974 31531
rect 9030 31475 9055 31531
rect 9111 31475 9136 31531
rect 9192 31475 9217 31531
rect 9273 31475 9298 31531
rect 9354 31475 9379 31531
rect 9435 31475 9460 31531
rect 9516 31475 9541 31531
rect 9597 31475 9622 31531
rect 9678 31475 9703 31531
rect 9759 31475 9767 31531
rect 8567 31443 9767 31475
rect 8567 31387 8572 31443
rect 8628 31387 8652 31443
rect 8708 31387 8732 31443
rect 8788 31387 8812 31443
rect 8868 31387 8893 31443
rect 8949 31387 8974 31443
rect 9030 31387 9055 31443
rect 9111 31387 9136 31443
rect 9192 31387 9217 31443
rect 9273 31387 9298 31443
rect 9354 31387 9379 31443
rect 9435 31387 9460 31443
rect 9516 31387 9541 31443
rect 9597 31387 9622 31443
rect 9678 31387 9703 31443
rect 9759 31387 9767 31443
rect 8567 29883 9767 31387
rect 8567 29827 8572 29883
rect 8628 29827 8652 29883
rect 8708 29827 8732 29883
rect 8788 29827 8812 29883
rect 8868 29827 8893 29883
rect 8949 29827 8974 29883
rect 9030 29827 9055 29883
rect 9111 29827 9136 29883
rect 9192 29827 9217 29883
rect 9273 29827 9298 29883
rect 9354 29827 9379 29883
rect 9435 29827 9460 29883
rect 9516 29827 9541 29883
rect 9597 29827 9622 29883
rect 9678 29827 9703 29883
rect 9759 29827 9767 29883
rect 8567 29795 9767 29827
rect 8567 29739 8572 29795
rect 8628 29739 8652 29795
rect 8708 29739 8732 29795
rect 8788 29739 8812 29795
rect 8868 29739 8893 29795
rect 8949 29739 8974 29795
rect 9030 29739 9055 29795
rect 9111 29739 9136 29795
rect 9192 29739 9217 29795
rect 9273 29739 9298 29795
rect 9354 29739 9379 29795
rect 9435 29739 9460 29795
rect 9516 29739 9541 29795
rect 9597 29739 9622 29795
rect 9678 29739 9703 29795
rect 9759 29739 9767 29795
rect 8567 29707 9767 29739
rect 8567 29651 8572 29707
rect 8628 29651 8652 29707
rect 8708 29651 8732 29707
rect 8788 29651 8812 29707
rect 8868 29651 8893 29707
rect 8949 29651 8974 29707
rect 9030 29651 9055 29707
rect 9111 29651 9136 29707
rect 9192 29651 9217 29707
rect 9273 29651 9298 29707
rect 9354 29651 9379 29707
rect 9435 29651 9460 29707
rect 9516 29651 9541 29707
rect 9597 29651 9622 29707
rect 9678 29651 9703 29707
rect 9759 29651 9767 29707
rect 8567 29619 9767 29651
rect 8567 29563 8572 29619
rect 8628 29563 8652 29619
rect 8708 29563 8732 29619
rect 8788 29563 8812 29619
rect 8868 29563 8893 29619
rect 8949 29563 8974 29619
rect 9030 29563 9055 29619
rect 9111 29563 9136 29619
rect 9192 29563 9217 29619
rect 9273 29563 9298 29619
rect 9354 29563 9379 29619
rect 9435 29563 9460 29619
rect 9516 29563 9541 29619
rect 9597 29563 9622 29619
rect 9678 29563 9703 29619
rect 9759 29563 9767 29619
rect 8567 29531 9767 29563
rect 8567 29475 8572 29531
rect 8628 29475 8652 29531
rect 8708 29475 8732 29531
rect 8788 29475 8812 29531
rect 8868 29475 8893 29531
rect 8949 29475 8974 29531
rect 9030 29475 9055 29531
rect 9111 29475 9136 29531
rect 9192 29475 9217 29531
rect 9273 29475 9298 29531
rect 9354 29475 9379 29531
rect 9435 29475 9460 29531
rect 9516 29475 9541 29531
rect 9597 29475 9622 29531
rect 9678 29475 9703 29531
rect 9759 29475 9767 29531
rect 8567 29443 9767 29475
rect 8567 29387 8572 29443
rect 8628 29387 8652 29443
rect 8708 29387 8732 29443
rect 8788 29387 8812 29443
rect 8868 29387 8893 29443
rect 8949 29387 8974 29443
rect 9030 29387 9055 29443
rect 9111 29387 9136 29443
rect 9192 29387 9217 29443
rect 9273 29387 9298 29443
rect 9354 29387 9379 29443
rect 9435 29387 9460 29443
rect 9516 29387 9541 29443
rect 9597 29387 9622 29443
rect 9678 29387 9703 29443
rect 9759 29387 9767 29443
rect 8567 27883 9767 29387
rect 8567 27827 8572 27883
rect 8628 27827 8652 27883
rect 8708 27827 8732 27883
rect 8788 27827 8812 27883
rect 8868 27827 8893 27883
rect 8949 27827 8974 27883
rect 9030 27827 9055 27883
rect 9111 27827 9136 27883
rect 9192 27827 9217 27883
rect 9273 27827 9298 27883
rect 9354 27827 9379 27883
rect 9435 27827 9460 27883
rect 9516 27827 9541 27883
rect 9597 27827 9622 27883
rect 9678 27827 9703 27883
rect 9759 27827 9767 27883
rect 8567 27795 9767 27827
rect 8567 27739 8572 27795
rect 8628 27739 8652 27795
rect 8708 27739 8732 27795
rect 8788 27739 8812 27795
rect 8868 27739 8893 27795
rect 8949 27739 8974 27795
rect 9030 27739 9055 27795
rect 9111 27739 9136 27795
rect 9192 27739 9217 27795
rect 9273 27739 9298 27795
rect 9354 27739 9379 27795
rect 9435 27739 9460 27795
rect 9516 27739 9541 27795
rect 9597 27739 9622 27795
rect 9678 27739 9703 27795
rect 9759 27739 9767 27795
rect 8567 27707 9767 27739
rect 8567 27651 8572 27707
rect 8628 27651 8652 27707
rect 8708 27651 8732 27707
rect 8788 27651 8812 27707
rect 8868 27651 8893 27707
rect 8949 27651 8974 27707
rect 9030 27651 9055 27707
rect 9111 27651 9136 27707
rect 9192 27651 9217 27707
rect 9273 27651 9298 27707
rect 9354 27651 9379 27707
rect 9435 27651 9460 27707
rect 9516 27651 9541 27707
rect 9597 27651 9622 27707
rect 9678 27651 9703 27707
rect 9759 27651 9767 27707
rect 8567 27619 9767 27651
rect 8567 27563 8572 27619
rect 8628 27563 8652 27619
rect 8708 27563 8732 27619
rect 8788 27563 8812 27619
rect 8868 27563 8893 27619
rect 8949 27563 8974 27619
rect 9030 27563 9055 27619
rect 9111 27563 9136 27619
rect 9192 27563 9217 27619
rect 9273 27563 9298 27619
rect 9354 27563 9379 27619
rect 9435 27563 9460 27619
rect 9516 27563 9541 27619
rect 9597 27563 9622 27619
rect 9678 27563 9703 27619
rect 9759 27563 9767 27619
rect 8567 27531 9767 27563
rect 8567 27475 8572 27531
rect 8628 27475 8652 27531
rect 8708 27475 8732 27531
rect 8788 27475 8812 27531
rect 8868 27475 8893 27531
rect 8949 27475 8974 27531
rect 9030 27475 9055 27531
rect 9111 27475 9136 27531
rect 9192 27475 9217 27531
rect 9273 27475 9298 27531
rect 9354 27475 9379 27531
rect 9435 27475 9460 27531
rect 9516 27475 9541 27531
rect 9597 27475 9622 27531
rect 9678 27475 9703 27531
rect 9759 27475 9767 27531
rect 8567 27443 9767 27475
rect 8567 27387 8572 27443
rect 8628 27387 8652 27443
rect 8708 27387 8732 27443
rect 8788 27387 8812 27443
rect 8868 27387 8893 27443
rect 8949 27387 8974 27443
rect 9030 27387 9055 27443
rect 9111 27387 9136 27443
rect 9192 27387 9217 27443
rect 9273 27387 9298 27443
rect 9354 27387 9379 27443
rect 9435 27387 9460 27443
rect 9516 27387 9541 27443
rect 9597 27387 9622 27443
rect 9678 27387 9703 27443
rect 9759 27387 9767 27443
rect 8567 25882 9767 27387
rect 8567 25826 8572 25882
rect 8628 25826 8652 25882
rect 8708 25826 8732 25882
rect 8788 25826 8812 25882
rect 8868 25826 8893 25882
rect 8949 25826 8974 25882
rect 9030 25826 9055 25882
rect 9111 25826 9136 25882
rect 9192 25826 9217 25882
rect 9273 25826 9298 25882
rect 9354 25826 9379 25882
rect 9435 25826 9460 25882
rect 9516 25826 9541 25882
rect 9597 25826 9622 25882
rect 9678 25826 9703 25882
rect 9759 25826 9767 25882
rect 8567 25794 9767 25826
rect 8567 25738 8572 25794
rect 8628 25738 8652 25794
rect 8708 25738 8732 25794
rect 8788 25738 8812 25794
rect 8868 25738 8893 25794
rect 8949 25738 8974 25794
rect 9030 25738 9055 25794
rect 9111 25738 9136 25794
rect 9192 25738 9217 25794
rect 9273 25738 9298 25794
rect 9354 25738 9379 25794
rect 9435 25738 9460 25794
rect 9516 25738 9541 25794
rect 9597 25738 9622 25794
rect 9678 25738 9703 25794
rect 9759 25738 9767 25794
rect 8567 25706 9767 25738
rect 8567 25650 8572 25706
rect 8628 25650 8652 25706
rect 8708 25650 8732 25706
rect 8788 25650 8812 25706
rect 8868 25650 8893 25706
rect 8949 25650 8974 25706
rect 9030 25650 9055 25706
rect 9111 25650 9136 25706
rect 9192 25650 9217 25706
rect 9273 25650 9298 25706
rect 9354 25650 9379 25706
rect 9435 25650 9460 25706
rect 9516 25650 9541 25706
rect 9597 25650 9622 25706
rect 9678 25650 9703 25706
rect 9759 25650 9767 25706
rect 8567 25618 9767 25650
rect 8567 25562 8572 25618
rect 8628 25562 8652 25618
rect 8708 25562 8732 25618
rect 8788 25562 8812 25618
rect 8868 25562 8893 25618
rect 8949 25562 8974 25618
rect 9030 25562 9055 25618
rect 9111 25562 9136 25618
rect 9192 25562 9217 25618
rect 9273 25562 9298 25618
rect 9354 25562 9379 25618
rect 9435 25562 9460 25618
rect 9516 25562 9541 25618
rect 9597 25562 9622 25618
rect 9678 25562 9703 25618
rect 9759 25562 9767 25618
rect 8567 25530 9767 25562
rect 8567 25474 8572 25530
rect 8628 25474 8652 25530
rect 8708 25474 8732 25530
rect 8788 25474 8812 25530
rect 8868 25474 8893 25530
rect 8949 25474 8974 25530
rect 9030 25474 9055 25530
rect 9111 25474 9136 25530
rect 9192 25474 9217 25530
rect 9273 25474 9298 25530
rect 9354 25474 9379 25530
rect 9435 25474 9460 25530
rect 9516 25474 9541 25530
rect 9597 25474 9622 25530
rect 9678 25474 9703 25530
rect 9759 25474 9767 25530
rect 8567 25442 9767 25474
rect 8567 25386 8572 25442
rect 8628 25386 8652 25442
rect 8708 25386 8732 25442
rect 8788 25386 8812 25442
rect 8868 25386 8893 25442
rect 8949 25386 8974 25442
rect 9030 25386 9055 25442
rect 9111 25386 9136 25442
rect 9192 25386 9217 25442
rect 9273 25386 9298 25442
rect 9354 25386 9379 25442
rect 9435 25386 9460 25442
rect 9516 25386 9541 25442
rect 9597 25386 9622 25442
rect 9678 25386 9703 25442
rect 9759 25386 9767 25442
rect 8567 19362 9767 25386
rect 10866 31883 12066 33373
rect 10866 31827 10871 31883
rect 10927 31827 10951 31883
rect 11007 31827 11031 31883
rect 11087 31827 11111 31883
rect 11167 31827 11192 31883
rect 11248 31827 11273 31883
rect 11329 31827 11354 31883
rect 11410 31827 11435 31883
rect 11491 31827 11516 31883
rect 11572 31827 11597 31883
rect 11653 31827 11678 31883
rect 11734 31827 11759 31883
rect 11815 31827 11840 31883
rect 11896 31827 11921 31883
rect 11977 31827 12002 31883
rect 12058 31827 12066 31883
rect 10866 31795 12066 31827
rect 10866 31739 10871 31795
rect 10927 31739 10951 31795
rect 11007 31739 11031 31795
rect 11087 31739 11111 31795
rect 11167 31739 11192 31795
rect 11248 31739 11273 31795
rect 11329 31739 11354 31795
rect 11410 31739 11435 31795
rect 11491 31739 11516 31795
rect 11572 31739 11597 31795
rect 11653 31739 11678 31795
rect 11734 31739 11759 31795
rect 11815 31739 11840 31795
rect 11896 31739 11921 31795
rect 11977 31739 12002 31795
rect 12058 31739 12066 31795
rect 10866 31707 12066 31739
rect 10866 31651 10871 31707
rect 10927 31651 10951 31707
rect 11007 31651 11031 31707
rect 11087 31651 11111 31707
rect 11167 31651 11192 31707
rect 11248 31651 11273 31707
rect 11329 31651 11354 31707
rect 11410 31651 11435 31707
rect 11491 31651 11516 31707
rect 11572 31651 11597 31707
rect 11653 31651 11678 31707
rect 11734 31651 11759 31707
rect 11815 31651 11840 31707
rect 11896 31651 11921 31707
rect 11977 31651 12002 31707
rect 12058 31651 12066 31707
rect 10866 31619 12066 31651
rect 10866 31563 10871 31619
rect 10927 31563 10951 31619
rect 11007 31563 11031 31619
rect 11087 31563 11111 31619
rect 11167 31563 11192 31619
rect 11248 31563 11273 31619
rect 11329 31563 11354 31619
rect 11410 31563 11435 31619
rect 11491 31563 11516 31619
rect 11572 31563 11597 31619
rect 11653 31563 11678 31619
rect 11734 31563 11759 31619
rect 11815 31563 11840 31619
rect 11896 31563 11921 31619
rect 11977 31563 12002 31619
rect 12058 31563 12066 31619
rect 10866 31531 12066 31563
rect 10866 31475 10871 31531
rect 10927 31475 10951 31531
rect 11007 31475 11031 31531
rect 11087 31475 11111 31531
rect 11167 31475 11192 31531
rect 11248 31475 11273 31531
rect 11329 31475 11354 31531
rect 11410 31475 11435 31531
rect 11491 31475 11516 31531
rect 11572 31475 11597 31531
rect 11653 31475 11678 31531
rect 11734 31475 11759 31531
rect 11815 31475 11840 31531
rect 11896 31475 11921 31531
rect 11977 31475 12002 31531
rect 12058 31475 12066 31531
rect 10866 31443 12066 31475
rect 10866 31387 10871 31443
rect 10927 31387 10951 31443
rect 11007 31387 11031 31443
rect 11087 31387 11111 31443
rect 11167 31387 11192 31443
rect 11248 31387 11273 31443
rect 11329 31387 11354 31443
rect 11410 31387 11435 31443
rect 11491 31387 11516 31443
rect 11572 31387 11597 31443
rect 11653 31387 11678 31443
rect 11734 31387 11759 31443
rect 11815 31387 11840 31443
rect 11896 31387 11921 31443
rect 11977 31387 12002 31443
rect 12058 31387 12066 31443
rect 10866 29883 12066 31387
rect 10866 29827 10871 29883
rect 10927 29827 10951 29883
rect 11007 29827 11031 29883
rect 11087 29827 11111 29883
rect 11167 29827 11192 29883
rect 11248 29827 11273 29883
rect 11329 29827 11354 29883
rect 11410 29827 11435 29883
rect 11491 29827 11516 29883
rect 11572 29827 11597 29883
rect 11653 29827 11678 29883
rect 11734 29827 11759 29883
rect 11815 29827 11840 29883
rect 11896 29827 11921 29883
rect 11977 29827 12002 29883
rect 12058 29827 12066 29883
rect 10866 29795 12066 29827
rect 10866 29739 10871 29795
rect 10927 29739 10951 29795
rect 11007 29739 11031 29795
rect 11087 29739 11111 29795
rect 11167 29739 11192 29795
rect 11248 29739 11273 29795
rect 11329 29739 11354 29795
rect 11410 29739 11435 29795
rect 11491 29739 11516 29795
rect 11572 29739 11597 29795
rect 11653 29739 11678 29795
rect 11734 29739 11759 29795
rect 11815 29739 11840 29795
rect 11896 29739 11921 29795
rect 11977 29739 12002 29795
rect 12058 29739 12066 29795
rect 10866 29707 12066 29739
rect 10866 29651 10871 29707
rect 10927 29651 10951 29707
rect 11007 29651 11031 29707
rect 11087 29651 11111 29707
rect 11167 29651 11192 29707
rect 11248 29651 11273 29707
rect 11329 29651 11354 29707
rect 11410 29651 11435 29707
rect 11491 29651 11516 29707
rect 11572 29651 11597 29707
rect 11653 29651 11678 29707
rect 11734 29651 11759 29707
rect 11815 29651 11840 29707
rect 11896 29651 11921 29707
rect 11977 29651 12002 29707
rect 12058 29651 12066 29707
rect 10866 29619 12066 29651
rect 10866 29563 10871 29619
rect 10927 29563 10951 29619
rect 11007 29563 11031 29619
rect 11087 29563 11111 29619
rect 11167 29563 11192 29619
rect 11248 29563 11273 29619
rect 11329 29563 11354 29619
rect 11410 29563 11435 29619
rect 11491 29563 11516 29619
rect 11572 29563 11597 29619
rect 11653 29563 11678 29619
rect 11734 29563 11759 29619
rect 11815 29563 11840 29619
rect 11896 29563 11921 29619
rect 11977 29563 12002 29619
rect 12058 29563 12066 29619
rect 10866 29531 12066 29563
rect 10866 29475 10871 29531
rect 10927 29475 10951 29531
rect 11007 29475 11031 29531
rect 11087 29475 11111 29531
rect 11167 29475 11192 29531
rect 11248 29475 11273 29531
rect 11329 29475 11354 29531
rect 11410 29475 11435 29531
rect 11491 29475 11516 29531
rect 11572 29475 11597 29531
rect 11653 29475 11678 29531
rect 11734 29475 11759 29531
rect 11815 29475 11840 29531
rect 11896 29475 11921 29531
rect 11977 29475 12002 29531
rect 12058 29475 12066 29531
rect 10866 29443 12066 29475
rect 10866 29387 10871 29443
rect 10927 29387 10951 29443
rect 11007 29387 11031 29443
rect 11087 29387 11111 29443
rect 11167 29387 11192 29443
rect 11248 29387 11273 29443
rect 11329 29387 11354 29443
rect 11410 29387 11435 29443
rect 11491 29387 11516 29443
rect 11572 29387 11597 29443
rect 11653 29387 11678 29443
rect 11734 29387 11759 29443
rect 11815 29387 11840 29443
rect 11896 29387 11921 29443
rect 11977 29387 12002 29443
rect 12058 29387 12066 29443
rect 10866 27883 12066 29387
rect 10866 27827 10871 27883
rect 10927 27827 10951 27883
rect 11007 27827 11031 27883
rect 11087 27827 11111 27883
rect 11167 27827 11192 27883
rect 11248 27827 11273 27883
rect 11329 27827 11354 27883
rect 11410 27827 11435 27883
rect 11491 27827 11516 27883
rect 11572 27827 11597 27883
rect 11653 27827 11678 27883
rect 11734 27827 11759 27883
rect 11815 27827 11840 27883
rect 11896 27827 11921 27883
rect 11977 27827 12002 27883
rect 12058 27827 12066 27883
rect 10866 27795 12066 27827
rect 10866 27739 10871 27795
rect 10927 27739 10951 27795
rect 11007 27739 11031 27795
rect 11087 27739 11111 27795
rect 11167 27739 11192 27795
rect 11248 27739 11273 27795
rect 11329 27739 11354 27795
rect 11410 27739 11435 27795
rect 11491 27739 11516 27795
rect 11572 27739 11597 27795
rect 11653 27739 11678 27795
rect 11734 27739 11759 27795
rect 11815 27739 11840 27795
rect 11896 27739 11921 27795
rect 11977 27739 12002 27795
rect 12058 27739 12066 27795
rect 10866 27707 12066 27739
rect 10866 27651 10871 27707
rect 10927 27651 10951 27707
rect 11007 27651 11031 27707
rect 11087 27651 11111 27707
rect 11167 27651 11192 27707
rect 11248 27651 11273 27707
rect 11329 27651 11354 27707
rect 11410 27651 11435 27707
rect 11491 27651 11516 27707
rect 11572 27651 11597 27707
rect 11653 27651 11678 27707
rect 11734 27651 11759 27707
rect 11815 27651 11840 27707
rect 11896 27651 11921 27707
rect 11977 27651 12002 27707
rect 12058 27651 12066 27707
rect 10866 27619 12066 27651
rect 10866 27563 10871 27619
rect 10927 27563 10951 27619
rect 11007 27563 11031 27619
rect 11087 27563 11111 27619
rect 11167 27563 11192 27619
rect 11248 27563 11273 27619
rect 11329 27563 11354 27619
rect 11410 27563 11435 27619
rect 11491 27563 11516 27619
rect 11572 27563 11597 27619
rect 11653 27563 11678 27619
rect 11734 27563 11759 27619
rect 11815 27563 11840 27619
rect 11896 27563 11921 27619
rect 11977 27563 12002 27619
rect 12058 27563 12066 27619
rect 10866 27531 12066 27563
rect 10866 27475 10871 27531
rect 10927 27475 10951 27531
rect 11007 27475 11031 27531
rect 11087 27475 11111 27531
rect 11167 27475 11192 27531
rect 11248 27475 11273 27531
rect 11329 27475 11354 27531
rect 11410 27475 11435 27531
rect 11491 27475 11516 27531
rect 11572 27475 11597 27531
rect 11653 27475 11678 27531
rect 11734 27475 11759 27531
rect 11815 27475 11840 27531
rect 11896 27475 11921 27531
rect 11977 27475 12002 27531
rect 12058 27475 12066 27531
rect 10866 27443 12066 27475
rect 10866 27387 10871 27443
rect 10927 27387 10951 27443
rect 11007 27387 11031 27443
rect 11087 27387 11111 27443
rect 11167 27387 11192 27443
rect 11248 27387 11273 27443
rect 11329 27387 11354 27443
rect 11410 27387 11435 27443
rect 11491 27387 11516 27443
rect 11572 27387 11597 27443
rect 11653 27387 11678 27443
rect 11734 27387 11759 27443
rect 11815 27387 11840 27443
rect 11896 27387 11921 27443
rect 11977 27387 12002 27443
rect 12058 27387 12066 27443
rect 10866 25882 12066 27387
rect 10866 25826 10871 25882
rect 10927 25826 10951 25882
rect 11007 25826 11031 25882
rect 11087 25826 11111 25882
rect 11167 25826 11192 25882
rect 11248 25826 11273 25882
rect 11329 25826 11354 25882
rect 11410 25826 11435 25882
rect 11491 25826 11516 25882
rect 11572 25826 11597 25882
rect 11653 25826 11678 25882
rect 11734 25826 11759 25882
rect 11815 25826 11840 25882
rect 11896 25826 11921 25882
rect 11977 25826 12002 25882
rect 12058 25826 12066 25882
rect 10866 25794 12066 25826
rect 10866 25738 10871 25794
rect 10927 25738 10951 25794
rect 11007 25738 11031 25794
rect 11087 25738 11111 25794
rect 11167 25738 11192 25794
rect 11248 25738 11273 25794
rect 11329 25738 11354 25794
rect 11410 25738 11435 25794
rect 11491 25738 11516 25794
rect 11572 25738 11597 25794
rect 11653 25738 11678 25794
rect 11734 25738 11759 25794
rect 11815 25738 11840 25794
rect 11896 25738 11921 25794
rect 11977 25738 12002 25794
rect 12058 25738 12066 25794
rect 10866 25706 12066 25738
rect 10866 25650 10871 25706
rect 10927 25650 10951 25706
rect 11007 25650 11031 25706
rect 11087 25650 11111 25706
rect 11167 25650 11192 25706
rect 11248 25650 11273 25706
rect 11329 25650 11354 25706
rect 11410 25650 11435 25706
rect 11491 25650 11516 25706
rect 11572 25650 11597 25706
rect 11653 25650 11678 25706
rect 11734 25650 11759 25706
rect 11815 25650 11840 25706
rect 11896 25650 11921 25706
rect 11977 25650 12002 25706
rect 12058 25650 12066 25706
rect 10866 25618 12066 25650
rect 10866 25562 10871 25618
rect 10927 25562 10951 25618
rect 11007 25562 11031 25618
rect 11087 25562 11111 25618
rect 11167 25562 11192 25618
rect 11248 25562 11273 25618
rect 11329 25562 11354 25618
rect 11410 25562 11435 25618
rect 11491 25562 11516 25618
rect 11572 25562 11597 25618
rect 11653 25562 11678 25618
rect 11734 25562 11759 25618
rect 11815 25562 11840 25618
rect 11896 25562 11921 25618
rect 11977 25562 12002 25618
rect 12058 25562 12066 25618
rect 10866 25530 12066 25562
rect 10866 25474 10871 25530
rect 10927 25474 10951 25530
rect 11007 25474 11031 25530
rect 11087 25474 11111 25530
rect 11167 25474 11192 25530
rect 11248 25474 11273 25530
rect 11329 25474 11354 25530
rect 11410 25474 11435 25530
rect 11491 25474 11516 25530
rect 11572 25474 11597 25530
rect 11653 25474 11678 25530
rect 11734 25474 11759 25530
rect 11815 25474 11840 25530
rect 11896 25474 11921 25530
rect 11977 25474 12002 25530
rect 12058 25474 12066 25530
rect 10866 25442 12066 25474
rect 10866 25386 10871 25442
rect 10927 25386 10951 25442
rect 11007 25386 11031 25442
rect 11087 25386 11111 25442
rect 11167 25386 11192 25442
rect 11248 25386 11273 25442
rect 11329 25386 11354 25442
rect 11410 25386 11435 25442
rect 11491 25386 11516 25442
rect 11572 25386 11597 25442
rect 11653 25386 11678 25442
rect 11734 25386 11759 25442
rect 11815 25386 11840 25442
rect 11896 25386 11921 25442
rect 11977 25386 12002 25442
rect 12058 25386 12066 25442
tri 10195 19362 10866 20033 se
rect 10866 19537 12066 25386
rect 10866 19362 11891 19537
tri 11891 19362 12066 19537 nw
rect 12409 34197 14940 34447
rect 12409 34133 12446 34197
rect 12510 34133 12554 34197
rect 12618 34133 14940 34197
rect 12409 34089 14940 34133
rect 12409 34025 12446 34089
rect 12510 34025 12554 34089
rect 12618 34045 14940 34089
rect 12618 34025 12646 34045
rect 12409 33981 12646 34025
rect 12710 33981 12737 34045
rect 12801 33981 12828 34045
rect 12892 33981 14940 34045
rect 12409 33917 12446 33981
rect 12510 33917 12554 33981
rect 12618 33917 14940 33981
rect 12409 33915 14940 33917
rect 12409 33897 12950 33915
rect 12409 33872 12646 33897
rect 12409 33808 12446 33872
rect 12510 33808 12554 33872
rect 12618 33833 12646 33872
rect 12710 33833 12737 33897
rect 12801 33833 12828 33897
rect 12892 33851 12950 33897
rect 13014 33851 14940 33915
rect 12892 33833 14940 33851
rect 12618 33808 14940 33833
rect 12409 33800 14940 33808
rect 12409 33763 12648 33800
rect 12409 33699 12446 33763
rect 12510 33699 12554 33763
rect 12618 33736 12648 33763
rect 12712 33736 12777 33800
rect 12841 33736 12906 33800
rect 12970 33736 13034 33800
rect 13098 33736 14940 33800
rect 12618 33699 14940 33736
rect 12409 33698 14940 33699
rect 12409 33634 12648 33698
rect 12712 33634 12777 33698
rect 12841 33634 12906 33698
rect 12970 33634 13034 33698
rect 13098 33683 14940 33698
rect 13098 33634 13182 33683
rect 12409 33619 13182 33634
rect 13246 33619 14940 33683
rect 12409 33594 14940 33619
rect 12409 33564 12870 33594
rect 12409 33500 12728 33564
rect 12792 33530 12870 33564
rect 12934 33530 12951 33594
rect 13015 33530 13033 33594
rect 13097 33530 13115 33594
rect 13179 33530 13197 33594
rect 13261 33530 13279 33594
rect 13343 33530 14940 33594
rect 12792 33500 14940 33530
rect 12409 33468 14940 33500
rect 12409 33446 13397 33468
rect 12409 33382 12870 33446
rect 12934 33382 12951 33446
rect 13015 33382 13033 33446
rect 13097 33382 13115 33446
rect 13179 33382 13197 33446
rect 13261 33382 13279 33446
rect 13343 33404 13397 33446
rect 13461 33404 14940 33468
rect 13343 33382 14940 33404
rect 12409 33366 14940 33382
rect 12409 33349 13068 33366
rect 12409 33285 12943 33349
rect 13007 33302 13068 33349
rect 13132 33302 13149 33366
rect 13213 33302 13231 33366
rect 13295 33302 13313 33366
rect 13377 33302 13395 33366
rect 13459 33302 13477 33366
rect 13541 33302 14940 33366
rect 13007 33285 14940 33302
rect 12409 33229 14940 33285
rect 12409 33218 13636 33229
rect 12409 33154 13068 33218
rect 13132 33154 13149 33218
rect 13213 33154 13231 33218
rect 13295 33154 13313 33218
rect 13377 33154 13395 33218
rect 13459 33154 13477 33218
rect 13541 33165 13636 33218
rect 13700 33165 14940 33229
rect 13541 33154 14940 33165
rect 12409 33138 14940 33154
rect 12409 33110 13324 33138
rect 12409 33046 13182 33110
rect 13246 33074 13324 33110
rect 13388 33074 13405 33138
rect 13469 33074 13487 33138
rect 13551 33074 13569 33138
rect 13633 33074 13651 33138
rect 13715 33074 13733 33138
rect 13797 33074 14940 33138
rect 13246 33046 14940 33074
rect 12409 33006 14940 33046
rect 12409 32990 13859 33006
rect 12409 32926 13324 32990
rect 13388 32926 13405 32990
rect 13469 32926 13487 32990
rect 13551 32926 13569 32990
rect 13633 32926 13651 32990
rect 13715 32926 13733 32990
rect 13797 32942 13859 32990
rect 13923 32942 14940 33006
rect 13797 32926 14940 32942
rect 12409 32887 14940 32926
rect 12409 32823 13405 32887
rect 13469 32869 14940 32887
rect 13469 32823 13506 32869
rect 12409 32805 13506 32823
rect 13570 32805 13598 32869
rect 13662 32805 13690 32869
rect 13754 32805 13782 32869
rect 13846 32805 13874 32869
rect 13938 32805 13966 32869
rect 14030 32805 14940 32869
rect 12409 32789 14940 32805
rect 12409 32725 13506 32789
rect 13570 32725 13598 32789
rect 13662 32725 13690 32789
rect 13754 32725 13782 32789
rect 13846 32725 13874 32789
rect 13938 32725 13966 32789
rect 14030 32725 14940 32789
rect 12409 32709 14940 32725
rect 12409 32645 13506 32709
rect 13570 32645 13598 32709
rect 13662 32645 13690 32709
rect 13754 32645 13782 32709
rect 13846 32645 13874 32709
rect 13938 32645 13966 32709
rect 14030 32645 14940 32709
rect 12409 32629 14940 32645
rect 12409 32565 13506 32629
rect 13570 32565 13598 32629
rect 13662 32565 13690 32629
rect 13754 32565 13782 32629
rect 13846 32565 13874 32629
rect 13938 32565 13966 32629
rect 14030 32565 14940 32629
rect 12409 32549 14940 32565
rect 12409 32485 13506 32549
rect 13570 32485 13598 32549
rect 13662 32485 13690 32549
rect 13754 32485 13782 32549
rect 13846 32485 13874 32549
rect 13938 32485 13966 32549
rect 14030 32485 14940 32549
rect 12409 32469 14940 32485
rect 12409 32405 13506 32469
rect 13570 32405 13598 32469
rect 13662 32405 13690 32469
rect 13754 32405 13782 32469
rect 13846 32405 13874 32469
rect 13938 32405 13966 32469
rect 14030 32405 14940 32469
rect 12409 32389 14940 32405
rect 12409 32325 13506 32389
rect 13570 32325 13598 32389
rect 13662 32325 13690 32389
rect 13754 32325 13782 32389
rect 13846 32325 13874 32389
rect 13938 32325 13966 32389
rect 14030 32325 14940 32389
rect 12409 32309 14940 32325
rect 12409 32245 13506 32309
rect 13570 32245 13598 32309
rect 13662 32245 13690 32309
rect 13754 32245 13782 32309
rect 13846 32245 13874 32309
rect 13938 32245 13966 32309
rect 14030 32245 14940 32309
rect 12409 32229 14940 32245
rect 12409 32165 13506 32229
rect 13570 32165 13598 32229
rect 13662 32165 13690 32229
rect 13754 32165 13782 32229
rect 13846 32165 13874 32229
rect 13938 32165 13966 32229
rect 14030 32165 14940 32229
rect 12409 32149 14940 32165
rect 12409 32085 13506 32149
rect 13570 32085 13598 32149
rect 13662 32085 13690 32149
rect 13754 32085 13782 32149
rect 13846 32085 13874 32149
rect 13938 32085 13966 32149
rect 14030 32085 14940 32149
rect 12409 32069 14940 32085
rect 12409 32005 13506 32069
rect 13570 32005 13598 32069
rect 13662 32005 13690 32069
rect 13754 32005 13782 32069
rect 13846 32005 13874 32069
rect 13938 32005 13966 32069
rect 14030 32005 14940 32069
rect 12409 31989 14940 32005
rect 12409 31925 13506 31989
rect 13570 31925 13598 31989
rect 13662 31925 13690 31989
rect 13754 31925 13782 31989
rect 13846 31925 13874 31989
rect 13938 31925 13966 31989
rect 14030 31925 14940 31989
rect 12409 31909 14940 31925
rect 12409 31845 13506 31909
rect 13570 31845 13598 31909
rect 13662 31845 13690 31909
rect 13754 31845 13782 31909
rect 13846 31845 13874 31909
rect 13938 31845 13966 31909
rect 14030 31845 14940 31909
rect 12409 31829 14940 31845
rect 12409 31765 13506 31829
rect 13570 31765 13598 31829
rect 13662 31765 13690 31829
rect 13754 31765 13782 31829
rect 13846 31765 13874 31829
rect 13938 31765 13966 31829
rect 14030 31765 14940 31829
rect 12409 31749 14940 31765
rect 12409 31685 13506 31749
rect 13570 31685 13598 31749
rect 13662 31685 13690 31749
rect 13754 31685 13782 31749
rect 13846 31685 13874 31749
rect 13938 31685 13966 31749
rect 14030 31685 14940 31749
rect 12409 31669 14940 31685
rect 12409 31605 13506 31669
rect 13570 31605 13598 31669
rect 13662 31605 13690 31669
rect 13754 31605 13782 31669
rect 13846 31605 13874 31669
rect 13938 31605 13966 31669
rect 14030 31605 14940 31669
rect 12409 31589 14940 31605
rect 12409 31525 13506 31589
rect 13570 31525 13598 31589
rect 13662 31525 13690 31589
rect 13754 31525 13782 31589
rect 13846 31525 13874 31589
rect 13938 31525 13966 31589
rect 14030 31525 14940 31589
rect 12409 31509 14940 31525
rect 12409 31445 13506 31509
rect 13570 31445 13598 31509
rect 13662 31445 13690 31509
rect 13754 31445 13782 31509
rect 13846 31445 13874 31509
rect 13938 31445 13966 31509
rect 14030 31445 14940 31509
rect 12409 31429 14940 31445
rect 12409 31365 13506 31429
rect 13570 31365 13598 31429
rect 13662 31365 13690 31429
rect 13754 31365 13782 31429
rect 13846 31365 13874 31429
rect 13938 31365 13966 31429
rect 14030 31365 14940 31429
rect 12409 31349 14940 31365
rect 12409 31285 13506 31349
rect 13570 31285 13598 31349
rect 13662 31285 13690 31349
rect 13754 31285 13782 31349
rect 13846 31285 13874 31349
rect 13938 31285 13966 31349
rect 14030 31285 14940 31349
rect 12409 31269 14940 31285
rect 12409 31205 13506 31269
rect 13570 31205 13598 31269
rect 13662 31205 13690 31269
rect 13754 31205 13782 31269
rect 13846 31205 13874 31269
rect 13938 31205 13966 31269
rect 14030 31205 14940 31269
rect 12409 31189 14940 31205
rect 12409 31125 13506 31189
rect 13570 31125 13598 31189
rect 13662 31125 13690 31189
rect 13754 31125 13782 31189
rect 13846 31125 13874 31189
rect 13938 31125 13966 31189
rect 14030 31125 14940 31189
rect 12409 31109 14940 31125
rect 12409 31045 13506 31109
rect 13570 31045 13598 31109
rect 13662 31045 13690 31109
rect 13754 31045 13782 31109
rect 13846 31045 13874 31109
rect 13938 31045 13966 31109
rect 14030 31045 14940 31109
rect 12409 31029 14940 31045
rect 12409 30965 13506 31029
rect 13570 30965 13598 31029
rect 13662 30965 13690 31029
rect 13754 30965 13782 31029
rect 13846 30965 13874 31029
rect 13938 30965 13966 31029
rect 14030 30965 14940 31029
rect 12409 30949 14940 30965
rect 12409 30885 13506 30949
rect 13570 30885 13598 30949
rect 13662 30885 13690 30949
rect 13754 30885 13782 30949
rect 13846 30885 13874 30949
rect 13938 30885 13966 30949
rect 14030 30885 14940 30949
rect 12409 30869 14940 30885
rect 12409 30805 13506 30869
rect 13570 30805 13598 30869
rect 13662 30805 13690 30869
rect 13754 30805 13782 30869
rect 13846 30805 13874 30869
rect 13938 30805 13966 30869
rect 14030 30805 14940 30869
rect 12409 30789 14940 30805
rect 12409 30725 13506 30789
rect 13570 30725 13598 30789
rect 13662 30725 13690 30789
rect 13754 30725 13782 30789
rect 13846 30725 13874 30789
rect 13938 30725 13966 30789
rect 14030 30725 14940 30789
rect 12409 30709 14940 30725
rect 12409 30645 13506 30709
rect 13570 30645 13598 30709
rect 13662 30645 13690 30709
rect 13754 30645 13782 30709
rect 13846 30645 13874 30709
rect 13938 30645 13966 30709
rect 14030 30645 14940 30709
rect 12409 30629 14940 30645
rect 12409 30565 13506 30629
rect 13570 30565 13598 30629
rect 13662 30565 13690 30629
rect 13754 30565 13782 30629
rect 13846 30565 13874 30629
rect 13938 30565 13966 30629
rect 14030 30565 14940 30629
rect 12409 30549 14940 30565
rect 12409 30485 13506 30549
rect 13570 30485 13598 30549
rect 13662 30485 13690 30549
rect 13754 30485 13782 30549
rect 13846 30485 13874 30549
rect 13938 30485 13966 30549
rect 14030 30485 14940 30549
rect 12409 30469 14940 30485
rect 12409 30405 13506 30469
rect 13570 30405 13598 30469
rect 13662 30405 13690 30469
rect 13754 30405 13782 30469
rect 13846 30405 13874 30469
rect 13938 30405 13966 30469
rect 14030 30405 14940 30469
rect 12409 30389 14940 30405
rect 12409 30325 13506 30389
rect 13570 30325 13598 30389
rect 13662 30325 13690 30389
rect 13754 30325 13782 30389
rect 13846 30325 13874 30389
rect 13938 30325 13966 30389
rect 14030 30325 14940 30389
rect 12409 30309 14940 30325
rect 12409 30245 13506 30309
rect 13570 30245 13598 30309
rect 13662 30245 13690 30309
rect 13754 30245 13782 30309
rect 13846 30245 13874 30309
rect 13938 30245 13966 30309
rect 14030 30245 14940 30309
rect 12409 30229 14940 30245
rect 12409 30165 13506 30229
rect 13570 30165 13598 30229
rect 13662 30165 13690 30229
rect 13754 30165 13782 30229
rect 13846 30165 13874 30229
rect 13938 30165 13966 30229
rect 14030 30165 14940 30229
rect 12409 30149 14940 30165
rect 12409 30085 13506 30149
rect 13570 30085 13598 30149
rect 13662 30085 13690 30149
rect 13754 30085 13782 30149
rect 13846 30085 13874 30149
rect 13938 30085 13966 30149
rect 14030 30085 14940 30149
rect 12409 30069 14940 30085
rect 12409 30005 13506 30069
rect 13570 30005 13598 30069
rect 13662 30005 13690 30069
rect 13754 30005 13782 30069
rect 13846 30005 13874 30069
rect 13938 30005 13966 30069
rect 14030 30005 14940 30069
rect 12409 29989 14940 30005
rect 12409 29925 13506 29989
rect 13570 29925 13598 29989
rect 13662 29925 13690 29989
rect 13754 29925 13782 29989
rect 13846 29925 13874 29989
rect 13938 29925 13966 29989
rect 14030 29925 14940 29989
rect 12409 29909 14940 29925
rect 12409 29845 13506 29909
rect 13570 29845 13598 29909
rect 13662 29845 13690 29909
rect 13754 29845 13782 29909
rect 13846 29845 13874 29909
rect 13938 29845 13966 29909
rect 14030 29845 14940 29909
rect 12409 29829 14940 29845
rect 12409 29765 13506 29829
rect 13570 29765 13598 29829
rect 13662 29765 13690 29829
rect 13754 29765 13782 29829
rect 13846 29765 13874 29829
rect 13938 29765 13966 29829
rect 14030 29765 14940 29829
rect 12409 29749 14940 29765
rect 12409 29685 13506 29749
rect 13570 29685 13598 29749
rect 13662 29685 13690 29749
rect 13754 29685 13782 29749
rect 13846 29685 13874 29749
rect 13938 29685 13966 29749
rect 14030 29685 14940 29749
rect 12409 29669 14940 29685
rect 12409 29605 13506 29669
rect 13570 29605 13598 29669
rect 13662 29605 13690 29669
rect 13754 29605 13782 29669
rect 13846 29605 13874 29669
rect 13938 29605 13966 29669
rect 14030 29605 14940 29669
rect 12409 29589 14940 29605
rect 12409 29525 13506 29589
rect 13570 29525 13598 29589
rect 13662 29525 13690 29589
rect 13754 29525 13782 29589
rect 13846 29525 13874 29589
rect 13938 29525 13966 29589
rect 14030 29525 14940 29589
rect 12409 29509 14940 29525
rect 12409 29445 13506 29509
rect 13570 29445 13598 29509
rect 13662 29445 13690 29509
rect 13754 29445 13782 29509
rect 13846 29445 13874 29509
rect 13938 29445 13966 29509
rect 14030 29445 14940 29509
rect 12409 29429 14940 29445
rect 12409 29365 13506 29429
rect 13570 29365 13598 29429
rect 13662 29365 13690 29429
rect 13754 29365 13782 29429
rect 13846 29365 13874 29429
rect 13938 29365 13966 29429
rect 14030 29365 14940 29429
rect 12409 29349 14940 29365
rect 12409 29285 13506 29349
rect 13570 29285 13598 29349
rect 13662 29285 13690 29349
rect 13754 29285 13782 29349
rect 13846 29285 13874 29349
rect 13938 29285 13966 29349
rect 14030 29285 14940 29349
rect 12409 29269 14940 29285
rect 12409 29205 13506 29269
rect 13570 29205 13598 29269
rect 13662 29205 13690 29269
rect 13754 29205 13782 29269
rect 13846 29205 13874 29269
rect 13938 29205 13966 29269
rect 14030 29205 14940 29269
rect 12409 29189 14940 29205
rect 12409 29125 13506 29189
rect 13570 29125 13598 29189
rect 13662 29125 13690 29189
rect 13754 29125 13782 29189
rect 13846 29125 13874 29189
rect 13938 29125 13966 29189
rect 14030 29125 14940 29189
rect 12409 29109 14940 29125
rect 12409 29045 13506 29109
rect 13570 29045 13598 29109
rect 13662 29045 13690 29109
rect 13754 29045 13782 29109
rect 13846 29045 13874 29109
rect 13938 29045 13966 29109
rect 14030 29045 14940 29109
rect 12409 29029 14940 29045
rect 12409 28965 13506 29029
rect 13570 28965 13598 29029
rect 13662 28965 13690 29029
rect 13754 28965 13782 29029
rect 13846 28965 13874 29029
rect 13938 28965 13966 29029
rect 14030 28965 14940 29029
rect 12409 28949 14940 28965
rect 12409 28885 13506 28949
rect 13570 28885 13598 28949
rect 13662 28885 13690 28949
rect 13754 28885 13782 28949
rect 13846 28885 13874 28949
rect 13938 28885 13966 28949
rect 14030 28885 14940 28949
rect 12409 28869 14940 28885
rect 12409 28805 13506 28869
rect 13570 28805 13598 28869
rect 13662 28805 13690 28869
rect 13754 28805 13782 28869
rect 13846 28805 13874 28869
rect 13938 28805 13966 28869
rect 14030 28805 14940 28869
rect 12409 28789 14940 28805
rect 12409 28725 13506 28789
rect 13570 28725 13598 28789
rect 13662 28725 13690 28789
rect 13754 28725 13782 28789
rect 13846 28725 13874 28789
rect 13938 28725 13966 28789
rect 14030 28725 14940 28789
rect 12409 28709 14940 28725
rect 12409 28645 13506 28709
rect 13570 28645 13598 28709
rect 13662 28645 13690 28709
rect 13754 28645 13782 28709
rect 13846 28645 13874 28709
rect 13938 28645 13966 28709
rect 14030 28645 14940 28709
rect 12409 28629 14940 28645
rect 12409 28565 13506 28629
rect 13570 28565 13598 28629
rect 13662 28565 13690 28629
rect 13754 28565 13782 28629
rect 13846 28565 13874 28629
rect 13938 28565 13966 28629
rect 14030 28565 14940 28629
rect 12409 28549 14940 28565
rect 12409 28485 13506 28549
rect 13570 28485 13598 28549
rect 13662 28485 13690 28549
rect 13754 28485 13782 28549
rect 13846 28485 13874 28549
rect 13938 28485 13966 28549
rect 14030 28485 14940 28549
rect 12409 28469 14940 28485
rect 12409 28405 13506 28469
rect 13570 28405 13598 28469
rect 13662 28405 13690 28469
rect 13754 28405 13782 28469
rect 13846 28405 13874 28469
rect 13938 28405 13966 28469
rect 14030 28405 14940 28469
rect 12409 28389 14940 28405
rect 12409 28325 13506 28389
rect 13570 28325 13598 28389
rect 13662 28325 13690 28389
rect 13754 28325 13782 28389
rect 13846 28325 13874 28389
rect 13938 28325 13966 28389
rect 14030 28325 14940 28389
rect 12409 28309 14940 28325
rect 12409 28245 13506 28309
rect 13570 28245 13598 28309
rect 13662 28245 13690 28309
rect 13754 28245 13782 28309
rect 13846 28245 13874 28309
rect 13938 28245 13966 28309
rect 14030 28245 14940 28309
rect 12409 28229 14940 28245
rect 12409 28165 13506 28229
rect 13570 28165 13598 28229
rect 13662 28165 13690 28229
rect 13754 28165 13782 28229
rect 13846 28165 13874 28229
rect 13938 28165 13966 28229
rect 14030 28165 14940 28229
rect 12409 28149 14940 28165
rect 12409 28085 13506 28149
rect 13570 28085 13598 28149
rect 13662 28085 13690 28149
rect 13754 28085 13782 28149
rect 13846 28085 13874 28149
rect 13938 28085 13966 28149
rect 14030 28085 14940 28149
rect 12409 28069 14940 28085
rect 12409 28005 13506 28069
rect 13570 28005 13598 28069
rect 13662 28005 13690 28069
rect 13754 28005 13782 28069
rect 13846 28005 13874 28069
rect 13938 28005 13966 28069
rect 14030 28005 14940 28069
rect 12409 27989 14940 28005
rect 12409 27925 13506 27989
rect 13570 27925 13598 27989
rect 13662 27925 13690 27989
rect 13754 27925 13782 27989
rect 13846 27925 13874 27989
rect 13938 27925 13966 27989
rect 14030 27925 14940 27989
rect 12409 27909 14940 27925
rect 12409 27845 13506 27909
rect 13570 27845 13598 27909
rect 13662 27845 13690 27909
rect 13754 27845 13782 27909
rect 13846 27845 13874 27909
rect 13938 27845 13966 27909
rect 14030 27845 14940 27909
rect 12409 27829 14940 27845
rect 12409 27765 13506 27829
rect 13570 27765 13598 27829
rect 13662 27765 13690 27829
rect 13754 27765 13782 27829
rect 13846 27765 13874 27829
rect 13938 27765 13966 27829
rect 14030 27765 14940 27829
rect 12409 27749 14940 27765
rect 12409 27685 13506 27749
rect 13570 27685 13598 27749
rect 13662 27685 13690 27749
rect 13754 27685 13782 27749
rect 13846 27685 13874 27749
rect 13938 27685 13966 27749
rect 14030 27685 14940 27749
rect 12409 27669 14940 27685
rect 12409 27605 13506 27669
rect 13570 27605 13598 27669
rect 13662 27605 13690 27669
rect 13754 27605 13782 27669
rect 13846 27605 13874 27669
rect 13938 27605 13966 27669
rect 14030 27605 14940 27669
rect 12409 27589 14940 27605
rect 12409 27525 13506 27589
rect 13570 27525 13598 27589
rect 13662 27525 13690 27589
rect 13754 27525 13782 27589
rect 13846 27525 13874 27589
rect 13938 27525 13966 27589
rect 14030 27525 14940 27589
rect 12409 27509 14940 27525
rect 12409 27445 13506 27509
rect 13570 27445 13598 27509
rect 13662 27445 13690 27509
rect 13754 27445 13782 27509
rect 13846 27445 13874 27509
rect 13938 27445 13966 27509
rect 14030 27445 14940 27509
rect 12409 27429 14940 27445
rect 12409 27365 13506 27429
rect 13570 27365 13598 27429
rect 13662 27365 13690 27429
rect 13754 27365 13782 27429
rect 13846 27365 13874 27429
rect 13938 27365 13966 27429
rect 14030 27365 14940 27429
rect 12409 27349 14940 27365
rect 12409 27285 13506 27349
rect 13570 27285 13598 27349
rect 13662 27285 13690 27349
rect 13754 27285 13782 27349
rect 13846 27285 13874 27349
rect 13938 27285 13966 27349
rect 14030 27285 14940 27349
rect 12409 27269 14940 27285
rect 12409 27205 13506 27269
rect 13570 27205 13598 27269
rect 13662 27205 13690 27269
rect 13754 27205 13782 27269
rect 13846 27205 13874 27269
rect 13938 27205 13966 27269
rect 14030 27205 14940 27269
rect 12409 27189 14940 27205
rect 12409 27125 13506 27189
rect 13570 27125 13598 27189
rect 13662 27125 13690 27189
rect 13754 27125 13782 27189
rect 13846 27125 13874 27189
rect 13938 27125 13966 27189
rect 14030 27125 14940 27189
rect 12409 27109 14940 27125
rect 12409 27045 13506 27109
rect 13570 27045 13598 27109
rect 13662 27045 13690 27109
rect 13754 27045 13782 27109
rect 13846 27045 13874 27109
rect 13938 27045 13966 27109
rect 14030 27045 14940 27109
rect 12409 27029 14940 27045
rect 12409 26965 13506 27029
rect 13570 26965 13598 27029
rect 13662 26965 13690 27029
rect 13754 26965 13782 27029
rect 13846 26965 13874 27029
rect 13938 26965 13966 27029
rect 14030 26965 14940 27029
rect 12409 26949 14940 26965
rect 12409 26885 13506 26949
rect 13570 26885 13598 26949
rect 13662 26885 13690 26949
rect 13754 26885 13782 26949
rect 13846 26885 13874 26949
rect 13938 26885 13966 26949
rect 14030 26885 14940 26949
rect 12409 26869 14940 26885
rect 12409 26805 13506 26869
rect 13570 26805 13598 26869
rect 13662 26805 13690 26869
rect 13754 26805 13782 26869
rect 13846 26805 13874 26869
rect 13938 26805 13966 26869
rect 14030 26805 14940 26869
rect 12409 26789 14940 26805
rect 12409 26725 13506 26789
rect 13570 26725 13598 26789
rect 13662 26725 13690 26789
rect 13754 26725 13782 26789
rect 13846 26725 13874 26789
rect 13938 26725 13966 26789
rect 14030 26725 14940 26789
rect 12409 26709 14940 26725
rect 12409 26645 13506 26709
rect 13570 26645 13598 26709
rect 13662 26645 13690 26709
rect 13754 26645 13782 26709
rect 13846 26645 13874 26709
rect 13938 26645 13966 26709
rect 14030 26645 14940 26709
rect 12409 26629 14940 26645
rect 12409 26565 13506 26629
rect 13570 26565 13598 26629
rect 13662 26565 13690 26629
rect 13754 26565 13782 26629
rect 13846 26565 13874 26629
rect 13938 26565 13966 26629
rect 14030 26565 14940 26629
rect 12409 26549 14940 26565
rect 12409 26485 13506 26549
rect 13570 26485 13598 26549
rect 13662 26485 13690 26549
rect 13754 26485 13782 26549
rect 13846 26485 13874 26549
rect 13938 26485 13966 26549
rect 14030 26485 14940 26549
rect 12409 26469 14940 26485
rect 12409 26405 13506 26469
rect 13570 26405 13598 26469
rect 13662 26405 13690 26469
rect 13754 26405 13782 26469
rect 13846 26405 13874 26469
rect 13938 26405 13966 26469
rect 14030 26405 14940 26469
rect 12409 26389 14940 26405
rect 12409 26325 13506 26389
rect 13570 26325 13598 26389
rect 13662 26325 13690 26389
rect 13754 26325 13782 26389
rect 13846 26325 13874 26389
rect 13938 26325 13966 26389
rect 14030 26325 14940 26389
rect 12409 26309 14940 26325
rect 12409 26245 13506 26309
rect 13570 26245 13598 26309
rect 13662 26245 13690 26309
rect 13754 26245 13782 26309
rect 13846 26245 13874 26309
rect 13938 26245 13966 26309
rect 14030 26245 14940 26309
rect 12409 26229 14940 26245
rect 12409 26165 13506 26229
rect 13570 26165 13598 26229
rect 13662 26165 13690 26229
rect 13754 26165 13782 26229
rect 13846 26165 13874 26229
rect 13938 26165 13966 26229
rect 14030 26165 14940 26229
rect 12409 26149 14940 26165
rect 12409 26085 13506 26149
rect 13570 26085 13598 26149
rect 13662 26085 13690 26149
rect 13754 26085 13782 26149
rect 13846 26085 13874 26149
rect 13938 26085 13966 26149
rect 14030 26085 14940 26149
rect 12409 26069 14940 26085
rect 12409 26005 13506 26069
rect 13570 26005 13598 26069
rect 13662 26005 13690 26069
rect 13754 26005 13782 26069
rect 13846 26005 13874 26069
rect 13938 26005 13966 26069
rect 14030 26005 14940 26069
rect 12409 25989 14940 26005
rect 12409 25925 13506 25989
rect 13570 25925 13598 25989
rect 13662 25925 13690 25989
rect 13754 25925 13782 25989
rect 13846 25925 13874 25989
rect 13938 25925 13966 25989
rect 14030 25925 14940 25989
rect 12409 25909 14940 25925
rect 12409 25845 13506 25909
rect 13570 25845 13598 25909
rect 13662 25845 13690 25909
rect 13754 25845 13782 25909
rect 13846 25845 13874 25909
rect 13938 25845 13966 25909
rect 14030 25845 14940 25909
rect 12409 25829 14940 25845
rect 12409 25765 13506 25829
rect 13570 25765 13598 25829
rect 13662 25765 13690 25829
rect 13754 25765 13782 25829
rect 13846 25765 13874 25829
rect 13938 25765 13966 25829
rect 14030 25765 14940 25829
rect 12409 25749 14940 25765
rect 12409 25685 13506 25749
rect 13570 25685 13598 25749
rect 13662 25685 13690 25749
rect 13754 25685 13782 25749
rect 13846 25685 13874 25749
rect 13938 25685 13966 25749
rect 14030 25685 14940 25749
rect 12409 25669 14940 25685
rect 12409 25605 13506 25669
rect 13570 25605 13598 25669
rect 13662 25605 13690 25669
rect 13754 25605 13782 25669
rect 13846 25605 13874 25669
rect 13938 25605 13966 25669
rect 14030 25605 14940 25669
rect 12409 25589 14940 25605
rect 12409 25525 13506 25589
rect 13570 25525 13598 25589
rect 13662 25525 13690 25589
rect 13754 25525 13782 25589
rect 13846 25525 13874 25589
rect 13938 25525 13966 25589
rect 14030 25525 14940 25589
rect 12409 25509 14940 25525
rect 12409 25445 13506 25509
rect 13570 25445 13598 25509
rect 13662 25445 13690 25509
rect 13754 25445 13782 25509
rect 13846 25445 13874 25509
rect 13938 25445 13966 25509
rect 14030 25445 14940 25509
rect 12409 25429 14940 25445
rect 12409 25365 13506 25429
rect 13570 25365 13598 25429
rect 13662 25365 13690 25429
rect 13754 25365 13782 25429
rect 13846 25365 13874 25429
rect 13938 25365 13966 25429
rect 14030 25365 14940 25429
rect 12409 25349 14940 25365
rect 12409 25285 13506 25349
rect 13570 25285 13598 25349
rect 13662 25285 13690 25349
rect 13754 25285 13782 25349
rect 13846 25285 13874 25349
rect 13938 25285 13966 25349
rect 14030 25285 14940 25349
rect 12409 25269 14940 25285
rect 12409 25205 13506 25269
rect 13570 25205 13598 25269
rect 13662 25205 13690 25269
rect 13754 25205 13782 25269
rect 13846 25205 13874 25269
rect 13938 25205 13966 25269
rect 14030 25205 14940 25269
rect 12409 25189 14940 25205
rect 12409 25125 13506 25189
rect 13570 25125 13598 25189
rect 13662 25125 13690 25189
rect 13754 25125 13782 25189
rect 13846 25125 13874 25189
rect 13938 25125 13966 25189
rect 14030 25125 14940 25189
rect 12409 25109 14940 25125
rect 12409 25045 13506 25109
rect 13570 25045 13598 25109
rect 13662 25045 13690 25109
rect 13754 25045 13782 25109
rect 13846 25045 13874 25109
rect 13938 25045 13966 25109
rect 14030 25045 14940 25109
rect 12409 25029 14940 25045
rect 12409 24965 13506 25029
rect 13570 24965 13598 25029
rect 13662 24965 13690 25029
rect 13754 24965 13782 25029
rect 13846 24965 13874 25029
rect 13938 24965 13966 25029
rect 14030 24965 14940 25029
rect 12409 24949 14940 24965
rect 12409 24885 13506 24949
rect 13570 24885 13598 24949
rect 13662 24885 13690 24949
rect 13754 24885 13782 24949
rect 13846 24885 13874 24949
rect 13938 24885 13966 24949
rect 14030 24885 14940 24949
rect 12409 24869 14940 24885
rect 12409 24805 13506 24869
rect 13570 24805 13598 24869
rect 13662 24805 13690 24869
rect 13754 24805 13782 24869
rect 13846 24805 13874 24869
rect 13938 24805 13966 24869
rect 14030 24805 14940 24869
rect 12409 24789 14940 24805
rect 12409 24725 13506 24789
rect 13570 24725 13598 24789
rect 13662 24725 13690 24789
rect 13754 24725 13782 24789
rect 13846 24725 13874 24789
rect 13938 24725 13966 24789
rect 14030 24725 14940 24789
rect 12409 24709 14940 24725
rect 12409 24645 13506 24709
rect 13570 24645 13598 24709
rect 13662 24645 13690 24709
rect 13754 24645 13782 24709
rect 13846 24645 13874 24709
rect 13938 24645 13966 24709
rect 14030 24645 14940 24709
rect 12409 24629 14940 24645
rect 12409 24565 13506 24629
rect 13570 24565 13598 24629
rect 13662 24565 13690 24629
rect 13754 24565 13782 24629
rect 13846 24565 13874 24629
rect 13938 24565 13966 24629
rect 14030 24565 14940 24629
rect 12409 24549 14940 24565
rect 12409 24485 13506 24549
rect 13570 24485 13598 24549
rect 13662 24485 13690 24549
rect 13754 24485 13782 24549
rect 13846 24485 13874 24549
rect 13938 24485 13966 24549
rect 14030 24485 14940 24549
rect 12409 24469 14940 24485
rect 12409 24405 13506 24469
rect 13570 24405 13598 24469
rect 13662 24405 13690 24469
rect 13754 24405 13782 24469
rect 13846 24405 13874 24469
rect 13938 24405 13966 24469
rect 14030 24405 14940 24469
rect 12409 24389 14940 24405
rect 12409 24325 13506 24389
rect 13570 24325 13598 24389
rect 13662 24325 13690 24389
rect 13754 24325 13782 24389
rect 13846 24325 13874 24389
rect 13938 24325 13966 24389
rect 14030 24325 14940 24389
rect 12409 24309 14940 24325
rect 12409 24245 13506 24309
rect 13570 24245 13598 24309
rect 13662 24245 13690 24309
rect 13754 24245 13782 24309
rect 13846 24245 13874 24309
rect 13938 24245 13966 24309
rect 14030 24245 14940 24309
rect 12409 24229 14940 24245
rect 12409 24165 13506 24229
rect 13570 24165 13598 24229
rect 13662 24165 13690 24229
rect 13754 24165 13782 24229
rect 13846 24165 13874 24229
rect 13938 24165 13966 24229
rect 14030 24165 14940 24229
rect 12409 24148 14940 24165
rect 12409 24084 13506 24148
rect 13570 24084 13598 24148
rect 13662 24084 13690 24148
rect 13754 24084 13782 24148
rect 13846 24084 13874 24148
rect 13938 24084 13966 24148
rect 14030 24084 14940 24148
rect 12409 24067 14940 24084
rect 12409 24003 13506 24067
rect 13570 24003 13598 24067
rect 13662 24003 13690 24067
rect 13754 24003 13782 24067
rect 13846 24003 13874 24067
rect 13938 24003 13966 24067
rect 14030 24003 14940 24067
rect 12409 23986 14940 24003
rect 12409 23922 13506 23986
rect 13570 23922 13598 23986
rect 13662 23922 13690 23986
rect 13754 23922 13782 23986
rect 13846 23922 13874 23986
rect 13938 23922 13966 23986
rect 14030 23922 14940 23986
rect 12409 23905 14940 23922
rect 12409 23841 13506 23905
rect 13570 23841 13598 23905
rect 13662 23841 13690 23905
rect 13754 23841 13782 23905
rect 13846 23841 13874 23905
rect 13938 23841 13966 23905
rect 14030 23841 14940 23905
rect 12409 23824 14940 23841
rect 12409 23760 13506 23824
rect 13570 23760 13598 23824
rect 13662 23760 13690 23824
rect 13754 23760 13782 23824
rect 13846 23760 13874 23824
rect 13938 23760 13966 23824
rect 14030 23760 14940 23824
rect 12409 23743 14940 23760
rect 12409 23679 13506 23743
rect 13570 23679 13598 23743
rect 13662 23679 13690 23743
rect 13754 23679 13782 23743
rect 13846 23679 13874 23743
rect 13938 23679 13966 23743
rect 14030 23679 14940 23743
rect 12409 23662 14940 23679
rect 12409 23598 13506 23662
rect 13570 23598 13598 23662
rect 13662 23598 13690 23662
rect 13754 23598 13782 23662
rect 13846 23598 13874 23662
rect 13938 23598 13966 23662
rect 14030 23598 14940 23662
rect 12409 23581 14940 23598
rect 12409 23517 13506 23581
rect 13570 23517 13598 23581
rect 13662 23517 13690 23581
rect 13754 23517 13782 23581
rect 13846 23517 13874 23581
rect 13938 23517 13966 23581
rect 14030 23517 14940 23581
rect 12409 23500 14940 23517
rect 12409 23436 13506 23500
rect 13570 23436 13598 23500
rect 13662 23436 13690 23500
rect 13754 23436 13782 23500
rect 13846 23436 13874 23500
rect 13938 23436 13966 23500
rect 14030 23436 14940 23500
rect 12409 23419 14940 23436
rect 12409 23355 13506 23419
rect 13570 23355 13598 23419
rect 13662 23355 13690 23419
rect 13754 23355 13782 23419
rect 13846 23355 13874 23419
rect 13938 23355 13966 23419
rect 14030 23355 14940 23419
rect 12409 23338 14940 23355
rect 12409 23274 13506 23338
rect 13570 23274 13598 23338
rect 13662 23274 13690 23338
rect 13754 23274 13782 23338
rect 13846 23274 13874 23338
rect 13938 23274 13966 23338
rect 14030 23274 14940 23338
rect 12409 23257 14940 23274
rect 12409 23193 13506 23257
rect 13570 23193 13598 23257
rect 13662 23193 13690 23257
rect 13754 23193 13782 23257
rect 13846 23193 13874 23257
rect 13938 23193 13966 23257
rect 14030 23193 14940 23257
rect 12409 23176 14940 23193
rect 12409 23112 13506 23176
rect 13570 23112 13598 23176
rect 13662 23112 13690 23176
rect 13754 23112 13782 23176
rect 13846 23112 13874 23176
rect 13938 23112 13966 23176
rect 14030 23112 14940 23176
rect 12409 23095 14940 23112
rect 12409 23031 13506 23095
rect 13570 23031 13598 23095
rect 13662 23031 13690 23095
rect 13754 23031 13782 23095
rect 13846 23031 13874 23095
rect 13938 23031 13966 23095
rect 14030 23031 14940 23095
rect 12409 23014 14940 23031
rect 12409 22950 13506 23014
rect 13570 22950 13598 23014
rect 13662 22950 13690 23014
rect 13754 22950 13782 23014
rect 13846 22950 13874 23014
rect 13938 22950 13966 23014
rect 14030 22950 14940 23014
rect 12409 22933 14940 22950
rect 12409 22869 13506 22933
rect 13570 22869 13598 22933
rect 13662 22869 13690 22933
rect 13754 22869 13782 22933
rect 13846 22869 13874 22933
rect 13938 22869 13966 22933
rect 14030 22869 14940 22933
rect 12409 22852 14940 22869
rect 12409 22788 13506 22852
rect 13570 22788 13598 22852
rect 13662 22788 13690 22852
rect 13754 22788 13782 22852
rect 13846 22788 13874 22852
rect 13938 22788 13966 22852
rect 14030 22788 14940 22852
rect 12409 22771 14940 22788
rect 12409 22707 13506 22771
rect 13570 22707 13598 22771
rect 13662 22707 13690 22771
rect 13754 22707 13782 22771
rect 13846 22707 13874 22771
rect 13938 22707 13966 22771
rect 14030 22707 14940 22771
rect 12409 22690 14940 22707
rect 12409 22626 13506 22690
rect 13570 22626 13598 22690
rect 13662 22626 13690 22690
rect 13754 22626 13782 22690
rect 13846 22626 13874 22690
rect 13938 22626 13966 22690
rect 14030 22626 14940 22690
rect 12409 22609 14940 22626
rect 12409 22545 13506 22609
rect 13570 22545 13598 22609
rect 13662 22545 13690 22609
rect 13754 22545 13782 22609
rect 13846 22545 13874 22609
rect 13938 22545 13966 22609
rect 14030 22545 14940 22609
rect 12409 22528 14940 22545
rect 12409 22464 13506 22528
rect 13570 22464 13598 22528
rect 13662 22464 13690 22528
rect 13754 22464 13782 22528
rect 13846 22464 13874 22528
rect 13938 22464 13966 22528
rect 14030 22464 14940 22528
rect 12409 22447 14940 22464
rect 12409 22383 13506 22447
rect 13570 22383 13598 22447
rect 13662 22383 13690 22447
rect 13754 22383 13782 22447
rect 13846 22383 13874 22447
rect 13938 22383 13966 22447
rect 14030 22383 14940 22447
rect 12409 22366 14940 22383
rect 12409 22302 13506 22366
rect 13570 22302 13598 22366
rect 13662 22302 13690 22366
rect 13754 22302 13782 22366
rect 13846 22302 13874 22366
rect 13938 22302 13966 22366
rect 14030 22302 14940 22366
rect 12409 22285 14940 22302
rect 12409 22221 13506 22285
rect 13570 22221 13598 22285
rect 13662 22221 13690 22285
rect 13754 22221 13782 22285
rect 13846 22221 13874 22285
rect 13938 22221 13966 22285
rect 14030 22221 14940 22285
rect 12409 22204 14940 22221
rect 12409 22140 13506 22204
rect 13570 22140 13598 22204
rect 13662 22140 13690 22204
rect 13754 22140 13782 22204
rect 13846 22140 13874 22204
rect 13938 22140 13966 22204
rect 14030 22140 14940 22204
rect 12409 22123 14940 22140
rect 12409 22059 13506 22123
rect 13570 22059 13598 22123
rect 13662 22059 13690 22123
rect 13754 22059 13782 22123
rect 13846 22059 13874 22123
rect 13938 22059 13966 22123
rect 14030 22059 14940 22123
rect 12409 22042 14940 22059
rect 12409 21978 13506 22042
rect 13570 21978 13598 22042
rect 13662 21978 13690 22042
rect 13754 21978 13782 22042
rect 13846 21978 13874 22042
rect 13938 21978 13966 22042
rect 14030 21978 14940 22042
rect 12409 21961 14940 21978
rect 12409 21897 13506 21961
rect 13570 21897 13598 21961
rect 13662 21897 13690 21961
rect 13754 21897 13782 21961
rect 13846 21897 13874 21961
rect 13938 21897 13966 21961
rect 14030 21897 14940 21961
rect 12409 21880 14940 21897
rect 12409 21816 13506 21880
rect 13570 21816 13598 21880
rect 13662 21816 13690 21880
rect 13754 21816 13782 21880
rect 13846 21816 13874 21880
rect 13938 21816 13966 21880
rect 14030 21816 14940 21880
rect 12409 21799 14940 21816
rect 12409 21735 13506 21799
rect 13570 21735 13598 21799
rect 13662 21735 13690 21799
rect 13754 21735 13782 21799
rect 13846 21735 13874 21799
rect 13938 21735 13966 21799
rect 14030 21735 14940 21799
rect 12409 21718 14940 21735
rect 12409 21654 13506 21718
rect 13570 21654 13598 21718
rect 13662 21654 13690 21718
rect 13754 21654 13782 21718
rect 13846 21654 13874 21718
rect 13938 21654 13966 21718
rect 14030 21654 14940 21718
rect 12409 21637 14940 21654
rect 12409 21573 13506 21637
rect 13570 21573 13598 21637
rect 13662 21573 13690 21637
rect 13754 21573 13782 21637
rect 13846 21573 13874 21637
rect 13938 21573 13966 21637
rect 14030 21573 14940 21637
rect 12409 21556 14940 21573
rect 12409 21492 13506 21556
rect 13570 21492 13598 21556
rect 13662 21492 13690 21556
rect 13754 21492 13782 21556
rect 13846 21492 13874 21556
rect 13938 21492 13966 21556
rect 14030 21492 14940 21556
rect 12409 21475 14940 21492
rect 12409 21411 13506 21475
rect 13570 21411 13598 21475
rect 13662 21411 13690 21475
rect 13754 21411 13782 21475
rect 13846 21411 13874 21475
rect 13938 21411 13966 21475
rect 14030 21411 14940 21475
rect 12409 21394 14940 21411
rect 12409 21330 13506 21394
rect 13570 21330 13598 21394
rect 13662 21330 13690 21394
rect 13754 21330 13782 21394
rect 13846 21330 13874 21394
rect 13938 21330 13966 21394
rect 14030 21330 14940 21394
rect 12409 21313 14940 21330
rect 12409 21249 13506 21313
rect 13570 21249 13598 21313
rect 13662 21249 13690 21313
rect 13754 21249 13782 21313
rect 13846 21249 13874 21313
rect 13938 21249 13966 21313
rect 14030 21249 14940 21313
rect 12409 21232 14940 21249
rect 12409 21168 13506 21232
rect 13570 21168 13598 21232
rect 13662 21168 13690 21232
rect 13754 21168 13782 21232
rect 13846 21168 13874 21232
rect 13938 21168 13966 21232
rect 14030 21168 14940 21232
rect 12409 21151 14940 21168
rect 12409 21087 13506 21151
rect 13570 21087 13598 21151
rect 13662 21087 13690 21151
rect 13754 21087 13782 21151
rect 13846 21087 13874 21151
rect 13938 21087 13966 21151
rect 14030 21087 14940 21151
rect 12409 21070 14940 21087
rect 12409 21006 13506 21070
rect 13570 21006 13598 21070
rect 13662 21006 13690 21070
rect 13754 21006 13782 21070
rect 13846 21006 13874 21070
rect 13938 21006 13966 21070
rect 14030 21006 14940 21070
rect 12409 20989 14940 21006
rect 12409 20925 13506 20989
rect 13570 20925 13598 20989
rect 13662 20925 13690 20989
rect 13754 20925 13782 20989
rect 13846 20925 13874 20989
rect 13938 20925 13966 20989
rect 14030 20925 14940 20989
rect 12409 20908 14940 20925
rect 12409 20844 13506 20908
rect 13570 20844 13598 20908
rect 13662 20844 13690 20908
rect 13754 20844 13782 20908
rect 13846 20844 13874 20908
rect 13938 20844 13966 20908
rect 14030 20844 14940 20908
rect 12409 20827 14940 20844
rect 12409 20763 13506 20827
rect 13570 20763 13598 20827
rect 13662 20763 13690 20827
rect 13754 20763 13782 20827
rect 13846 20763 13874 20827
rect 13938 20763 13966 20827
rect 14030 20763 14940 20827
rect 12409 20746 14940 20763
rect 12409 20682 13506 20746
rect 13570 20682 13598 20746
rect 13662 20682 13690 20746
rect 13754 20682 13782 20746
rect 13846 20682 13874 20746
rect 13938 20682 13966 20746
rect 14030 20682 14940 20746
rect 12409 20665 14940 20682
rect 12409 20601 13506 20665
rect 13570 20601 13598 20665
rect 13662 20601 13690 20665
rect 13754 20601 13782 20665
rect 13846 20601 13874 20665
rect 13938 20601 13966 20665
rect 14030 20601 14940 20665
rect 12409 20534 14940 20601
rect 12409 20470 13405 20534
rect 13469 20470 13497 20534
rect 13561 20470 13589 20534
rect 13653 20470 13681 20534
rect 13745 20470 13773 20534
rect 13837 20470 13865 20534
rect 13929 20470 13957 20534
rect 14021 20470 14940 20534
rect 12409 20431 14940 20470
rect 12409 20367 13324 20431
rect 13388 20367 13405 20431
rect 13469 20367 13487 20431
rect 13551 20367 13569 20431
rect 13633 20367 13651 20431
rect 13715 20367 13733 20431
rect 13797 20415 14940 20431
rect 13797 20367 13859 20415
rect 12409 20351 13859 20367
rect 13923 20351 14940 20415
rect 12409 20311 14940 20351
rect 12409 20247 13182 20311
rect 13246 20283 14940 20311
rect 13246 20247 13324 20283
rect 12409 20219 13324 20247
rect 13388 20219 13405 20283
rect 13469 20219 13487 20283
rect 13551 20219 13569 20283
rect 13633 20219 13651 20283
rect 13715 20219 13733 20283
rect 13797 20219 14940 20283
rect 12409 20203 14940 20219
rect 12409 20139 13068 20203
rect 13132 20139 13149 20203
rect 13213 20139 13231 20203
rect 13295 20139 13313 20203
rect 13377 20139 13395 20203
rect 13459 20139 13477 20203
rect 13541 20192 14940 20203
rect 13541 20139 13636 20192
rect 12409 20128 13636 20139
rect 13700 20128 14940 20192
rect 12409 20072 14940 20128
rect 12409 20008 12943 20072
rect 13007 20055 14940 20072
rect 13007 20008 13068 20055
rect 12409 19991 13068 20008
rect 13132 19991 13149 20055
rect 13213 19991 13231 20055
rect 13295 19991 13313 20055
rect 13377 19991 13395 20055
rect 13459 19991 13477 20055
rect 13541 19991 14940 20055
rect 12409 19975 14940 19991
rect 12409 19911 12870 19975
rect 12934 19911 12951 19975
rect 13015 19911 13033 19975
rect 13097 19911 13115 19975
rect 13179 19911 13197 19975
rect 13261 19911 13279 19975
rect 13343 19953 14940 19975
rect 13343 19911 13397 19953
rect 12409 19889 13397 19911
rect 13461 19889 14940 19953
rect 12409 19857 14940 19889
rect 12409 19793 12728 19857
rect 12792 19827 14940 19857
rect 12792 19793 12870 19827
rect 12409 19763 12870 19793
rect 12934 19763 12951 19827
rect 13015 19763 13033 19827
rect 13097 19763 13115 19827
rect 13179 19763 13197 19827
rect 13261 19763 13279 19827
rect 13343 19763 14940 19827
rect 12409 19742 14940 19763
rect 12409 19678 12646 19742
rect 12710 19678 12727 19742
rect 12791 19678 12809 19742
rect 12873 19678 12891 19742
rect 12955 19678 12973 19742
rect 13037 19678 13055 19742
rect 13119 19738 14940 19742
rect 13119 19678 13182 19738
rect 12409 19674 13182 19678
rect 13246 19674 14940 19738
rect 12409 19658 14940 19674
rect 12409 19594 12446 19658
rect 12510 19594 12554 19658
rect 12618 19594 14940 19658
rect 12409 19549 12646 19594
rect 12409 19485 12446 19549
rect 12510 19485 12554 19549
rect 12618 19530 12646 19549
rect 12710 19530 12727 19594
rect 12791 19530 12809 19594
rect 12873 19530 12891 19594
rect 12955 19530 12973 19594
rect 13037 19530 13055 19594
rect 13119 19530 14940 19594
rect 12618 19508 14940 19530
rect 12618 19485 12646 19508
rect 12409 19444 12646 19485
rect 12710 19444 12737 19508
rect 12801 19444 12828 19508
rect 12892 19499 14940 19508
rect 12892 19444 12950 19499
rect 12409 19440 12950 19444
rect 12409 19376 12446 19440
rect 12510 19376 12554 19440
rect 12618 19435 12950 19440
rect 13014 19435 14940 19499
rect 12618 19376 14940 19435
rect 3121 18862 4779 18900
tri 3121 18852 3131 18862 ne
rect 3131 18852 4779 18862
tri 4779 18852 4827 18900 sw
tri 5207 18852 5255 18900 ne
rect 5255 18852 6407 18900
tri 8336 18852 8567 19083 se
rect 8567 18934 9339 19362
tri 9339 18934 9767 19362 nw
tri 9984 19151 10195 19362 se
rect 10195 19151 11680 19362
tri 11680 19151 11891 19362 nw
rect 12409 19360 14940 19376
rect 12409 19332 12646 19360
rect 12409 19268 12446 19332
rect 12510 19268 12554 19332
rect 12618 19296 12646 19332
rect 12710 19296 12737 19360
rect 12801 19296 12828 19360
rect 12892 19296 14940 19360
rect 12618 19268 14940 19296
rect 12409 19224 14940 19268
rect 12409 19160 12446 19224
rect 12510 19160 12554 19224
rect 12618 19160 14940 19224
rect 12409 19151 14940 19160
tri 9767 18934 9984 19151 se
rect 9984 18934 10951 19151
rect 8567 18852 9257 18934
tri 9257 18852 9339 18934 nw
tri 9685 18852 9767 18934 se
rect 9767 18852 10951 18934
tri 2580 18472 2960 18852 sw
tri 3131 18472 3511 18852 ne
rect 3511 18678 4827 18852
tri 4827 18678 5001 18852 sw
tri 5255 18678 5429 18852 ne
rect 5429 18678 6407 18852
tri 8162 18678 8336 18852 se
rect 8336 18838 9243 18852
tri 9243 18838 9257 18852 nw
tri 9671 18838 9685 18852 se
rect 9685 18838 10951 18852
rect 8336 18678 8815 18838
rect 3511 18472 5001 18678
tri 5001 18472 5207 18678 sw
tri 5429 18472 5635 18678 ne
rect 5635 18472 6407 18678
rect 100 18311 2960 18472
tri 2960 18311 3121 18472 sw
tri 3511 18311 3672 18472 ne
rect 3672 18311 5207 18472
rect 100 18213 3121 18311
tri 3121 18213 3219 18311 sw
tri 3672 18213 3770 18311 ne
rect 3770 18213 5207 18311
rect 100 17662 3219 18213
tri 3219 17662 3770 18213 sw
tri 3770 17662 4321 18213 ne
rect 4321 18075 5207 18213
tri 5207 18075 5604 18472 sw
tri 5635 18075 6032 18472 ne
rect 6032 18410 6407 18472
tri 6407 18410 6675 18678 sw
tri 7894 18410 8162 18678 se
rect 8162 18410 8815 18678
tri 8815 18410 9243 18838 nw
tri 9243 18410 9671 18838 se
rect 9671 18422 10951 18838
tri 10951 18422 11680 19151 nw
rect 9671 18410 10933 18422
rect 6032 18075 6675 18410
tri 6675 18075 7010 18410 sw
tri 7559 18075 7894 18410 se
rect 7894 18075 8387 18410
rect 4321 17700 5604 18075
tri 5604 17700 5979 18075 sw
tri 6032 17700 6407 18075 ne
rect 6407 17982 8387 18075
tri 8387 17982 8815 18410 nw
tri 8815 17982 9243 18410 se
rect 9243 18404 10933 18410
tri 10933 18404 10951 18422 nw
tri 11662 18404 11680 18422 se
rect 11680 18404 14940 19151
rect 9243 17982 10204 18404
rect 6407 17917 8322 17982
tri 8322 17917 8387 17982 nw
tri 8750 17917 8815 17982 se
rect 8815 17917 10204 17982
rect 6407 17700 7894 17917
rect 4321 17662 5979 17700
rect 100 17213 3770 17662
tri 3770 17213 4219 17662 sw
tri 4321 17272 4711 17662 ne
rect 4711 17489 5979 17662
tri 5979 17489 6190 17700 sw
tri 6407 17489 6618 17700 ne
rect 6618 17489 7894 17700
tri 7894 17489 8322 17917 nw
tri 8322 17489 8750 17917 se
rect 8750 17489 10204 17917
tri 10204 17675 10933 18404 nw
rect 10933 17675 14940 18404
rect 4711 17472 6190 17489
tri 6190 17472 6207 17489 sw
tri 6618 17472 6635 17489 ne
rect 6635 17472 7877 17489
tri 7877 17472 7894 17489 nw
rect 4711 17272 6207 17472
tri 6207 17272 6407 17472 sw
tri 6635 17272 6835 17472 ne
rect 6835 17272 7877 17472
tri 4711 17250 4733 17272 ne
rect 4733 17250 6407 17272
tri 6407 17250 6429 17272 sw
tri 4733 17213 4770 17250 ne
rect 100 16930 4219 17213
tri 4219 16930 4502 17213 sw
rect 4770 16930 6429 17250
tri 6835 17206 6901 17272 ne
rect 100 16662 4502 16930
tri 4502 16662 4770 16930 sw
tri 4770 16796 4904 16930 ne
rect 4904 16796 6429 16930
tri 6429 16796 6571 16938 sw
tri 6759 16796 6901 16938 se
rect 6901 16796 7877 17272
rect 8322 17392 10204 17489
rect 8322 17339 10151 17392
tri 10151 17339 10204 17392 nw
rect 8322 17206 10018 17339
tri 10018 17206 10151 17339 nw
tri 7877 16796 8019 16938 sw
tri 8180 16796 8322 16938 se
rect 8322 16796 9774 17206
tri 9774 16962 10018 17206 nw
rect 10220 16962 14940 17675
tri 4904 16662 5038 16796 ne
rect 5038 16662 9774 16796
rect 100 16532 4770 16662
tri 4770 16532 4900 16662 sw
rect 100 0 4900 16532
tri 5038 16500 5200 16662 ne
rect 5200 15363 9774 16662
rect 5200 14948 9359 15363
tri 9359 14948 9774 15363 nw
rect 5008 8286 5074 8293
rect 5072 8222 5074 8286
rect 5008 8198 5074 8222
rect 5072 8134 5074 8198
rect 5008 8110 5074 8134
rect 5072 8046 5074 8110
rect 5008 8022 5074 8046
rect 5072 7958 5074 8022
rect 5008 5201 5074 7958
rect 5008 5145 5013 5201
rect 5069 5145 5074 5201
rect 5008 5121 5074 5145
rect 5008 5065 5013 5121
rect 5069 5065 5074 5121
rect 5008 5054 5074 5065
rect 5008 4867 5092 4877
rect 5008 4811 5022 4867
rect 5078 4811 5092 4867
rect 5008 4785 5092 4811
rect 5008 4729 5022 4785
rect 5078 4729 5092 4785
rect 5008 4702 5092 4729
rect 5008 4646 5022 4702
rect 5078 4646 5092 4702
rect 5008 4449 5092 4646
rect 5008 4385 5018 4449
rect 5082 4385 5092 4449
rect 5008 4366 5092 4385
rect 5008 4302 5018 4366
rect 5082 4302 5092 4366
rect 5008 4284 5092 4302
rect 5008 4220 5018 4284
rect 5082 4220 5092 4284
rect 5008 4202 5092 4220
rect 5008 4138 5018 4202
rect 5082 4138 5092 4202
rect 5008 4120 5092 4138
rect 5008 4056 5018 4120
rect 5082 4056 5092 4120
rect 5008 4038 5092 4056
rect 5008 3974 5018 4038
rect 5082 3974 5092 4038
rect 5008 3956 5092 3974
rect 5008 3892 5018 3956
rect 5082 3892 5092 3956
rect 5008 3874 5092 3892
rect 5008 3810 5018 3874
rect 5082 3810 5092 3874
rect 5008 3792 5092 3810
rect 5008 3728 5018 3792
rect 5082 3728 5092 3792
rect 5008 3710 5092 3728
rect 5008 3646 5018 3710
rect 5082 3646 5092 3710
rect 5008 3628 5092 3646
rect 5008 3564 5018 3628
rect 5082 3564 5092 3628
rect 5008 3558 5092 3564
rect 5200 4220 7376 14948
tri 7376 14221 8103 14948 nw
rect 5200 4164 5212 4220
rect 5268 4164 5347 4220
rect 5403 4164 5481 4220
rect 5537 4164 5615 4220
rect 5671 4164 5749 4220
rect 5805 4164 5883 4220
rect 5939 4164 7376 4220
rect 5200 4100 7376 4164
rect 5200 4044 5212 4100
rect 5268 4044 5347 4100
rect 5403 4044 5481 4100
rect 5537 4044 5615 4100
rect 5671 4044 5749 4100
rect 5805 4044 5883 4100
rect 5939 4044 7376 4100
rect 5200 0 7376 4044
rect 7676 13877 9851 13898
rect 7676 13821 7691 13877
rect 7747 13821 7775 13877
rect 7831 13821 7858 13877
rect 7914 13821 7941 13877
rect 7997 13821 8024 13877
rect 8080 13821 8107 13877
rect 8163 13821 8190 13877
rect 8246 13821 8273 13877
rect 8329 13821 8356 13877
rect 8412 13821 8439 13877
rect 8495 13821 8522 13877
rect 8578 13821 8605 13877
rect 8661 13821 8688 13877
rect 8744 13821 8771 13877
rect 8827 13821 8854 13877
rect 8910 13821 8937 13877
rect 8993 13821 9020 13877
rect 9076 13821 9103 13877
rect 9159 13821 9186 13877
rect 9242 13821 9269 13877
rect 9325 13821 9352 13877
rect 9408 13821 9435 13877
rect 9491 13821 9518 13877
rect 9574 13821 9601 13877
rect 9657 13821 9684 13877
rect 9740 13821 9767 13877
rect 9823 13821 9851 13877
rect 7676 13789 9851 13821
rect 7676 13733 7691 13789
rect 7747 13733 7775 13789
rect 7831 13733 7858 13789
rect 7914 13733 7941 13789
rect 7997 13733 8024 13789
rect 8080 13733 8107 13789
rect 8163 13733 8190 13789
rect 8246 13733 8273 13789
rect 8329 13733 8356 13789
rect 8412 13733 8439 13789
rect 8495 13733 8522 13789
rect 8578 13733 8605 13789
rect 8661 13733 8688 13789
rect 8744 13733 8771 13789
rect 8827 13733 8854 13789
rect 8910 13733 8937 13789
rect 8993 13733 9020 13789
rect 9076 13733 9103 13789
rect 9159 13733 9186 13789
rect 9242 13733 9269 13789
rect 9325 13733 9352 13789
rect 9408 13733 9435 13789
rect 9491 13733 9518 13789
rect 9574 13733 9601 13789
rect 9657 13733 9684 13789
rect 9740 13733 9767 13789
rect 9823 13733 9851 13789
rect 7676 13701 9851 13733
rect 7676 13645 7691 13701
rect 7747 13645 7775 13701
rect 7831 13645 7858 13701
rect 7914 13645 7941 13701
rect 7997 13645 8024 13701
rect 8080 13645 8107 13701
rect 8163 13645 8190 13701
rect 8246 13645 8273 13701
rect 8329 13645 8356 13701
rect 8412 13645 8439 13701
rect 8495 13645 8522 13701
rect 8578 13645 8605 13701
rect 8661 13645 8688 13701
rect 8744 13645 8771 13701
rect 8827 13645 8854 13701
rect 8910 13645 8937 13701
rect 8993 13645 9020 13701
rect 9076 13645 9103 13701
rect 9159 13645 9186 13701
rect 9242 13645 9269 13701
rect 9325 13645 9352 13701
rect 9408 13645 9435 13701
rect 9491 13645 9518 13701
rect 9574 13645 9601 13701
rect 9657 13645 9684 13701
rect 9740 13645 9767 13701
rect 9823 13645 9851 13701
rect 7676 13613 9851 13645
rect 7676 13557 7691 13613
rect 7747 13557 7775 13613
rect 7831 13557 7858 13613
rect 7914 13557 7941 13613
rect 7997 13557 8024 13613
rect 8080 13557 8107 13613
rect 8163 13557 8190 13613
rect 8246 13557 8273 13613
rect 8329 13557 8356 13613
rect 8412 13557 8439 13613
rect 8495 13557 8522 13613
rect 8578 13557 8605 13613
rect 8661 13557 8688 13613
rect 8744 13557 8771 13613
rect 8827 13557 8854 13613
rect 8910 13557 8937 13613
rect 8993 13557 9020 13613
rect 9076 13557 9103 13613
rect 9159 13557 9186 13613
rect 9242 13557 9269 13613
rect 9325 13557 9352 13613
rect 9408 13557 9435 13613
rect 9491 13557 9518 13613
rect 9574 13557 9601 13613
rect 9657 13557 9684 13613
rect 9740 13557 9767 13613
rect 9823 13557 9851 13613
rect 7676 13525 9851 13557
rect 7676 13469 7691 13525
rect 7747 13469 7775 13525
rect 7831 13469 7858 13525
rect 7914 13469 7941 13525
rect 7997 13469 8024 13525
rect 8080 13469 8107 13525
rect 8163 13469 8190 13525
rect 8246 13469 8273 13525
rect 8329 13469 8356 13525
rect 8412 13469 8439 13525
rect 8495 13469 8522 13525
rect 8578 13469 8605 13525
rect 8661 13469 8688 13525
rect 8744 13469 8771 13525
rect 8827 13469 8854 13525
rect 8910 13469 8937 13525
rect 8993 13469 9020 13525
rect 9076 13469 9103 13525
rect 9159 13469 9186 13525
rect 9242 13469 9269 13525
rect 9325 13469 9352 13525
rect 9408 13469 9435 13525
rect 9491 13469 9518 13525
rect 9574 13469 9601 13525
rect 9657 13469 9684 13525
rect 9740 13469 9767 13525
rect 9823 13469 9851 13525
rect 7676 13437 9851 13469
rect 7676 13381 7691 13437
rect 7747 13381 7775 13437
rect 7831 13381 7858 13437
rect 7914 13381 7941 13437
rect 7997 13381 8024 13437
rect 8080 13381 8107 13437
rect 8163 13381 8190 13437
rect 8246 13381 8273 13437
rect 8329 13381 8356 13437
rect 8412 13381 8439 13437
rect 8495 13381 8522 13437
rect 8578 13381 8605 13437
rect 8661 13381 8688 13437
rect 8744 13381 8771 13437
rect 8827 13381 8854 13437
rect 8910 13381 8937 13437
rect 8993 13381 9020 13437
rect 9076 13381 9103 13437
rect 9159 13381 9186 13437
rect 9242 13381 9269 13437
rect 9325 13381 9352 13437
rect 9408 13381 9435 13437
rect 9491 13381 9518 13437
rect 9574 13381 9601 13437
rect 9657 13381 9684 13437
rect 9740 13381 9767 13437
rect 9823 13381 9851 13437
rect 7676 11882 9851 13381
rect 7676 11826 7691 11882
rect 7747 11826 7775 11882
rect 7831 11826 7858 11882
rect 7914 11826 7941 11882
rect 7997 11826 8024 11882
rect 8080 11826 8107 11882
rect 8163 11826 8190 11882
rect 8246 11826 8273 11882
rect 8329 11826 8356 11882
rect 8412 11826 8439 11882
rect 8495 11826 8522 11882
rect 8578 11826 8605 11882
rect 8661 11826 8688 11882
rect 8744 11826 8771 11882
rect 8827 11826 8854 11882
rect 8910 11826 8937 11882
rect 8993 11826 9020 11882
rect 9076 11826 9103 11882
rect 9159 11826 9186 11882
rect 9242 11826 9269 11882
rect 9325 11826 9352 11882
rect 9408 11826 9435 11882
rect 9491 11826 9518 11882
rect 9574 11826 9601 11882
rect 9657 11826 9684 11882
rect 9740 11826 9767 11882
rect 9823 11826 9851 11882
rect 7676 11794 9851 11826
rect 7676 11738 7691 11794
rect 7747 11738 7775 11794
rect 7831 11738 7858 11794
rect 7914 11738 7941 11794
rect 7997 11738 8024 11794
rect 8080 11738 8107 11794
rect 8163 11738 8190 11794
rect 8246 11738 8273 11794
rect 8329 11738 8356 11794
rect 8412 11738 8439 11794
rect 8495 11738 8522 11794
rect 8578 11738 8605 11794
rect 8661 11738 8688 11794
rect 8744 11738 8771 11794
rect 8827 11738 8854 11794
rect 8910 11738 8937 11794
rect 8993 11738 9020 11794
rect 9076 11738 9103 11794
rect 9159 11738 9186 11794
rect 9242 11738 9269 11794
rect 9325 11738 9352 11794
rect 9408 11738 9435 11794
rect 9491 11738 9518 11794
rect 9574 11738 9601 11794
rect 9657 11738 9684 11794
rect 9740 11738 9767 11794
rect 9823 11738 9851 11794
rect 7676 11706 9851 11738
rect 7676 11650 7691 11706
rect 7747 11650 7775 11706
rect 7831 11650 7858 11706
rect 7914 11650 7941 11706
rect 7997 11650 8024 11706
rect 8080 11650 8107 11706
rect 8163 11650 8190 11706
rect 8246 11650 8273 11706
rect 8329 11650 8356 11706
rect 8412 11650 8439 11706
rect 8495 11650 8522 11706
rect 8578 11650 8605 11706
rect 8661 11650 8688 11706
rect 8744 11650 8771 11706
rect 8827 11650 8854 11706
rect 8910 11650 8937 11706
rect 8993 11650 9020 11706
rect 9076 11650 9103 11706
rect 9159 11650 9186 11706
rect 9242 11650 9269 11706
rect 9325 11650 9352 11706
rect 9408 11650 9435 11706
rect 9491 11650 9518 11706
rect 9574 11650 9601 11706
rect 9657 11650 9684 11706
rect 9740 11650 9767 11706
rect 9823 11650 9851 11706
rect 7676 11618 9851 11650
rect 7676 11562 7691 11618
rect 7747 11562 7775 11618
rect 7831 11562 7858 11618
rect 7914 11562 7941 11618
rect 7997 11562 8024 11618
rect 8080 11562 8107 11618
rect 8163 11562 8190 11618
rect 8246 11562 8273 11618
rect 8329 11562 8356 11618
rect 8412 11562 8439 11618
rect 8495 11562 8522 11618
rect 8578 11562 8605 11618
rect 8661 11562 8688 11618
rect 8744 11562 8771 11618
rect 8827 11562 8854 11618
rect 8910 11562 8937 11618
rect 8993 11562 9020 11618
rect 9076 11562 9103 11618
rect 9159 11562 9186 11618
rect 9242 11562 9269 11618
rect 9325 11562 9352 11618
rect 9408 11562 9435 11618
rect 9491 11562 9518 11618
rect 9574 11562 9601 11618
rect 9657 11562 9684 11618
rect 9740 11562 9767 11618
rect 9823 11562 9851 11618
rect 7676 11530 9851 11562
rect 7676 11474 7691 11530
rect 7747 11474 7775 11530
rect 7831 11474 7858 11530
rect 7914 11474 7941 11530
rect 7997 11474 8024 11530
rect 8080 11474 8107 11530
rect 8163 11474 8190 11530
rect 8246 11474 8273 11530
rect 8329 11474 8356 11530
rect 8412 11474 8439 11530
rect 8495 11474 8522 11530
rect 8578 11474 8605 11530
rect 8661 11474 8688 11530
rect 8744 11474 8771 11530
rect 8827 11474 8854 11530
rect 8910 11474 8937 11530
rect 8993 11474 9020 11530
rect 9076 11474 9103 11530
rect 9159 11474 9186 11530
rect 9242 11474 9269 11530
rect 9325 11474 9352 11530
rect 9408 11474 9435 11530
rect 9491 11474 9518 11530
rect 9574 11474 9601 11530
rect 9657 11474 9684 11530
rect 9740 11474 9767 11530
rect 9823 11474 9851 11530
rect 7676 11442 9851 11474
rect 7676 11386 7691 11442
rect 7747 11386 7775 11442
rect 7831 11386 7858 11442
rect 7914 11386 7941 11442
rect 7997 11386 8024 11442
rect 8080 11386 8107 11442
rect 8163 11386 8190 11442
rect 8246 11386 8273 11442
rect 8329 11386 8356 11442
rect 8412 11386 8439 11442
rect 8495 11386 8522 11442
rect 8578 11386 8605 11442
rect 8661 11386 8688 11442
rect 8744 11386 8771 11442
rect 8827 11386 8854 11442
rect 8910 11386 8937 11442
rect 8993 11386 9020 11442
rect 9076 11386 9103 11442
rect 9159 11386 9186 11442
rect 9242 11386 9269 11442
rect 9325 11386 9352 11442
rect 9408 11386 9435 11442
rect 9491 11386 9518 11442
rect 9574 11386 9601 11442
rect 9657 11386 9684 11442
rect 9740 11386 9767 11442
rect 9823 11386 9851 11442
rect 7676 9877 9851 11386
rect 7676 9821 7691 9877
rect 7747 9821 7775 9877
rect 7831 9821 7858 9877
rect 7914 9821 7941 9877
rect 7997 9821 8024 9877
rect 8080 9821 8107 9877
rect 8163 9821 8190 9877
rect 8246 9821 8273 9877
rect 8329 9821 8356 9877
rect 8412 9821 8439 9877
rect 8495 9821 8522 9877
rect 8578 9821 8605 9877
rect 8661 9821 8688 9877
rect 8744 9821 8771 9877
rect 8827 9821 8854 9877
rect 8910 9821 8937 9877
rect 8993 9821 9020 9877
rect 9076 9821 9103 9877
rect 9159 9821 9186 9877
rect 9242 9821 9269 9877
rect 9325 9821 9352 9877
rect 9408 9821 9435 9877
rect 9491 9821 9518 9877
rect 9574 9821 9601 9877
rect 9657 9821 9684 9877
rect 9740 9821 9767 9877
rect 9823 9821 9851 9877
rect 7676 9789 9851 9821
rect 7676 9733 7691 9789
rect 7747 9733 7775 9789
rect 7831 9733 7858 9789
rect 7914 9733 7941 9789
rect 7997 9733 8024 9789
rect 8080 9733 8107 9789
rect 8163 9733 8190 9789
rect 8246 9733 8273 9789
rect 8329 9733 8356 9789
rect 8412 9733 8439 9789
rect 8495 9733 8522 9789
rect 8578 9733 8605 9789
rect 8661 9733 8688 9789
rect 8744 9733 8771 9789
rect 8827 9733 8854 9789
rect 8910 9733 8937 9789
rect 8993 9733 9020 9789
rect 9076 9733 9103 9789
rect 9159 9733 9186 9789
rect 9242 9733 9269 9789
rect 9325 9733 9352 9789
rect 9408 9733 9435 9789
rect 9491 9733 9518 9789
rect 9574 9733 9601 9789
rect 9657 9733 9684 9789
rect 9740 9733 9767 9789
rect 9823 9733 9851 9789
rect 7676 9701 9851 9733
rect 7676 9645 7691 9701
rect 7747 9645 7775 9701
rect 7831 9645 7858 9701
rect 7914 9645 7941 9701
rect 7997 9645 8024 9701
rect 8080 9645 8107 9701
rect 8163 9645 8190 9701
rect 8246 9645 8273 9701
rect 8329 9645 8356 9701
rect 8412 9645 8439 9701
rect 8495 9645 8522 9701
rect 8578 9645 8605 9701
rect 8661 9645 8688 9701
rect 8744 9645 8771 9701
rect 8827 9645 8854 9701
rect 8910 9645 8937 9701
rect 8993 9645 9020 9701
rect 9076 9645 9103 9701
rect 9159 9645 9186 9701
rect 9242 9645 9269 9701
rect 9325 9645 9352 9701
rect 9408 9645 9435 9701
rect 9491 9645 9518 9701
rect 9574 9645 9601 9701
rect 9657 9645 9684 9701
rect 9740 9645 9767 9701
rect 9823 9645 9851 9701
rect 7676 9613 9851 9645
rect 7676 9557 7691 9613
rect 7747 9557 7775 9613
rect 7831 9557 7858 9613
rect 7914 9557 7941 9613
rect 7997 9557 8024 9613
rect 8080 9557 8107 9613
rect 8163 9557 8190 9613
rect 8246 9557 8273 9613
rect 8329 9557 8356 9613
rect 8412 9557 8439 9613
rect 8495 9557 8522 9613
rect 8578 9557 8605 9613
rect 8661 9557 8688 9613
rect 8744 9557 8771 9613
rect 8827 9557 8854 9613
rect 8910 9557 8937 9613
rect 8993 9557 9020 9613
rect 9076 9557 9103 9613
rect 9159 9557 9186 9613
rect 9242 9557 9269 9613
rect 9325 9557 9352 9613
rect 9408 9557 9435 9613
rect 9491 9557 9518 9613
rect 9574 9557 9601 9613
rect 9657 9557 9684 9613
rect 9740 9557 9767 9613
rect 9823 9557 9851 9613
rect 7676 9525 9851 9557
rect 7676 9469 7691 9525
rect 7747 9469 7775 9525
rect 7831 9469 7858 9525
rect 7914 9469 7941 9525
rect 7997 9469 8024 9525
rect 8080 9469 8107 9525
rect 8163 9469 8190 9525
rect 8246 9469 8273 9525
rect 8329 9469 8356 9525
rect 8412 9469 8439 9525
rect 8495 9469 8522 9525
rect 8578 9469 8605 9525
rect 8661 9469 8688 9525
rect 8744 9469 8771 9525
rect 8827 9469 8854 9525
rect 8910 9469 8937 9525
rect 8993 9469 9020 9525
rect 9076 9469 9103 9525
rect 9159 9469 9186 9525
rect 9242 9469 9269 9525
rect 9325 9469 9352 9525
rect 9408 9469 9435 9525
rect 9491 9469 9518 9525
rect 9574 9469 9601 9525
rect 9657 9469 9684 9525
rect 9740 9469 9767 9525
rect 9823 9469 9851 9525
rect 7676 9437 9851 9469
rect 7676 9381 7691 9437
rect 7747 9381 7775 9437
rect 7831 9381 7858 9437
rect 7914 9381 7941 9437
rect 7997 9381 8024 9437
rect 8080 9381 8107 9437
rect 8163 9381 8190 9437
rect 8246 9381 8273 9437
rect 8329 9381 8356 9437
rect 8412 9381 8439 9437
rect 8495 9381 8522 9437
rect 8578 9381 8605 9437
rect 8661 9381 8688 9437
rect 8744 9381 8771 9437
rect 8827 9381 8854 9437
rect 8910 9381 8937 9437
rect 8993 9381 9020 9437
rect 9076 9381 9103 9437
rect 9159 9381 9186 9437
rect 9242 9381 9269 9437
rect 9325 9381 9352 9437
rect 9408 9381 9435 9437
rect 9491 9381 9518 9437
rect 9574 9381 9601 9437
rect 9657 9381 9684 9437
rect 9740 9381 9767 9437
rect 9823 9381 9851 9437
rect 7676 7882 9851 9381
rect 7676 7826 7691 7882
rect 7747 7826 7775 7882
rect 7831 7826 7858 7882
rect 7914 7826 7941 7882
rect 7997 7826 8024 7882
rect 8080 7826 8107 7882
rect 8163 7826 8190 7882
rect 8246 7826 8273 7882
rect 8329 7826 8356 7882
rect 8412 7826 8439 7882
rect 8495 7826 8522 7882
rect 8578 7826 8605 7882
rect 8661 7826 8688 7882
rect 8744 7826 8771 7882
rect 8827 7826 8854 7882
rect 8910 7826 8937 7882
rect 8993 7826 9020 7882
rect 9076 7826 9103 7882
rect 9159 7826 9186 7882
rect 9242 7826 9269 7882
rect 9325 7826 9352 7882
rect 9408 7826 9435 7882
rect 9491 7826 9518 7882
rect 9574 7826 9601 7882
rect 9657 7826 9684 7882
rect 9740 7826 9767 7882
rect 9823 7826 9851 7882
rect 7676 7794 9851 7826
rect 7676 7738 7691 7794
rect 7747 7738 7775 7794
rect 7831 7738 7858 7794
rect 7914 7738 7941 7794
rect 7997 7738 8024 7794
rect 8080 7738 8107 7794
rect 8163 7738 8190 7794
rect 8246 7738 8273 7794
rect 8329 7738 8356 7794
rect 8412 7738 8439 7794
rect 8495 7738 8522 7794
rect 8578 7738 8605 7794
rect 8661 7738 8688 7794
rect 8744 7738 8771 7794
rect 8827 7738 8854 7794
rect 8910 7738 8937 7794
rect 8993 7738 9020 7794
rect 9076 7738 9103 7794
rect 9159 7738 9186 7794
rect 9242 7738 9269 7794
rect 9325 7738 9352 7794
rect 9408 7738 9435 7794
rect 9491 7738 9518 7794
rect 9574 7738 9601 7794
rect 9657 7738 9684 7794
rect 9740 7738 9767 7794
rect 9823 7738 9851 7794
rect 7676 7706 9851 7738
rect 7676 7650 7691 7706
rect 7747 7650 7775 7706
rect 7831 7650 7858 7706
rect 7914 7650 7941 7706
rect 7997 7650 8024 7706
rect 8080 7650 8107 7706
rect 8163 7650 8190 7706
rect 8246 7650 8273 7706
rect 8329 7650 8356 7706
rect 8412 7650 8439 7706
rect 8495 7650 8522 7706
rect 8578 7650 8605 7706
rect 8661 7650 8688 7706
rect 8744 7650 8771 7706
rect 8827 7650 8854 7706
rect 8910 7650 8937 7706
rect 8993 7650 9020 7706
rect 9076 7650 9103 7706
rect 9159 7650 9186 7706
rect 9242 7650 9269 7706
rect 9325 7650 9352 7706
rect 9408 7650 9435 7706
rect 9491 7650 9518 7706
rect 9574 7650 9601 7706
rect 9657 7650 9684 7706
rect 9740 7650 9767 7706
rect 9823 7650 9851 7706
rect 7676 7618 9851 7650
rect 7676 7562 7691 7618
rect 7747 7562 7775 7618
rect 7831 7562 7858 7618
rect 7914 7562 7941 7618
rect 7997 7562 8024 7618
rect 8080 7562 8107 7618
rect 8163 7562 8190 7618
rect 8246 7562 8273 7618
rect 8329 7562 8356 7618
rect 8412 7562 8439 7618
rect 8495 7562 8522 7618
rect 8578 7562 8605 7618
rect 8661 7562 8688 7618
rect 8744 7562 8771 7618
rect 8827 7562 8854 7618
rect 8910 7562 8937 7618
rect 8993 7562 9020 7618
rect 9076 7562 9103 7618
rect 9159 7562 9186 7618
rect 9242 7562 9269 7618
rect 9325 7562 9352 7618
rect 9408 7562 9435 7618
rect 9491 7562 9518 7618
rect 9574 7562 9601 7618
rect 9657 7562 9684 7618
rect 9740 7562 9767 7618
rect 9823 7562 9851 7618
rect 7676 7530 9851 7562
rect 7676 7474 7691 7530
rect 7747 7474 7775 7530
rect 7831 7474 7858 7530
rect 7914 7474 7941 7530
rect 7997 7474 8024 7530
rect 8080 7474 8107 7530
rect 8163 7474 8190 7530
rect 8246 7474 8273 7530
rect 8329 7474 8356 7530
rect 8412 7474 8439 7530
rect 8495 7474 8522 7530
rect 8578 7474 8605 7530
rect 8661 7474 8688 7530
rect 8744 7474 8771 7530
rect 8827 7474 8854 7530
rect 8910 7474 8937 7530
rect 8993 7474 9020 7530
rect 9076 7474 9103 7530
rect 9159 7474 9186 7530
rect 9242 7474 9269 7530
rect 9325 7474 9352 7530
rect 9408 7474 9435 7530
rect 9491 7474 9518 7530
rect 9574 7474 9601 7530
rect 9657 7474 9684 7530
rect 9740 7474 9767 7530
rect 9823 7474 9851 7530
rect 7676 7442 9851 7474
rect 7676 7386 7691 7442
rect 7747 7386 7775 7442
rect 7831 7386 7858 7442
rect 7914 7386 7941 7442
rect 7997 7386 8024 7442
rect 8080 7386 8107 7442
rect 8163 7386 8190 7442
rect 8246 7386 8273 7442
rect 8329 7386 8356 7442
rect 8412 7386 8439 7442
rect 8495 7386 8522 7442
rect 8578 7386 8605 7442
rect 8661 7386 8688 7442
rect 8744 7386 8771 7442
rect 8827 7386 8854 7442
rect 8910 7386 8937 7442
rect 8993 7386 9020 7442
rect 9076 7386 9103 7442
rect 9159 7386 9186 7442
rect 9242 7386 9269 7442
rect 9325 7386 9352 7442
rect 9408 7386 9435 7442
rect 9491 7386 9518 7442
rect 9574 7386 9601 7442
rect 9657 7386 9684 7442
rect 9740 7386 9767 7442
rect 9823 7386 9851 7442
rect 7676 5877 9851 7386
rect 7676 5821 7691 5877
rect 7747 5821 7775 5877
rect 7831 5821 7858 5877
rect 7914 5821 7941 5877
rect 7997 5821 8024 5877
rect 8080 5821 8107 5877
rect 8163 5821 8190 5877
rect 8246 5821 8273 5877
rect 8329 5821 8356 5877
rect 8412 5821 8439 5877
rect 8495 5821 8522 5877
rect 8578 5821 8605 5877
rect 8661 5821 8688 5877
rect 8744 5821 8771 5877
rect 8827 5821 8854 5877
rect 8910 5821 8937 5877
rect 8993 5821 9020 5877
rect 9076 5821 9103 5877
rect 9159 5821 9186 5877
rect 9242 5821 9269 5877
rect 9325 5821 9352 5877
rect 9408 5821 9435 5877
rect 9491 5821 9518 5877
rect 9574 5821 9601 5877
rect 9657 5821 9684 5877
rect 9740 5821 9767 5877
rect 9823 5821 9851 5877
rect 7676 5789 9851 5821
rect 7676 5733 7691 5789
rect 7747 5733 7775 5789
rect 7831 5733 7858 5789
rect 7914 5733 7941 5789
rect 7997 5733 8024 5789
rect 8080 5733 8107 5789
rect 8163 5733 8190 5789
rect 8246 5733 8273 5789
rect 8329 5733 8356 5789
rect 8412 5733 8439 5789
rect 8495 5733 8522 5789
rect 8578 5733 8605 5789
rect 8661 5733 8688 5789
rect 8744 5733 8771 5789
rect 8827 5733 8854 5789
rect 8910 5733 8937 5789
rect 8993 5733 9020 5789
rect 9076 5733 9103 5789
rect 9159 5733 9186 5789
rect 9242 5733 9269 5789
rect 9325 5733 9352 5789
rect 9408 5733 9435 5789
rect 9491 5733 9518 5789
rect 9574 5733 9601 5789
rect 9657 5733 9684 5789
rect 9740 5733 9767 5789
rect 9823 5733 9851 5789
rect 7676 5701 9851 5733
rect 7676 5645 7691 5701
rect 7747 5645 7775 5701
rect 7831 5645 7858 5701
rect 7914 5645 7941 5701
rect 7997 5645 8024 5701
rect 8080 5645 8107 5701
rect 8163 5645 8190 5701
rect 8246 5645 8273 5701
rect 8329 5645 8356 5701
rect 8412 5645 8439 5701
rect 8495 5645 8522 5701
rect 8578 5645 8605 5701
rect 8661 5645 8688 5701
rect 8744 5645 8771 5701
rect 8827 5645 8854 5701
rect 8910 5645 8937 5701
rect 8993 5645 9020 5701
rect 9076 5645 9103 5701
rect 9159 5645 9186 5701
rect 9242 5645 9269 5701
rect 9325 5645 9352 5701
rect 9408 5645 9435 5701
rect 9491 5645 9518 5701
rect 9574 5645 9601 5701
rect 9657 5645 9684 5701
rect 9740 5645 9767 5701
rect 9823 5645 9851 5701
rect 7676 5613 9851 5645
rect 7676 5557 7691 5613
rect 7747 5557 7775 5613
rect 7831 5557 7858 5613
rect 7914 5557 7941 5613
rect 7997 5557 8024 5613
rect 8080 5557 8107 5613
rect 8163 5557 8190 5613
rect 8246 5557 8273 5613
rect 8329 5557 8356 5613
rect 8412 5557 8439 5613
rect 8495 5557 8522 5613
rect 8578 5557 8605 5613
rect 8661 5557 8688 5613
rect 8744 5557 8771 5613
rect 8827 5557 8854 5613
rect 8910 5557 8937 5613
rect 8993 5557 9020 5613
rect 9076 5557 9103 5613
rect 9159 5557 9186 5613
rect 9242 5557 9269 5613
rect 9325 5557 9352 5613
rect 9408 5557 9435 5613
rect 9491 5557 9518 5613
rect 9574 5557 9601 5613
rect 9657 5557 9684 5613
rect 9740 5557 9767 5613
rect 9823 5557 9851 5613
rect 7676 5525 9851 5557
rect 7676 5469 7691 5525
rect 7747 5469 7775 5525
rect 7831 5469 7858 5525
rect 7914 5469 7941 5525
rect 7997 5469 8024 5525
rect 8080 5469 8107 5525
rect 8163 5469 8190 5525
rect 8246 5469 8273 5525
rect 8329 5469 8356 5525
rect 8412 5469 8439 5525
rect 8495 5469 8522 5525
rect 8578 5469 8605 5525
rect 8661 5469 8688 5525
rect 8744 5469 8771 5525
rect 8827 5469 8854 5525
rect 8910 5469 8937 5525
rect 8993 5469 9020 5525
rect 9076 5469 9103 5525
rect 9159 5469 9186 5525
rect 9242 5469 9269 5525
rect 9325 5469 9352 5525
rect 9408 5469 9435 5525
rect 9491 5469 9518 5525
rect 9574 5469 9601 5525
rect 9657 5469 9684 5525
rect 9740 5469 9767 5525
rect 9823 5469 9851 5525
rect 7676 5437 9851 5469
rect 7676 5381 7691 5437
rect 7747 5381 7775 5437
rect 7831 5381 7858 5437
rect 7914 5381 7941 5437
rect 7997 5381 8024 5437
rect 8080 5381 8107 5437
rect 8163 5381 8190 5437
rect 8246 5381 8273 5437
rect 8329 5381 8356 5437
rect 8412 5381 8439 5437
rect 8495 5381 8522 5437
rect 8578 5381 8605 5437
rect 8661 5381 8688 5437
rect 8744 5381 8771 5437
rect 8827 5381 8854 5437
rect 8910 5381 8937 5437
rect 8993 5381 9020 5437
rect 9076 5381 9103 5437
rect 9159 5381 9186 5437
rect 9242 5381 9269 5437
rect 9325 5381 9352 5437
rect 9408 5381 9435 5437
rect 9491 5381 9518 5437
rect 9574 5381 9601 5437
rect 9657 5381 9684 5437
rect 9740 5381 9767 5437
rect 9823 5381 9851 5437
rect 7676 4724 9851 5381
rect 7676 4668 7692 4724
rect 7748 4668 7853 4724
rect 7909 4668 8014 4724
rect 8070 4668 8175 4724
rect 8231 4668 8336 4724
rect 8392 4668 8497 4724
rect 8553 4668 8658 4724
rect 8714 4668 8819 4724
rect 8875 4668 8980 4724
rect 9036 4668 9141 4724
rect 9197 4668 9302 4724
rect 9358 4668 9462 4724
rect 9518 4668 9622 4724
rect 9678 4668 9782 4724
rect 9838 4668 9851 4724
rect 7676 4636 9851 4668
rect 7676 4580 7692 4636
rect 7748 4580 7853 4636
rect 7909 4580 8014 4636
rect 8070 4580 8175 4636
rect 8231 4580 8336 4636
rect 8392 4580 8497 4636
rect 8553 4580 8658 4636
rect 8714 4580 8819 4636
rect 8875 4580 8980 4636
rect 9036 4580 9141 4636
rect 9197 4580 9302 4636
rect 9358 4580 9462 4636
rect 9518 4580 9622 4636
rect 9678 4580 9782 4636
rect 9838 4580 9851 4636
rect 7676 0 9851 4580
rect 10151 0 14940 16962
<< via3 >>
rect 2220 34073 2284 34137
rect 2305 34073 2369 34137
rect 2394 34133 2458 34197
rect 2502 34133 2566 34197
rect 2123 33987 2187 34051
rect 2204 33987 2268 34051
rect 2284 33987 2348 34051
rect 2394 34025 2458 34089
rect 2502 34025 2566 34089
rect 1998 33851 2062 33915
rect 2123 33869 2187 33933
rect 2204 33869 2268 33933
rect 2284 33869 2348 33933
rect 2394 33917 2458 33981
rect 2502 33917 2566 33981
rect 1893 33754 1957 33818
rect 1975 33754 2039 33818
rect 2057 33754 2121 33818
rect 2139 33754 2203 33818
rect 2221 33754 2285 33818
rect 2302 33754 2366 33818
rect 2394 33808 2458 33872
rect 2502 33808 2566 33872
rect 2394 33699 2458 33763
rect 2502 33699 2566 33763
rect 1766 33619 1830 33683
rect 1893 33606 1957 33670
rect 1975 33606 2039 33670
rect 2057 33606 2121 33670
rect 2139 33606 2203 33670
rect 2221 33606 2285 33670
rect 2302 33606 2366 33670
rect 1684 33508 1748 33572
rect 1782 33508 1846 33572
rect 1880 33508 1944 33572
rect 1978 33508 2042 33572
rect 2075 33508 2139 33572
rect 2220 33500 2284 33564
rect 1551 33404 1615 33468
rect 1684 33384 1748 33448
rect 1782 33384 1846 33448
rect 1880 33384 1944 33448
rect 1978 33384 2042 33448
rect 2075 33384 2139 33448
rect 1471 33302 1535 33366
rect 1553 33302 1617 33366
rect 1635 33302 1699 33366
rect 1717 33302 1781 33366
rect 1799 33302 1863 33366
rect 1880 33302 1944 33366
rect 2005 33285 2069 33349
rect 1312 33165 1376 33229
rect 1471 33154 1535 33218
rect 1553 33154 1617 33218
rect 1635 33154 1699 33218
rect 1717 33154 1781 33218
rect 1799 33154 1863 33218
rect 1880 33154 1944 33218
rect 1215 33074 1279 33138
rect 1297 33074 1361 33138
rect 1379 33074 1443 33138
rect 1461 33074 1525 33138
rect 1543 33074 1607 33138
rect 1624 33074 1688 33138
rect 1766 33046 1830 33110
rect 1089 32942 1153 33006
rect 1215 32926 1279 32990
rect 1297 32926 1361 32990
rect 1379 32926 1443 32990
rect 1461 32926 1525 32990
rect 1543 32926 1607 32990
rect 1624 32926 1688 32990
rect 967 32844 1031 32908
rect 1059 32844 1123 32908
rect 1151 32844 1215 32908
rect 1243 32844 1307 32908
rect 1335 32844 1399 32908
rect 1427 32844 1491 32908
rect 967 32764 1031 32828
rect 1059 32764 1123 32828
rect 1151 32764 1215 32828
rect 1243 32764 1307 32828
rect 1335 32764 1399 32828
rect 1427 32764 1491 32828
rect 1543 32823 1607 32887
rect 967 32684 1031 32748
rect 1059 32684 1123 32748
rect 1151 32684 1215 32748
rect 1243 32684 1307 32748
rect 1335 32684 1399 32748
rect 1427 32684 1491 32748
rect 967 32604 1031 32668
rect 1059 32604 1123 32668
rect 1151 32604 1215 32668
rect 1243 32604 1307 32668
rect 1335 32604 1399 32668
rect 1427 32604 1491 32668
rect 967 32524 1031 32588
rect 1059 32524 1123 32588
rect 1151 32524 1215 32588
rect 1243 32524 1307 32588
rect 1335 32524 1399 32588
rect 1427 32524 1491 32588
rect 967 32444 1031 32508
rect 1059 32444 1123 32508
rect 1151 32444 1215 32508
rect 1243 32444 1307 32508
rect 1335 32444 1399 32508
rect 1427 32444 1491 32508
rect 967 32364 1031 32428
rect 1059 32364 1123 32428
rect 1151 32364 1215 32428
rect 1243 32364 1307 32428
rect 1335 32364 1399 32428
rect 1427 32364 1491 32428
rect 967 32284 1031 32348
rect 1059 32284 1123 32348
rect 1151 32284 1215 32348
rect 1243 32284 1307 32348
rect 1335 32284 1399 32348
rect 1427 32284 1491 32348
rect 967 32204 1031 32268
rect 1059 32204 1123 32268
rect 1151 32204 1215 32268
rect 1243 32204 1307 32268
rect 1335 32204 1399 32268
rect 1427 32204 1491 32268
rect 967 32124 1031 32188
rect 1059 32124 1123 32188
rect 1151 32124 1215 32188
rect 1243 32124 1307 32188
rect 1335 32124 1399 32188
rect 1427 32124 1491 32188
rect 967 32044 1031 32108
rect 1059 32044 1123 32108
rect 1151 32044 1215 32108
rect 1243 32044 1307 32108
rect 1335 32044 1399 32108
rect 1427 32044 1491 32108
rect 967 31964 1031 32028
rect 1059 31964 1123 32028
rect 1151 31964 1215 32028
rect 1243 31964 1307 32028
rect 1335 31964 1399 32028
rect 1427 31964 1491 32028
rect 967 31884 1031 31948
rect 1059 31884 1123 31948
rect 1151 31884 1215 31948
rect 1243 31884 1307 31948
rect 1335 31884 1399 31948
rect 1427 31884 1491 31948
rect 967 31804 1031 31868
rect 1059 31804 1123 31868
rect 1151 31804 1215 31868
rect 1243 31804 1307 31868
rect 1335 31804 1399 31868
rect 1427 31804 1491 31868
rect 967 31724 1031 31788
rect 1059 31724 1123 31788
rect 1151 31724 1215 31788
rect 1243 31724 1307 31788
rect 1335 31724 1399 31788
rect 1427 31724 1491 31788
rect 967 31644 1031 31708
rect 1059 31644 1123 31708
rect 1151 31644 1215 31708
rect 1243 31644 1307 31708
rect 1335 31644 1399 31708
rect 1427 31644 1491 31708
rect 967 31564 1031 31628
rect 1059 31564 1123 31628
rect 1151 31564 1215 31628
rect 1243 31564 1307 31628
rect 1335 31564 1399 31628
rect 1427 31564 1491 31628
rect 967 31484 1031 31548
rect 1059 31484 1123 31548
rect 1151 31484 1215 31548
rect 1243 31484 1307 31548
rect 1335 31484 1399 31548
rect 1427 31484 1491 31548
rect 967 31404 1031 31468
rect 1059 31404 1123 31468
rect 1151 31404 1215 31468
rect 1243 31404 1307 31468
rect 1335 31404 1399 31468
rect 1427 31404 1491 31468
rect 967 31324 1031 31388
rect 1059 31324 1123 31388
rect 1151 31324 1215 31388
rect 1243 31324 1307 31388
rect 1335 31324 1399 31388
rect 1427 31324 1491 31388
rect 967 31244 1031 31308
rect 1059 31244 1123 31308
rect 1151 31244 1215 31308
rect 1243 31244 1307 31308
rect 1335 31244 1399 31308
rect 1427 31244 1491 31308
rect 967 31164 1031 31228
rect 1059 31164 1123 31228
rect 1151 31164 1215 31228
rect 1243 31164 1307 31228
rect 1335 31164 1399 31228
rect 1427 31164 1491 31228
rect 967 31084 1031 31148
rect 1059 31084 1123 31148
rect 1151 31084 1215 31148
rect 1243 31084 1307 31148
rect 1335 31084 1399 31148
rect 1427 31084 1491 31148
rect 967 31004 1031 31068
rect 1059 31004 1123 31068
rect 1151 31004 1215 31068
rect 1243 31004 1307 31068
rect 1335 31004 1399 31068
rect 1427 31004 1491 31068
rect 967 30924 1031 30988
rect 1059 30924 1123 30988
rect 1151 30924 1215 30988
rect 1243 30924 1307 30988
rect 1335 30924 1399 30988
rect 1427 30924 1491 30988
rect 967 30844 1031 30908
rect 1059 30844 1123 30908
rect 1151 30844 1215 30908
rect 1243 30844 1307 30908
rect 1335 30844 1399 30908
rect 1427 30844 1491 30908
rect 967 30764 1031 30828
rect 1059 30764 1123 30828
rect 1151 30764 1215 30828
rect 1243 30764 1307 30828
rect 1335 30764 1399 30828
rect 1427 30764 1491 30828
rect 967 30684 1031 30748
rect 1059 30684 1123 30748
rect 1151 30684 1215 30748
rect 1243 30684 1307 30748
rect 1335 30684 1399 30748
rect 1427 30684 1491 30748
rect 967 30604 1031 30668
rect 1059 30604 1123 30668
rect 1151 30604 1215 30668
rect 1243 30604 1307 30668
rect 1335 30604 1399 30668
rect 1427 30604 1491 30668
rect 967 30524 1031 30588
rect 1059 30524 1123 30588
rect 1151 30524 1215 30588
rect 1243 30524 1307 30588
rect 1335 30524 1399 30588
rect 1427 30524 1491 30588
rect 967 30444 1031 30508
rect 1059 30444 1123 30508
rect 1151 30444 1215 30508
rect 1243 30444 1307 30508
rect 1335 30444 1399 30508
rect 1427 30444 1491 30508
rect 967 30364 1031 30428
rect 1059 30364 1123 30428
rect 1151 30364 1215 30428
rect 1243 30364 1307 30428
rect 1335 30364 1399 30428
rect 1427 30364 1491 30428
rect 967 30284 1031 30348
rect 1059 30284 1123 30348
rect 1151 30284 1215 30348
rect 1243 30284 1307 30348
rect 1335 30284 1399 30348
rect 1427 30284 1491 30348
rect 967 30204 1031 30268
rect 1059 30204 1123 30268
rect 1151 30204 1215 30268
rect 1243 30204 1307 30268
rect 1335 30204 1399 30268
rect 1427 30204 1491 30268
rect 967 30124 1031 30188
rect 1059 30124 1123 30188
rect 1151 30124 1215 30188
rect 1243 30124 1307 30188
rect 1335 30124 1399 30188
rect 1427 30124 1491 30188
rect 967 30044 1031 30108
rect 1059 30044 1123 30108
rect 1151 30044 1215 30108
rect 1243 30044 1307 30108
rect 1335 30044 1399 30108
rect 1427 30044 1491 30108
rect 967 29964 1031 30028
rect 1059 29964 1123 30028
rect 1151 29964 1215 30028
rect 1243 29964 1307 30028
rect 1335 29964 1399 30028
rect 1427 29964 1491 30028
rect 967 29884 1031 29948
rect 1059 29884 1123 29948
rect 1151 29884 1215 29948
rect 1243 29884 1307 29948
rect 1335 29884 1399 29948
rect 1427 29884 1491 29948
rect 967 29804 1031 29868
rect 1059 29804 1123 29868
rect 1151 29804 1215 29868
rect 1243 29804 1307 29868
rect 1335 29804 1399 29868
rect 1427 29804 1491 29868
rect 967 29724 1031 29788
rect 1059 29724 1123 29788
rect 1151 29724 1215 29788
rect 1243 29724 1307 29788
rect 1335 29724 1399 29788
rect 1427 29724 1491 29788
rect 967 29644 1031 29708
rect 1059 29644 1123 29708
rect 1151 29644 1215 29708
rect 1243 29644 1307 29708
rect 1335 29644 1399 29708
rect 1427 29644 1491 29708
rect 967 29564 1031 29628
rect 1059 29564 1123 29628
rect 1151 29564 1215 29628
rect 1243 29564 1307 29628
rect 1335 29564 1399 29628
rect 1427 29564 1491 29628
rect 967 29484 1031 29548
rect 1059 29484 1123 29548
rect 1151 29484 1215 29548
rect 1243 29484 1307 29548
rect 1335 29484 1399 29548
rect 1427 29484 1491 29548
rect 967 29404 1031 29468
rect 1059 29404 1123 29468
rect 1151 29404 1215 29468
rect 1243 29404 1307 29468
rect 1335 29404 1399 29468
rect 1427 29404 1491 29468
rect 967 29324 1031 29388
rect 1059 29324 1123 29388
rect 1151 29324 1215 29388
rect 1243 29324 1307 29388
rect 1335 29324 1399 29388
rect 1427 29324 1491 29388
rect 967 29244 1031 29308
rect 1059 29244 1123 29308
rect 1151 29244 1215 29308
rect 1243 29244 1307 29308
rect 1335 29244 1399 29308
rect 1427 29244 1491 29308
rect 967 29164 1031 29228
rect 1059 29164 1123 29228
rect 1151 29164 1215 29228
rect 1243 29164 1307 29228
rect 1335 29164 1399 29228
rect 1427 29164 1491 29228
rect 967 29084 1031 29148
rect 1059 29084 1123 29148
rect 1151 29084 1215 29148
rect 1243 29084 1307 29148
rect 1335 29084 1399 29148
rect 1427 29084 1491 29148
rect 967 29004 1031 29068
rect 1059 29004 1123 29068
rect 1151 29004 1215 29068
rect 1243 29004 1307 29068
rect 1335 29004 1399 29068
rect 1427 29004 1491 29068
rect 967 28924 1031 28988
rect 1059 28924 1123 28988
rect 1151 28924 1215 28988
rect 1243 28924 1307 28988
rect 1335 28924 1399 28988
rect 1427 28924 1491 28988
rect 967 28844 1031 28908
rect 1059 28844 1123 28908
rect 1151 28844 1215 28908
rect 1243 28844 1307 28908
rect 1335 28844 1399 28908
rect 1427 28844 1491 28908
rect 967 28764 1031 28828
rect 1059 28764 1123 28828
rect 1151 28764 1215 28828
rect 1243 28764 1307 28828
rect 1335 28764 1399 28828
rect 1427 28764 1491 28828
rect 967 28684 1031 28748
rect 1059 28684 1123 28748
rect 1151 28684 1215 28748
rect 1243 28684 1307 28748
rect 1335 28684 1399 28748
rect 1427 28684 1491 28748
rect 967 28604 1031 28668
rect 1059 28604 1123 28668
rect 1151 28604 1215 28668
rect 1243 28604 1307 28668
rect 1335 28604 1399 28668
rect 1427 28604 1491 28668
rect 967 28524 1031 28588
rect 1059 28524 1123 28588
rect 1151 28524 1215 28588
rect 1243 28524 1307 28588
rect 1335 28524 1399 28588
rect 1427 28524 1491 28588
rect 967 28444 1031 28508
rect 1059 28444 1123 28508
rect 1151 28444 1215 28508
rect 1243 28444 1307 28508
rect 1335 28444 1399 28508
rect 1427 28444 1491 28508
rect 967 28364 1031 28428
rect 1059 28364 1123 28428
rect 1151 28364 1215 28428
rect 1243 28364 1307 28428
rect 1335 28364 1399 28428
rect 1427 28364 1491 28428
rect 967 28284 1031 28348
rect 1059 28284 1123 28348
rect 1151 28284 1215 28348
rect 1243 28284 1307 28348
rect 1335 28284 1399 28348
rect 1427 28284 1491 28348
rect 967 28204 1031 28268
rect 1059 28204 1123 28268
rect 1151 28204 1215 28268
rect 1243 28204 1307 28268
rect 1335 28204 1399 28268
rect 1427 28204 1491 28268
rect 967 28124 1031 28188
rect 1059 28124 1123 28188
rect 1151 28124 1215 28188
rect 1243 28124 1307 28188
rect 1335 28124 1399 28188
rect 1427 28124 1491 28188
rect 967 28044 1031 28108
rect 1059 28044 1123 28108
rect 1151 28044 1215 28108
rect 1243 28044 1307 28108
rect 1335 28044 1399 28108
rect 1427 28044 1491 28108
rect 967 27964 1031 28028
rect 1059 27964 1123 28028
rect 1151 27964 1215 28028
rect 1243 27964 1307 28028
rect 1335 27964 1399 28028
rect 1427 27964 1491 28028
rect 967 27884 1031 27948
rect 1059 27884 1123 27948
rect 1151 27884 1215 27948
rect 1243 27884 1307 27948
rect 1335 27884 1399 27948
rect 1427 27884 1491 27948
rect 967 27804 1031 27868
rect 1059 27804 1123 27868
rect 1151 27804 1215 27868
rect 1243 27804 1307 27868
rect 1335 27804 1399 27868
rect 1427 27804 1491 27868
rect 967 27724 1031 27788
rect 1059 27724 1123 27788
rect 1151 27724 1215 27788
rect 1243 27724 1307 27788
rect 1335 27724 1399 27788
rect 1427 27724 1491 27788
rect 967 27644 1031 27708
rect 1059 27644 1123 27708
rect 1151 27644 1215 27708
rect 1243 27644 1307 27708
rect 1335 27644 1399 27708
rect 1427 27644 1491 27708
rect 967 27564 1031 27628
rect 1059 27564 1123 27628
rect 1151 27564 1215 27628
rect 1243 27564 1307 27628
rect 1335 27564 1399 27628
rect 1427 27564 1491 27628
rect 967 27484 1031 27548
rect 1059 27484 1123 27548
rect 1151 27484 1215 27548
rect 1243 27484 1307 27548
rect 1335 27484 1399 27548
rect 1427 27484 1491 27548
rect 967 27404 1031 27468
rect 1059 27404 1123 27468
rect 1151 27404 1215 27468
rect 1243 27404 1307 27468
rect 1335 27404 1399 27468
rect 1427 27404 1491 27468
rect 967 27324 1031 27388
rect 1059 27324 1123 27388
rect 1151 27324 1215 27388
rect 1243 27324 1307 27388
rect 1335 27324 1399 27388
rect 1427 27324 1491 27388
rect 967 27244 1031 27308
rect 1059 27244 1123 27308
rect 1151 27244 1215 27308
rect 1243 27244 1307 27308
rect 1335 27244 1399 27308
rect 1427 27244 1491 27308
rect 967 27164 1031 27228
rect 1059 27164 1123 27228
rect 1151 27164 1215 27228
rect 1243 27164 1307 27228
rect 1335 27164 1399 27228
rect 1427 27164 1491 27228
rect 967 27084 1031 27148
rect 1059 27084 1123 27148
rect 1151 27084 1215 27148
rect 1243 27084 1307 27148
rect 1335 27084 1399 27148
rect 1427 27084 1491 27148
rect 967 27004 1031 27068
rect 1059 27004 1123 27068
rect 1151 27004 1215 27068
rect 1243 27004 1307 27068
rect 1335 27004 1399 27068
rect 1427 27004 1491 27068
rect 967 26924 1031 26988
rect 1059 26924 1123 26988
rect 1151 26924 1215 26988
rect 1243 26924 1307 26988
rect 1335 26924 1399 26988
rect 1427 26924 1491 26988
rect 967 26844 1031 26908
rect 1059 26844 1123 26908
rect 1151 26844 1215 26908
rect 1243 26844 1307 26908
rect 1335 26844 1399 26908
rect 1427 26844 1491 26908
rect 967 26764 1031 26828
rect 1059 26764 1123 26828
rect 1151 26764 1215 26828
rect 1243 26764 1307 26828
rect 1335 26764 1399 26828
rect 1427 26764 1491 26828
rect 967 26684 1031 26748
rect 1059 26684 1123 26748
rect 1151 26684 1215 26748
rect 1243 26684 1307 26748
rect 1335 26684 1399 26748
rect 1427 26684 1491 26748
rect 967 26604 1031 26668
rect 1059 26604 1123 26668
rect 1151 26604 1215 26668
rect 1243 26604 1307 26668
rect 1335 26604 1399 26668
rect 1427 26604 1491 26668
rect 967 26524 1031 26588
rect 1059 26524 1123 26588
rect 1151 26524 1215 26588
rect 1243 26524 1307 26588
rect 1335 26524 1399 26588
rect 1427 26524 1491 26588
rect 967 26444 1031 26508
rect 1059 26444 1123 26508
rect 1151 26444 1215 26508
rect 1243 26444 1307 26508
rect 1335 26444 1399 26508
rect 1427 26444 1491 26508
rect 967 26364 1031 26428
rect 1059 26364 1123 26428
rect 1151 26364 1215 26428
rect 1243 26364 1307 26428
rect 1335 26364 1399 26428
rect 1427 26364 1491 26428
rect 967 26284 1031 26348
rect 1059 26284 1123 26348
rect 1151 26284 1215 26348
rect 1243 26284 1307 26348
rect 1335 26284 1399 26348
rect 1427 26284 1491 26348
rect 967 26204 1031 26268
rect 1059 26204 1123 26268
rect 1151 26204 1215 26268
rect 1243 26204 1307 26268
rect 1335 26204 1399 26268
rect 1427 26204 1491 26268
rect 967 26124 1031 26188
rect 1059 26124 1123 26188
rect 1151 26124 1215 26188
rect 1243 26124 1307 26188
rect 1335 26124 1399 26188
rect 1427 26124 1491 26188
rect 967 26044 1031 26108
rect 1059 26044 1123 26108
rect 1151 26044 1215 26108
rect 1243 26044 1307 26108
rect 1335 26044 1399 26108
rect 1427 26044 1491 26108
rect 967 25964 1031 26028
rect 1059 25964 1123 26028
rect 1151 25964 1215 26028
rect 1243 25964 1307 26028
rect 1335 25964 1399 26028
rect 1427 25964 1491 26028
rect 967 25884 1031 25948
rect 1059 25884 1123 25948
rect 1151 25884 1215 25948
rect 1243 25884 1307 25948
rect 1335 25884 1399 25948
rect 1427 25884 1491 25948
rect 967 25804 1031 25868
rect 1059 25804 1123 25868
rect 1151 25804 1215 25868
rect 1243 25804 1307 25868
rect 1335 25804 1399 25868
rect 1427 25804 1491 25868
rect 967 25724 1031 25788
rect 1059 25724 1123 25788
rect 1151 25724 1215 25788
rect 1243 25724 1307 25788
rect 1335 25724 1399 25788
rect 1427 25724 1491 25788
rect 967 25644 1031 25708
rect 1059 25644 1123 25708
rect 1151 25644 1215 25708
rect 1243 25644 1307 25708
rect 1335 25644 1399 25708
rect 1427 25644 1491 25708
rect 967 25564 1031 25628
rect 1059 25564 1123 25628
rect 1151 25564 1215 25628
rect 1243 25564 1307 25628
rect 1335 25564 1399 25628
rect 1427 25564 1491 25628
rect 967 25483 1031 25547
rect 1059 25483 1123 25547
rect 1151 25483 1215 25547
rect 1243 25483 1307 25547
rect 1335 25483 1399 25547
rect 1427 25483 1491 25547
rect 967 25402 1031 25466
rect 1059 25402 1123 25466
rect 1151 25402 1215 25466
rect 1243 25402 1307 25466
rect 1335 25402 1399 25466
rect 1427 25402 1491 25466
rect 967 25321 1031 25385
rect 1059 25321 1123 25385
rect 1151 25321 1215 25385
rect 1243 25321 1307 25385
rect 1335 25321 1399 25385
rect 1427 25321 1491 25385
rect 967 25240 1031 25304
rect 1059 25240 1123 25304
rect 1151 25240 1215 25304
rect 1243 25240 1307 25304
rect 1335 25240 1399 25304
rect 1427 25240 1491 25304
rect 967 25159 1031 25223
rect 1059 25159 1123 25223
rect 1151 25159 1215 25223
rect 1243 25159 1307 25223
rect 1335 25159 1399 25223
rect 1427 25159 1491 25223
rect 967 25078 1031 25142
rect 1059 25078 1123 25142
rect 1151 25078 1215 25142
rect 1243 25078 1307 25142
rect 1335 25078 1399 25142
rect 1427 25078 1491 25142
rect 967 24997 1031 25061
rect 1059 24997 1123 25061
rect 1151 24997 1215 25061
rect 1243 24997 1307 25061
rect 1335 24997 1399 25061
rect 1427 24997 1491 25061
rect 967 24916 1031 24980
rect 1059 24916 1123 24980
rect 1151 24916 1215 24980
rect 1243 24916 1307 24980
rect 1335 24916 1399 24980
rect 1427 24916 1491 24980
rect 967 24835 1031 24899
rect 1059 24835 1123 24899
rect 1151 24835 1215 24899
rect 1243 24835 1307 24899
rect 1335 24835 1399 24899
rect 1427 24835 1491 24899
rect 967 24754 1031 24818
rect 1059 24754 1123 24818
rect 1151 24754 1215 24818
rect 1243 24754 1307 24818
rect 1335 24754 1399 24818
rect 1427 24754 1491 24818
rect 967 24673 1031 24737
rect 1059 24673 1123 24737
rect 1151 24673 1215 24737
rect 1243 24673 1307 24737
rect 1335 24673 1399 24737
rect 1427 24673 1491 24737
rect 967 24592 1031 24656
rect 1059 24592 1123 24656
rect 1151 24592 1215 24656
rect 1243 24592 1307 24656
rect 1335 24592 1399 24656
rect 1427 24592 1491 24656
rect 967 24511 1031 24575
rect 1059 24511 1123 24575
rect 1151 24511 1215 24575
rect 1243 24511 1307 24575
rect 1335 24511 1399 24575
rect 1427 24511 1491 24575
rect 967 24430 1031 24494
rect 1059 24430 1123 24494
rect 1151 24430 1215 24494
rect 1243 24430 1307 24494
rect 1335 24430 1399 24494
rect 1427 24430 1491 24494
rect 967 24349 1031 24413
rect 1059 24349 1123 24413
rect 1151 24349 1215 24413
rect 1243 24349 1307 24413
rect 1335 24349 1399 24413
rect 1427 24349 1491 24413
rect 967 24268 1031 24332
rect 1059 24268 1123 24332
rect 1151 24268 1215 24332
rect 1243 24268 1307 24332
rect 1335 24268 1399 24332
rect 1427 24268 1491 24332
rect 967 24187 1031 24251
rect 1059 24187 1123 24251
rect 1151 24187 1215 24251
rect 1243 24187 1307 24251
rect 1335 24187 1399 24251
rect 1427 24187 1491 24251
rect 967 24106 1031 24170
rect 1059 24106 1123 24170
rect 1151 24106 1215 24170
rect 1243 24106 1307 24170
rect 1335 24106 1399 24170
rect 1427 24106 1491 24170
rect 967 24025 1031 24089
rect 1059 24025 1123 24089
rect 1151 24025 1215 24089
rect 1243 24025 1307 24089
rect 1335 24025 1399 24089
rect 1427 24025 1491 24089
rect 967 23944 1031 24008
rect 1059 23944 1123 24008
rect 1151 23944 1215 24008
rect 1243 23944 1307 24008
rect 1335 23944 1399 24008
rect 1427 23944 1491 24008
rect 967 23863 1031 23927
rect 1059 23863 1123 23927
rect 1151 23863 1215 23927
rect 1243 23863 1307 23927
rect 1335 23863 1399 23927
rect 1427 23863 1491 23927
rect 967 23782 1031 23846
rect 1059 23782 1123 23846
rect 1151 23782 1215 23846
rect 1243 23782 1307 23846
rect 1335 23782 1399 23846
rect 1427 23782 1491 23846
rect 967 23701 1031 23765
rect 1059 23701 1123 23765
rect 1151 23701 1215 23765
rect 1243 23701 1307 23765
rect 1335 23701 1399 23765
rect 1427 23701 1491 23765
rect 967 23620 1031 23684
rect 1059 23620 1123 23684
rect 1151 23620 1215 23684
rect 1243 23620 1307 23684
rect 1335 23620 1399 23684
rect 1427 23620 1491 23684
rect 967 23539 1031 23603
rect 1059 23539 1123 23603
rect 1151 23539 1215 23603
rect 1243 23539 1307 23603
rect 1335 23539 1399 23603
rect 1427 23539 1491 23603
rect 967 23458 1031 23522
rect 1059 23458 1123 23522
rect 1151 23458 1215 23522
rect 1243 23458 1307 23522
rect 1335 23458 1399 23522
rect 1427 23458 1491 23522
rect 967 23377 1031 23441
rect 1059 23377 1123 23441
rect 1151 23377 1215 23441
rect 1243 23377 1307 23441
rect 1335 23377 1399 23441
rect 1427 23377 1491 23441
rect 967 23296 1031 23360
rect 1059 23296 1123 23360
rect 1151 23296 1215 23360
rect 1243 23296 1307 23360
rect 1335 23296 1399 23360
rect 1427 23296 1491 23360
rect 967 23215 1031 23279
rect 1059 23215 1123 23279
rect 1151 23215 1215 23279
rect 1243 23215 1307 23279
rect 1335 23215 1399 23279
rect 1427 23215 1491 23279
rect 967 23134 1031 23198
rect 1059 23134 1123 23198
rect 1151 23134 1215 23198
rect 1243 23134 1307 23198
rect 1335 23134 1399 23198
rect 1427 23134 1491 23198
rect 967 23053 1031 23117
rect 1059 23053 1123 23117
rect 1151 23053 1215 23117
rect 1243 23053 1307 23117
rect 1335 23053 1399 23117
rect 1427 23053 1491 23117
rect 967 22972 1031 23036
rect 1059 22972 1123 23036
rect 1151 22972 1215 23036
rect 1243 22972 1307 23036
rect 1335 22972 1399 23036
rect 1427 22972 1491 23036
rect 967 22891 1031 22955
rect 1059 22891 1123 22955
rect 1151 22891 1215 22955
rect 1243 22891 1307 22955
rect 1335 22891 1399 22955
rect 1427 22891 1491 22955
rect 967 22810 1031 22874
rect 1059 22810 1123 22874
rect 1151 22810 1215 22874
rect 1243 22810 1307 22874
rect 1335 22810 1399 22874
rect 1427 22810 1491 22874
rect 967 22729 1031 22793
rect 1059 22729 1123 22793
rect 1151 22729 1215 22793
rect 1243 22729 1307 22793
rect 1335 22729 1399 22793
rect 1427 22729 1491 22793
rect 967 22648 1031 22712
rect 1059 22648 1123 22712
rect 1151 22648 1215 22712
rect 1243 22648 1307 22712
rect 1335 22648 1399 22712
rect 1427 22648 1491 22712
rect 967 22567 1031 22631
rect 1059 22567 1123 22631
rect 1151 22567 1215 22631
rect 1243 22567 1307 22631
rect 1335 22567 1399 22631
rect 1427 22567 1491 22631
rect 967 22486 1031 22550
rect 1059 22486 1123 22550
rect 1151 22486 1215 22550
rect 1243 22486 1307 22550
rect 1335 22486 1399 22550
rect 1427 22486 1491 22550
rect 967 22405 1031 22469
rect 1059 22405 1123 22469
rect 1151 22405 1215 22469
rect 1243 22405 1307 22469
rect 1335 22405 1399 22469
rect 1427 22405 1491 22469
rect 967 22324 1031 22388
rect 1059 22324 1123 22388
rect 1151 22324 1215 22388
rect 1243 22324 1307 22388
rect 1335 22324 1399 22388
rect 1427 22324 1491 22388
rect 967 22243 1031 22307
rect 1059 22243 1123 22307
rect 1151 22243 1215 22307
rect 1243 22243 1307 22307
rect 1335 22243 1399 22307
rect 1427 22243 1491 22307
rect 967 22162 1031 22226
rect 1059 22162 1123 22226
rect 1151 22162 1215 22226
rect 1243 22162 1307 22226
rect 1335 22162 1399 22226
rect 1427 22162 1491 22226
rect 967 22081 1031 22145
rect 1059 22081 1123 22145
rect 1151 22081 1215 22145
rect 1243 22081 1307 22145
rect 1335 22081 1399 22145
rect 1427 22081 1491 22145
rect 967 22000 1031 22064
rect 1059 22000 1123 22064
rect 1151 22000 1215 22064
rect 1243 22000 1307 22064
rect 1335 22000 1399 22064
rect 1427 22000 1491 22064
rect 967 21919 1031 21983
rect 1059 21919 1123 21983
rect 1151 21919 1215 21983
rect 1243 21919 1307 21983
rect 1335 21919 1399 21983
rect 1427 21919 1491 21983
rect 967 21838 1031 21902
rect 1059 21838 1123 21902
rect 1151 21838 1215 21902
rect 1243 21838 1307 21902
rect 1335 21838 1399 21902
rect 1427 21838 1491 21902
rect 967 21757 1031 21821
rect 1059 21757 1123 21821
rect 1151 21757 1215 21821
rect 1243 21757 1307 21821
rect 1335 21757 1399 21821
rect 1427 21757 1491 21821
rect 967 21676 1031 21740
rect 1059 21676 1123 21740
rect 1151 21676 1215 21740
rect 1243 21676 1307 21740
rect 1335 21676 1399 21740
rect 1427 21676 1491 21740
rect 967 21595 1031 21659
rect 1059 21595 1123 21659
rect 1151 21595 1215 21659
rect 1243 21595 1307 21659
rect 1335 21595 1399 21659
rect 1427 21595 1491 21659
rect 967 21514 1031 21578
rect 1059 21514 1123 21578
rect 1151 21514 1215 21578
rect 1243 21514 1307 21578
rect 1335 21514 1399 21578
rect 1427 21514 1491 21578
rect 967 21433 1031 21497
rect 1059 21433 1123 21497
rect 1151 21433 1215 21497
rect 1243 21433 1307 21497
rect 1335 21433 1399 21497
rect 1427 21433 1491 21497
rect 967 21352 1031 21416
rect 1059 21352 1123 21416
rect 1151 21352 1215 21416
rect 1243 21352 1307 21416
rect 1335 21352 1399 21416
rect 1427 21352 1491 21416
rect 967 21271 1031 21335
rect 1059 21271 1123 21335
rect 1151 21271 1215 21335
rect 1243 21271 1307 21335
rect 1335 21271 1399 21335
rect 1427 21271 1491 21335
rect 967 21190 1031 21254
rect 1059 21190 1123 21254
rect 1151 21190 1215 21254
rect 1243 21190 1307 21254
rect 1335 21190 1399 21254
rect 1427 21190 1491 21254
rect 967 21109 1031 21173
rect 1059 21109 1123 21173
rect 1151 21109 1215 21173
rect 1243 21109 1307 21173
rect 1335 21109 1399 21173
rect 1427 21109 1491 21173
rect 967 21028 1031 21092
rect 1059 21028 1123 21092
rect 1151 21028 1215 21092
rect 1243 21028 1307 21092
rect 1335 21028 1399 21092
rect 1427 21028 1491 21092
rect 967 20947 1031 21011
rect 1059 20947 1123 21011
rect 1151 20947 1215 21011
rect 1243 20947 1307 21011
rect 1335 20947 1399 21011
rect 1427 20947 1491 21011
rect 967 20866 1031 20930
rect 1059 20866 1123 20930
rect 1151 20866 1215 20930
rect 1243 20866 1307 20930
rect 1335 20866 1399 20930
rect 1427 20866 1491 20930
rect 967 20785 1031 20849
rect 1059 20785 1123 20849
rect 1151 20785 1215 20849
rect 1243 20785 1307 20849
rect 1335 20785 1399 20849
rect 1427 20785 1491 20849
rect 967 20704 1031 20768
rect 1059 20704 1123 20768
rect 1151 20704 1215 20768
rect 1243 20704 1307 20768
rect 1335 20704 1399 20768
rect 1427 20704 1491 20768
rect 967 20623 1031 20687
rect 1059 20623 1123 20687
rect 1151 20623 1215 20687
rect 1243 20623 1307 20687
rect 1335 20623 1399 20687
rect 1427 20623 1491 20687
rect 967 20542 1031 20606
rect 1059 20542 1123 20606
rect 1151 20542 1215 20606
rect 1243 20542 1307 20606
rect 1335 20542 1399 20606
rect 1427 20542 1491 20606
rect 967 20461 1031 20525
rect 1059 20461 1123 20525
rect 1151 20461 1215 20525
rect 1243 20461 1307 20525
rect 1335 20461 1399 20525
rect 1427 20461 1491 20525
rect 1543 20470 1607 20534
rect 1089 20351 1153 20415
rect 1215 20367 1279 20431
rect 1297 20367 1361 20431
rect 1379 20367 1443 20431
rect 1461 20367 1525 20431
rect 1543 20367 1607 20431
rect 1624 20367 1688 20431
rect 1215 20219 1279 20283
rect 1297 20219 1361 20283
rect 1379 20219 1443 20283
rect 1461 20219 1525 20283
rect 1543 20219 1607 20283
rect 1624 20219 1688 20283
rect 1766 20247 1830 20311
rect 1312 20128 1376 20192
rect 1471 20139 1535 20203
rect 1553 20139 1617 20203
rect 1635 20139 1699 20203
rect 1717 20139 1781 20203
rect 1799 20139 1863 20203
rect 1880 20139 1944 20203
rect 1471 19991 1535 20055
rect 1553 19991 1617 20055
rect 1635 19991 1699 20055
rect 1717 19991 1781 20055
rect 1799 19991 1863 20055
rect 1880 19991 1944 20055
rect 2005 20008 2069 20072
rect 1551 19889 1615 19953
rect 1669 19911 1733 19975
rect 1751 19911 1815 19975
rect 1833 19911 1897 19975
rect 1915 19911 1979 19975
rect 1997 19911 2061 19975
rect 2078 19911 2142 19975
rect 1669 19763 1733 19827
rect 1751 19763 1815 19827
rect 1833 19763 1897 19827
rect 1915 19763 1979 19827
rect 1997 19763 2061 19827
rect 2078 19763 2142 19827
rect 2220 19793 2284 19857
rect 1766 19674 1830 19738
rect 1893 19678 1957 19742
rect 1975 19678 2039 19742
rect 2057 19678 2121 19742
rect 2139 19678 2203 19742
rect 2221 19678 2285 19742
rect 2302 19678 2366 19742
rect 2394 19594 2458 19658
rect 2502 19594 2566 19658
rect 1893 19530 1957 19594
rect 1975 19530 2039 19594
rect 2057 19530 2121 19594
rect 2139 19530 2203 19594
rect 2221 19530 2285 19594
rect 2302 19530 2366 19594
rect 1998 19435 2062 19499
rect 2120 19444 2184 19508
rect 2211 19444 2275 19508
rect 2302 19444 2366 19508
rect 2394 19485 2458 19549
rect 2502 19485 2566 19549
rect 2394 19376 2458 19440
rect 2502 19376 2566 19440
rect 2120 19296 2184 19360
rect 2211 19296 2275 19360
rect 2302 19296 2366 19360
rect 2220 19211 2284 19275
rect 2305 19211 2369 19275
rect 2394 19268 2458 19332
rect 2502 19268 2566 19332
rect 2394 19160 2458 19224
rect 2502 19160 2566 19224
rect 12446 34133 12510 34197
rect 12554 34133 12618 34197
rect 12446 34025 12510 34089
rect 12554 34025 12618 34089
rect 12646 33981 12710 34045
rect 12737 33981 12801 34045
rect 12828 33981 12892 34045
rect 12446 33917 12510 33981
rect 12554 33917 12618 33981
rect 12446 33808 12510 33872
rect 12554 33808 12618 33872
rect 12646 33833 12710 33897
rect 12737 33833 12801 33897
rect 12828 33833 12892 33897
rect 12950 33851 13014 33915
rect 12446 33699 12510 33763
rect 12554 33699 12618 33763
rect 12648 33736 12712 33800
rect 12777 33736 12841 33800
rect 12906 33736 12970 33800
rect 13034 33736 13098 33800
rect 12648 33634 12712 33698
rect 12777 33634 12841 33698
rect 12906 33634 12970 33698
rect 13034 33634 13098 33698
rect 13182 33619 13246 33683
rect 12728 33500 12792 33564
rect 12870 33530 12934 33594
rect 12951 33530 13015 33594
rect 13033 33530 13097 33594
rect 13115 33530 13179 33594
rect 13197 33530 13261 33594
rect 13279 33530 13343 33594
rect 12870 33382 12934 33446
rect 12951 33382 13015 33446
rect 13033 33382 13097 33446
rect 13115 33382 13179 33446
rect 13197 33382 13261 33446
rect 13279 33382 13343 33446
rect 13397 33404 13461 33468
rect 12943 33285 13007 33349
rect 13068 33302 13132 33366
rect 13149 33302 13213 33366
rect 13231 33302 13295 33366
rect 13313 33302 13377 33366
rect 13395 33302 13459 33366
rect 13477 33302 13541 33366
rect 13068 33154 13132 33218
rect 13149 33154 13213 33218
rect 13231 33154 13295 33218
rect 13313 33154 13377 33218
rect 13395 33154 13459 33218
rect 13477 33154 13541 33218
rect 13636 33165 13700 33229
rect 13182 33046 13246 33110
rect 13324 33074 13388 33138
rect 13405 33074 13469 33138
rect 13487 33074 13551 33138
rect 13569 33074 13633 33138
rect 13651 33074 13715 33138
rect 13733 33074 13797 33138
rect 13324 32926 13388 32990
rect 13405 32926 13469 32990
rect 13487 32926 13551 32990
rect 13569 32926 13633 32990
rect 13651 32926 13715 32990
rect 13733 32926 13797 32990
rect 13859 32942 13923 33006
rect 13405 32823 13469 32887
rect 13506 32805 13570 32869
rect 13598 32805 13662 32869
rect 13690 32805 13754 32869
rect 13782 32805 13846 32869
rect 13874 32805 13938 32869
rect 13966 32805 14030 32869
rect 13506 32725 13570 32789
rect 13598 32725 13662 32789
rect 13690 32725 13754 32789
rect 13782 32725 13846 32789
rect 13874 32725 13938 32789
rect 13966 32725 14030 32789
rect 13506 32645 13570 32709
rect 13598 32645 13662 32709
rect 13690 32645 13754 32709
rect 13782 32645 13846 32709
rect 13874 32645 13938 32709
rect 13966 32645 14030 32709
rect 13506 32565 13570 32629
rect 13598 32565 13662 32629
rect 13690 32565 13754 32629
rect 13782 32565 13846 32629
rect 13874 32565 13938 32629
rect 13966 32565 14030 32629
rect 13506 32485 13570 32549
rect 13598 32485 13662 32549
rect 13690 32485 13754 32549
rect 13782 32485 13846 32549
rect 13874 32485 13938 32549
rect 13966 32485 14030 32549
rect 13506 32405 13570 32469
rect 13598 32405 13662 32469
rect 13690 32405 13754 32469
rect 13782 32405 13846 32469
rect 13874 32405 13938 32469
rect 13966 32405 14030 32469
rect 13506 32325 13570 32389
rect 13598 32325 13662 32389
rect 13690 32325 13754 32389
rect 13782 32325 13846 32389
rect 13874 32325 13938 32389
rect 13966 32325 14030 32389
rect 13506 32245 13570 32309
rect 13598 32245 13662 32309
rect 13690 32245 13754 32309
rect 13782 32245 13846 32309
rect 13874 32245 13938 32309
rect 13966 32245 14030 32309
rect 13506 32165 13570 32229
rect 13598 32165 13662 32229
rect 13690 32165 13754 32229
rect 13782 32165 13846 32229
rect 13874 32165 13938 32229
rect 13966 32165 14030 32229
rect 13506 32085 13570 32149
rect 13598 32085 13662 32149
rect 13690 32085 13754 32149
rect 13782 32085 13846 32149
rect 13874 32085 13938 32149
rect 13966 32085 14030 32149
rect 13506 32005 13570 32069
rect 13598 32005 13662 32069
rect 13690 32005 13754 32069
rect 13782 32005 13846 32069
rect 13874 32005 13938 32069
rect 13966 32005 14030 32069
rect 13506 31925 13570 31989
rect 13598 31925 13662 31989
rect 13690 31925 13754 31989
rect 13782 31925 13846 31989
rect 13874 31925 13938 31989
rect 13966 31925 14030 31989
rect 13506 31845 13570 31909
rect 13598 31845 13662 31909
rect 13690 31845 13754 31909
rect 13782 31845 13846 31909
rect 13874 31845 13938 31909
rect 13966 31845 14030 31909
rect 13506 31765 13570 31829
rect 13598 31765 13662 31829
rect 13690 31765 13754 31829
rect 13782 31765 13846 31829
rect 13874 31765 13938 31829
rect 13966 31765 14030 31829
rect 13506 31685 13570 31749
rect 13598 31685 13662 31749
rect 13690 31685 13754 31749
rect 13782 31685 13846 31749
rect 13874 31685 13938 31749
rect 13966 31685 14030 31749
rect 13506 31605 13570 31669
rect 13598 31605 13662 31669
rect 13690 31605 13754 31669
rect 13782 31605 13846 31669
rect 13874 31605 13938 31669
rect 13966 31605 14030 31669
rect 13506 31525 13570 31589
rect 13598 31525 13662 31589
rect 13690 31525 13754 31589
rect 13782 31525 13846 31589
rect 13874 31525 13938 31589
rect 13966 31525 14030 31589
rect 13506 31445 13570 31509
rect 13598 31445 13662 31509
rect 13690 31445 13754 31509
rect 13782 31445 13846 31509
rect 13874 31445 13938 31509
rect 13966 31445 14030 31509
rect 13506 31365 13570 31429
rect 13598 31365 13662 31429
rect 13690 31365 13754 31429
rect 13782 31365 13846 31429
rect 13874 31365 13938 31429
rect 13966 31365 14030 31429
rect 13506 31285 13570 31349
rect 13598 31285 13662 31349
rect 13690 31285 13754 31349
rect 13782 31285 13846 31349
rect 13874 31285 13938 31349
rect 13966 31285 14030 31349
rect 13506 31205 13570 31269
rect 13598 31205 13662 31269
rect 13690 31205 13754 31269
rect 13782 31205 13846 31269
rect 13874 31205 13938 31269
rect 13966 31205 14030 31269
rect 13506 31125 13570 31189
rect 13598 31125 13662 31189
rect 13690 31125 13754 31189
rect 13782 31125 13846 31189
rect 13874 31125 13938 31189
rect 13966 31125 14030 31189
rect 13506 31045 13570 31109
rect 13598 31045 13662 31109
rect 13690 31045 13754 31109
rect 13782 31045 13846 31109
rect 13874 31045 13938 31109
rect 13966 31045 14030 31109
rect 13506 30965 13570 31029
rect 13598 30965 13662 31029
rect 13690 30965 13754 31029
rect 13782 30965 13846 31029
rect 13874 30965 13938 31029
rect 13966 30965 14030 31029
rect 13506 30885 13570 30949
rect 13598 30885 13662 30949
rect 13690 30885 13754 30949
rect 13782 30885 13846 30949
rect 13874 30885 13938 30949
rect 13966 30885 14030 30949
rect 13506 30805 13570 30869
rect 13598 30805 13662 30869
rect 13690 30805 13754 30869
rect 13782 30805 13846 30869
rect 13874 30805 13938 30869
rect 13966 30805 14030 30869
rect 13506 30725 13570 30789
rect 13598 30725 13662 30789
rect 13690 30725 13754 30789
rect 13782 30725 13846 30789
rect 13874 30725 13938 30789
rect 13966 30725 14030 30789
rect 13506 30645 13570 30709
rect 13598 30645 13662 30709
rect 13690 30645 13754 30709
rect 13782 30645 13846 30709
rect 13874 30645 13938 30709
rect 13966 30645 14030 30709
rect 13506 30565 13570 30629
rect 13598 30565 13662 30629
rect 13690 30565 13754 30629
rect 13782 30565 13846 30629
rect 13874 30565 13938 30629
rect 13966 30565 14030 30629
rect 13506 30485 13570 30549
rect 13598 30485 13662 30549
rect 13690 30485 13754 30549
rect 13782 30485 13846 30549
rect 13874 30485 13938 30549
rect 13966 30485 14030 30549
rect 13506 30405 13570 30469
rect 13598 30405 13662 30469
rect 13690 30405 13754 30469
rect 13782 30405 13846 30469
rect 13874 30405 13938 30469
rect 13966 30405 14030 30469
rect 13506 30325 13570 30389
rect 13598 30325 13662 30389
rect 13690 30325 13754 30389
rect 13782 30325 13846 30389
rect 13874 30325 13938 30389
rect 13966 30325 14030 30389
rect 13506 30245 13570 30309
rect 13598 30245 13662 30309
rect 13690 30245 13754 30309
rect 13782 30245 13846 30309
rect 13874 30245 13938 30309
rect 13966 30245 14030 30309
rect 13506 30165 13570 30229
rect 13598 30165 13662 30229
rect 13690 30165 13754 30229
rect 13782 30165 13846 30229
rect 13874 30165 13938 30229
rect 13966 30165 14030 30229
rect 13506 30085 13570 30149
rect 13598 30085 13662 30149
rect 13690 30085 13754 30149
rect 13782 30085 13846 30149
rect 13874 30085 13938 30149
rect 13966 30085 14030 30149
rect 13506 30005 13570 30069
rect 13598 30005 13662 30069
rect 13690 30005 13754 30069
rect 13782 30005 13846 30069
rect 13874 30005 13938 30069
rect 13966 30005 14030 30069
rect 13506 29925 13570 29989
rect 13598 29925 13662 29989
rect 13690 29925 13754 29989
rect 13782 29925 13846 29989
rect 13874 29925 13938 29989
rect 13966 29925 14030 29989
rect 13506 29845 13570 29909
rect 13598 29845 13662 29909
rect 13690 29845 13754 29909
rect 13782 29845 13846 29909
rect 13874 29845 13938 29909
rect 13966 29845 14030 29909
rect 13506 29765 13570 29829
rect 13598 29765 13662 29829
rect 13690 29765 13754 29829
rect 13782 29765 13846 29829
rect 13874 29765 13938 29829
rect 13966 29765 14030 29829
rect 13506 29685 13570 29749
rect 13598 29685 13662 29749
rect 13690 29685 13754 29749
rect 13782 29685 13846 29749
rect 13874 29685 13938 29749
rect 13966 29685 14030 29749
rect 13506 29605 13570 29669
rect 13598 29605 13662 29669
rect 13690 29605 13754 29669
rect 13782 29605 13846 29669
rect 13874 29605 13938 29669
rect 13966 29605 14030 29669
rect 13506 29525 13570 29589
rect 13598 29525 13662 29589
rect 13690 29525 13754 29589
rect 13782 29525 13846 29589
rect 13874 29525 13938 29589
rect 13966 29525 14030 29589
rect 13506 29445 13570 29509
rect 13598 29445 13662 29509
rect 13690 29445 13754 29509
rect 13782 29445 13846 29509
rect 13874 29445 13938 29509
rect 13966 29445 14030 29509
rect 13506 29365 13570 29429
rect 13598 29365 13662 29429
rect 13690 29365 13754 29429
rect 13782 29365 13846 29429
rect 13874 29365 13938 29429
rect 13966 29365 14030 29429
rect 13506 29285 13570 29349
rect 13598 29285 13662 29349
rect 13690 29285 13754 29349
rect 13782 29285 13846 29349
rect 13874 29285 13938 29349
rect 13966 29285 14030 29349
rect 13506 29205 13570 29269
rect 13598 29205 13662 29269
rect 13690 29205 13754 29269
rect 13782 29205 13846 29269
rect 13874 29205 13938 29269
rect 13966 29205 14030 29269
rect 13506 29125 13570 29189
rect 13598 29125 13662 29189
rect 13690 29125 13754 29189
rect 13782 29125 13846 29189
rect 13874 29125 13938 29189
rect 13966 29125 14030 29189
rect 13506 29045 13570 29109
rect 13598 29045 13662 29109
rect 13690 29045 13754 29109
rect 13782 29045 13846 29109
rect 13874 29045 13938 29109
rect 13966 29045 14030 29109
rect 13506 28965 13570 29029
rect 13598 28965 13662 29029
rect 13690 28965 13754 29029
rect 13782 28965 13846 29029
rect 13874 28965 13938 29029
rect 13966 28965 14030 29029
rect 13506 28885 13570 28949
rect 13598 28885 13662 28949
rect 13690 28885 13754 28949
rect 13782 28885 13846 28949
rect 13874 28885 13938 28949
rect 13966 28885 14030 28949
rect 13506 28805 13570 28869
rect 13598 28805 13662 28869
rect 13690 28805 13754 28869
rect 13782 28805 13846 28869
rect 13874 28805 13938 28869
rect 13966 28805 14030 28869
rect 13506 28725 13570 28789
rect 13598 28725 13662 28789
rect 13690 28725 13754 28789
rect 13782 28725 13846 28789
rect 13874 28725 13938 28789
rect 13966 28725 14030 28789
rect 13506 28645 13570 28709
rect 13598 28645 13662 28709
rect 13690 28645 13754 28709
rect 13782 28645 13846 28709
rect 13874 28645 13938 28709
rect 13966 28645 14030 28709
rect 13506 28565 13570 28629
rect 13598 28565 13662 28629
rect 13690 28565 13754 28629
rect 13782 28565 13846 28629
rect 13874 28565 13938 28629
rect 13966 28565 14030 28629
rect 13506 28485 13570 28549
rect 13598 28485 13662 28549
rect 13690 28485 13754 28549
rect 13782 28485 13846 28549
rect 13874 28485 13938 28549
rect 13966 28485 14030 28549
rect 13506 28405 13570 28469
rect 13598 28405 13662 28469
rect 13690 28405 13754 28469
rect 13782 28405 13846 28469
rect 13874 28405 13938 28469
rect 13966 28405 14030 28469
rect 13506 28325 13570 28389
rect 13598 28325 13662 28389
rect 13690 28325 13754 28389
rect 13782 28325 13846 28389
rect 13874 28325 13938 28389
rect 13966 28325 14030 28389
rect 13506 28245 13570 28309
rect 13598 28245 13662 28309
rect 13690 28245 13754 28309
rect 13782 28245 13846 28309
rect 13874 28245 13938 28309
rect 13966 28245 14030 28309
rect 13506 28165 13570 28229
rect 13598 28165 13662 28229
rect 13690 28165 13754 28229
rect 13782 28165 13846 28229
rect 13874 28165 13938 28229
rect 13966 28165 14030 28229
rect 13506 28085 13570 28149
rect 13598 28085 13662 28149
rect 13690 28085 13754 28149
rect 13782 28085 13846 28149
rect 13874 28085 13938 28149
rect 13966 28085 14030 28149
rect 13506 28005 13570 28069
rect 13598 28005 13662 28069
rect 13690 28005 13754 28069
rect 13782 28005 13846 28069
rect 13874 28005 13938 28069
rect 13966 28005 14030 28069
rect 13506 27925 13570 27989
rect 13598 27925 13662 27989
rect 13690 27925 13754 27989
rect 13782 27925 13846 27989
rect 13874 27925 13938 27989
rect 13966 27925 14030 27989
rect 13506 27845 13570 27909
rect 13598 27845 13662 27909
rect 13690 27845 13754 27909
rect 13782 27845 13846 27909
rect 13874 27845 13938 27909
rect 13966 27845 14030 27909
rect 13506 27765 13570 27829
rect 13598 27765 13662 27829
rect 13690 27765 13754 27829
rect 13782 27765 13846 27829
rect 13874 27765 13938 27829
rect 13966 27765 14030 27829
rect 13506 27685 13570 27749
rect 13598 27685 13662 27749
rect 13690 27685 13754 27749
rect 13782 27685 13846 27749
rect 13874 27685 13938 27749
rect 13966 27685 14030 27749
rect 13506 27605 13570 27669
rect 13598 27605 13662 27669
rect 13690 27605 13754 27669
rect 13782 27605 13846 27669
rect 13874 27605 13938 27669
rect 13966 27605 14030 27669
rect 13506 27525 13570 27589
rect 13598 27525 13662 27589
rect 13690 27525 13754 27589
rect 13782 27525 13846 27589
rect 13874 27525 13938 27589
rect 13966 27525 14030 27589
rect 13506 27445 13570 27509
rect 13598 27445 13662 27509
rect 13690 27445 13754 27509
rect 13782 27445 13846 27509
rect 13874 27445 13938 27509
rect 13966 27445 14030 27509
rect 13506 27365 13570 27429
rect 13598 27365 13662 27429
rect 13690 27365 13754 27429
rect 13782 27365 13846 27429
rect 13874 27365 13938 27429
rect 13966 27365 14030 27429
rect 13506 27285 13570 27349
rect 13598 27285 13662 27349
rect 13690 27285 13754 27349
rect 13782 27285 13846 27349
rect 13874 27285 13938 27349
rect 13966 27285 14030 27349
rect 13506 27205 13570 27269
rect 13598 27205 13662 27269
rect 13690 27205 13754 27269
rect 13782 27205 13846 27269
rect 13874 27205 13938 27269
rect 13966 27205 14030 27269
rect 13506 27125 13570 27189
rect 13598 27125 13662 27189
rect 13690 27125 13754 27189
rect 13782 27125 13846 27189
rect 13874 27125 13938 27189
rect 13966 27125 14030 27189
rect 13506 27045 13570 27109
rect 13598 27045 13662 27109
rect 13690 27045 13754 27109
rect 13782 27045 13846 27109
rect 13874 27045 13938 27109
rect 13966 27045 14030 27109
rect 13506 26965 13570 27029
rect 13598 26965 13662 27029
rect 13690 26965 13754 27029
rect 13782 26965 13846 27029
rect 13874 26965 13938 27029
rect 13966 26965 14030 27029
rect 13506 26885 13570 26949
rect 13598 26885 13662 26949
rect 13690 26885 13754 26949
rect 13782 26885 13846 26949
rect 13874 26885 13938 26949
rect 13966 26885 14030 26949
rect 13506 26805 13570 26869
rect 13598 26805 13662 26869
rect 13690 26805 13754 26869
rect 13782 26805 13846 26869
rect 13874 26805 13938 26869
rect 13966 26805 14030 26869
rect 13506 26725 13570 26789
rect 13598 26725 13662 26789
rect 13690 26725 13754 26789
rect 13782 26725 13846 26789
rect 13874 26725 13938 26789
rect 13966 26725 14030 26789
rect 13506 26645 13570 26709
rect 13598 26645 13662 26709
rect 13690 26645 13754 26709
rect 13782 26645 13846 26709
rect 13874 26645 13938 26709
rect 13966 26645 14030 26709
rect 13506 26565 13570 26629
rect 13598 26565 13662 26629
rect 13690 26565 13754 26629
rect 13782 26565 13846 26629
rect 13874 26565 13938 26629
rect 13966 26565 14030 26629
rect 13506 26485 13570 26549
rect 13598 26485 13662 26549
rect 13690 26485 13754 26549
rect 13782 26485 13846 26549
rect 13874 26485 13938 26549
rect 13966 26485 14030 26549
rect 13506 26405 13570 26469
rect 13598 26405 13662 26469
rect 13690 26405 13754 26469
rect 13782 26405 13846 26469
rect 13874 26405 13938 26469
rect 13966 26405 14030 26469
rect 13506 26325 13570 26389
rect 13598 26325 13662 26389
rect 13690 26325 13754 26389
rect 13782 26325 13846 26389
rect 13874 26325 13938 26389
rect 13966 26325 14030 26389
rect 13506 26245 13570 26309
rect 13598 26245 13662 26309
rect 13690 26245 13754 26309
rect 13782 26245 13846 26309
rect 13874 26245 13938 26309
rect 13966 26245 14030 26309
rect 13506 26165 13570 26229
rect 13598 26165 13662 26229
rect 13690 26165 13754 26229
rect 13782 26165 13846 26229
rect 13874 26165 13938 26229
rect 13966 26165 14030 26229
rect 13506 26085 13570 26149
rect 13598 26085 13662 26149
rect 13690 26085 13754 26149
rect 13782 26085 13846 26149
rect 13874 26085 13938 26149
rect 13966 26085 14030 26149
rect 13506 26005 13570 26069
rect 13598 26005 13662 26069
rect 13690 26005 13754 26069
rect 13782 26005 13846 26069
rect 13874 26005 13938 26069
rect 13966 26005 14030 26069
rect 13506 25925 13570 25989
rect 13598 25925 13662 25989
rect 13690 25925 13754 25989
rect 13782 25925 13846 25989
rect 13874 25925 13938 25989
rect 13966 25925 14030 25989
rect 13506 25845 13570 25909
rect 13598 25845 13662 25909
rect 13690 25845 13754 25909
rect 13782 25845 13846 25909
rect 13874 25845 13938 25909
rect 13966 25845 14030 25909
rect 13506 25765 13570 25829
rect 13598 25765 13662 25829
rect 13690 25765 13754 25829
rect 13782 25765 13846 25829
rect 13874 25765 13938 25829
rect 13966 25765 14030 25829
rect 13506 25685 13570 25749
rect 13598 25685 13662 25749
rect 13690 25685 13754 25749
rect 13782 25685 13846 25749
rect 13874 25685 13938 25749
rect 13966 25685 14030 25749
rect 13506 25605 13570 25669
rect 13598 25605 13662 25669
rect 13690 25605 13754 25669
rect 13782 25605 13846 25669
rect 13874 25605 13938 25669
rect 13966 25605 14030 25669
rect 13506 25525 13570 25589
rect 13598 25525 13662 25589
rect 13690 25525 13754 25589
rect 13782 25525 13846 25589
rect 13874 25525 13938 25589
rect 13966 25525 14030 25589
rect 13506 25445 13570 25509
rect 13598 25445 13662 25509
rect 13690 25445 13754 25509
rect 13782 25445 13846 25509
rect 13874 25445 13938 25509
rect 13966 25445 14030 25509
rect 13506 25365 13570 25429
rect 13598 25365 13662 25429
rect 13690 25365 13754 25429
rect 13782 25365 13846 25429
rect 13874 25365 13938 25429
rect 13966 25365 14030 25429
rect 13506 25285 13570 25349
rect 13598 25285 13662 25349
rect 13690 25285 13754 25349
rect 13782 25285 13846 25349
rect 13874 25285 13938 25349
rect 13966 25285 14030 25349
rect 13506 25205 13570 25269
rect 13598 25205 13662 25269
rect 13690 25205 13754 25269
rect 13782 25205 13846 25269
rect 13874 25205 13938 25269
rect 13966 25205 14030 25269
rect 13506 25125 13570 25189
rect 13598 25125 13662 25189
rect 13690 25125 13754 25189
rect 13782 25125 13846 25189
rect 13874 25125 13938 25189
rect 13966 25125 14030 25189
rect 13506 25045 13570 25109
rect 13598 25045 13662 25109
rect 13690 25045 13754 25109
rect 13782 25045 13846 25109
rect 13874 25045 13938 25109
rect 13966 25045 14030 25109
rect 13506 24965 13570 25029
rect 13598 24965 13662 25029
rect 13690 24965 13754 25029
rect 13782 24965 13846 25029
rect 13874 24965 13938 25029
rect 13966 24965 14030 25029
rect 13506 24885 13570 24949
rect 13598 24885 13662 24949
rect 13690 24885 13754 24949
rect 13782 24885 13846 24949
rect 13874 24885 13938 24949
rect 13966 24885 14030 24949
rect 13506 24805 13570 24869
rect 13598 24805 13662 24869
rect 13690 24805 13754 24869
rect 13782 24805 13846 24869
rect 13874 24805 13938 24869
rect 13966 24805 14030 24869
rect 13506 24725 13570 24789
rect 13598 24725 13662 24789
rect 13690 24725 13754 24789
rect 13782 24725 13846 24789
rect 13874 24725 13938 24789
rect 13966 24725 14030 24789
rect 13506 24645 13570 24709
rect 13598 24645 13662 24709
rect 13690 24645 13754 24709
rect 13782 24645 13846 24709
rect 13874 24645 13938 24709
rect 13966 24645 14030 24709
rect 13506 24565 13570 24629
rect 13598 24565 13662 24629
rect 13690 24565 13754 24629
rect 13782 24565 13846 24629
rect 13874 24565 13938 24629
rect 13966 24565 14030 24629
rect 13506 24485 13570 24549
rect 13598 24485 13662 24549
rect 13690 24485 13754 24549
rect 13782 24485 13846 24549
rect 13874 24485 13938 24549
rect 13966 24485 14030 24549
rect 13506 24405 13570 24469
rect 13598 24405 13662 24469
rect 13690 24405 13754 24469
rect 13782 24405 13846 24469
rect 13874 24405 13938 24469
rect 13966 24405 14030 24469
rect 13506 24325 13570 24389
rect 13598 24325 13662 24389
rect 13690 24325 13754 24389
rect 13782 24325 13846 24389
rect 13874 24325 13938 24389
rect 13966 24325 14030 24389
rect 13506 24245 13570 24309
rect 13598 24245 13662 24309
rect 13690 24245 13754 24309
rect 13782 24245 13846 24309
rect 13874 24245 13938 24309
rect 13966 24245 14030 24309
rect 13506 24165 13570 24229
rect 13598 24165 13662 24229
rect 13690 24165 13754 24229
rect 13782 24165 13846 24229
rect 13874 24165 13938 24229
rect 13966 24165 14030 24229
rect 13506 24084 13570 24148
rect 13598 24084 13662 24148
rect 13690 24084 13754 24148
rect 13782 24084 13846 24148
rect 13874 24084 13938 24148
rect 13966 24084 14030 24148
rect 13506 24003 13570 24067
rect 13598 24003 13662 24067
rect 13690 24003 13754 24067
rect 13782 24003 13846 24067
rect 13874 24003 13938 24067
rect 13966 24003 14030 24067
rect 13506 23922 13570 23986
rect 13598 23922 13662 23986
rect 13690 23922 13754 23986
rect 13782 23922 13846 23986
rect 13874 23922 13938 23986
rect 13966 23922 14030 23986
rect 13506 23841 13570 23905
rect 13598 23841 13662 23905
rect 13690 23841 13754 23905
rect 13782 23841 13846 23905
rect 13874 23841 13938 23905
rect 13966 23841 14030 23905
rect 13506 23760 13570 23824
rect 13598 23760 13662 23824
rect 13690 23760 13754 23824
rect 13782 23760 13846 23824
rect 13874 23760 13938 23824
rect 13966 23760 14030 23824
rect 13506 23679 13570 23743
rect 13598 23679 13662 23743
rect 13690 23679 13754 23743
rect 13782 23679 13846 23743
rect 13874 23679 13938 23743
rect 13966 23679 14030 23743
rect 13506 23598 13570 23662
rect 13598 23598 13662 23662
rect 13690 23598 13754 23662
rect 13782 23598 13846 23662
rect 13874 23598 13938 23662
rect 13966 23598 14030 23662
rect 13506 23517 13570 23581
rect 13598 23517 13662 23581
rect 13690 23517 13754 23581
rect 13782 23517 13846 23581
rect 13874 23517 13938 23581
rect 13966 23517 14030 23581
rect 13506 23436 13570 23500
rect 13598 23436 13662 23500
rect 13690 23436 13754 23500
rect 13782 23436 13846 23500
rect 13874 23436 13938 23500
rect 13966 23436 14030 23500
rect 13506 23355 13570 23419
rect 13598 23355 13662 23419
rect 13690 23355 13754 23419
rect 13782 23355 13846 23419
rect 13874 23355 13938 23419
rect 13966 23355 14030 23419
rect 13506 23274 13570 23338
rect 13598 23274 13662 23338
rect 13690 23274 13754 23338
rect 13782 23274 13846 23338
rect 13874 23274 13938 23338
rect 13966 23274 14030 23338
rect 13506 23193 13570 23257
rect 13598 23193 13662 23257
rect 13690 23193 13754 23257
rect 13782 23193 13846 23257
rect 13874 23193 13938 23257
rect 13966 23193 14030 23257
rect 13506 23112 13570 23176
rect 13598 23112 13662 23176
rect 13690 23112 13754 23176
rect 13782 23112 13846 23176
rect 13874 23112 13938 23176
rect 13966 23112 14030 23176
rect 13506 23031 13570 23095
rect 13598 23031 13662 23095
rect 13690 23031 13754 23095
rect 13782 23031 13846 23095
rect 13874 23031 13938 23095
rect 13966 23031 14030 23095
rect 13506 22950 13570 23014
rect 13598 22950 13662 23014
rect 13690 22950 13754 23014
rect 13782 22950 13846 23014
rect 13874 22950 13938 23014
rect 13966 22950 14030 23014
rect 13506 22869 13570 22933
rect 13598 22869 13662 22933
rect 13690 22869 13754 22933
rect 13782 22869 13846 22933
rect 13874 22869 13938 22933
rect 13966 22869 14030 22933
rect 13506 22788 13570 22852
rect 13598 22788 13662 22852
rect 13690 22788 13754 22852
rect 13782 22788 13846 22852
rect 13874 22788 13938 22852
rect 13966 22788 14030 22852
rect 13506 22707 13570 22771
rect 13598 22707 13662 22771
rect 13690 22707 13754 22771
rect 13782 22707 13846 22771
rect 13874 22707 13938 22771
rect 13966 22707 14030 22771
rect 13506 22626 13570 22690
rect 13598 22626 13662 22690
rect 13690 22626 13754 22690
rect 13782 22626 13846 22690
rect 13874 22626 13938 22690
rect 13966 22626 14030 22690
rect 13506 22545 13570 22609
rect 13598 22545 13662 22609
rect 13690 22545 13754 22609
rect 13782 22545 13846 22609
rect 13874 22545 13938 22609
rect 13966 22545 14030 22609
rect 13506 22464 13570 22528
rect 13598 22464 13662 22528
rect 13690 22464 13754 22528
rect 13782 22464 13846 22528
rect 13874 22464 13938 22528
rect 13966 22464 14030 22528
rect 13506 22383 13570 22447
rect 13598 22383 13662 22447
rect 13690 22383 13754 22447
rect 13782 22383 13846 22447
rect 13874 22383 13938 22447
rect 13966 22383 14030 22447
rect 13506 22302 13570 22366
rect 13598 22302 13662 22366
rect 13690 22302 13754 22366
rect 13782 22302 13846 22366
rect 13874 22302 13938 22366
rect 13966 22302 14030 22366
rect 13506 22221 13570 22285
rect 13598 22221 13662 22285
rect 13690 22221 13754 22285
rect 13782 22221 13846 22285
rect 13874 22221 13938 22285
rect 13966 22221 14030 22285
rect 13506 22140 13570 22204
rect 13598 22140 13662 22204
rect 13690 22140 13754 22204
rect 13782 22140 13846 22204
rect 13874 22140 13938 22204
rect 13966 22140 14030 22204
rect 13506 22059 13570 22123
rect 13598 22059 13662 22123
rect 13690 22059 13754 22123
rect 13782 22059 13846 22123
rect 13874 22059 13938 22123
rect 13966 22059 14030 22123
rect 13506 21978 13570 22042
rect 13598 21978 13662 22042
rect 13690 21978 13754 22042
rect 13782 21978 13846 22042
rect 13874 21978 13938 22042
rect 13966 21978 14030 22042
rect 13506 21897 13570 21961
rect 13598 21897 13662 21961
rect 13690 21897 13754 21961
rect 13782 21897 13846 21961
rect 13874 21897 13938 21961
rect 13966 21897 14030 21961
rect 13506 21816 13570 21880
rect 13598 21816 13662 21880
rect 13690 21816 13754 21880
rect 13782 21816 13846 21880
rect 13874 21816 13938 21880
rect 13966 21816 14030 21880
rect 13506 21735 13570 21799
rect 13598 21735 13662 21799
rect 13690 21735 13754 21799
rect 13782 21735 13846 21799
rect 13874 21735 13938 21799
rect 13966 21735 14030 21799
rect 13506 21654 13570 21718
rect 13598 21654 13662 21718
rect 13690 21654 13754 21718
rect 13782 21654 13846 21718
rect 13874 21654 13938 21718
rect 13966 21654 14030 21718
rect 13506 21573 13570 21637
rect 13598 21573 13662 21637
rect 13690 21573 13754 21637
rect 13782 21573 13846 21637
rect 13874 21573 13938 21637
rect 13966 21573 14030 21637
rect 13506 21492 13570 21556
rect 13598 21492 13662 21556
rect 13690 21492 13754 21556
rect 13782 21492 13846 21556
rect 13874 21492 13938 21556
rect 13966 21492 14030 21556
rect 13506 21411 13570 21475
rect 13598 21411 13662 21475
rect 13690 21411 13754 21475
rect 13782 21411 13846 21475
rect 13874 21411 13938 21475
rect 13966 21411 14030 21475
rect 13506 21330 13570 21394
rect 13598 21330 13662 21394
rect 13690 21330 13754 21394
rect 13782 21330 13846 21394
rect 13874 21330 13938 21394
rect 13966 21330 14030 21394
rect 13506 21249 13570 21313
rect 13598 21249 13662 21313
rect 13690 21249 13754 21313
rect 13782 21249 13846 21313
rect 13874 21249 13938 21313
rect 13966 21249 14030 21313
rect 13506 21168 13570 21232
rect 13598 21168 13662 21232
rect 13690 21168 13754 21232
rect 13782 21168 13846 21232
rect 13874 21168 13938 21232
rect 13966 21168 14030 21232
rect 13506 21087 13570 21151
rect 13598 21087 13662 21151
rect 13690 21087 13754 21151
rect 13782 21087 13846 21151
rect 13874 21087 13938 21151
rect 13966 21087 14030 21151
rect 13506 21006 13570 21070
rect 13598 21006 13662 21070
rect 13690 21006 13754 21070
rect 13782 21006 13846 21070
rect 13874 21006 13938 21070
rect 13966 21006 14030 21070
rect 13506 20925 13570 20989
rect 13598 20925 13662 20989
rect 13690 20925 13754 20989
rect 13782 20925 13846 20989
rect 13874 20925 13938 20989
rect 13966 20925 14030 20989
rect 13506 20844 13570 20908
rect 13598 20844 13662 20908
rect 13690 20844 13754 20908
rect 13782 20844 13846 20908
rect 13874 20844 13938 20908
rect 13966 20844 14030 20908
rect 13506 20763 13570 20827
rect 13598 20763 13662 20827
rect 13690 20763 13754 20827
rect 13782 20763 13846 20827
rect 13874 20763 13938 20827
rect 13966 20763 14030 20827
rect 13506 20682 13570 20746
rect 13598 20682 13662 20746
rect 13690 20682 13754 20746
rect 13782 20682 13846 20746
rect 13874 20682 13938 20746
rect 13966 20682 14030 20746
rect 13506 20601 13570 20665
rect 13598 20601 13662 20665
rect 13690 20601 13754 20665
rect 13782 20601 13846 20665
rect 13874 20601 13938 20665
rect 13966 20601 14030 20665
rect 13405 20470 13469 20534
rect 13497 20470 13561 20534
rect 13589 20470 13653 20534
rect 13681 20470 13745 20534
rect 13773 20470 13837 20534
rect 13865 20470 13929 20534
rect 13957 20470 14021 20534
rect 13324 20367 13388 20431
rect 13405 20367 13469 20431
rect 13487 20367 13551 20431
rect 13569 20367 13633 20431
rect 13651 20367 13715 20431
rect 13733 20367 13797 20431
rect 13859 20351 13923 20415
rect 13182 20247 13246 20311
rect 13324 20219 13388 20283
rect 13405 20219 13469 20283
rect 13487 20219 13551 20283
rect 13569 20219 13633 20283
rect 13651 20219 13715 20283
rect 13733 20219 13797 20283
rect 13068 20139 13132 20203
rect 13149 20139 13213 20203
rect 13231 20139 13295 20203
rect 13313 20139 13377 20203
rect 13395 20139 13459 20203
rect 13477 20139 13541 20203
rect 13636 20128 13700 20192
rect 12943 20008 13007 20072
rect 13068 19991 13132 20055
rect 13149 19991 13213 20055
rect 13231 19991 13295 20055
rect 13313 19991 13377 20055
rect 13395 19991 13459 20055
rect 13477 19991 13541 20055
rect 12870 19911 12934 19975
rect 12951 19911 13015 19975
rect 13033 19911 13097 19975
rect 13115 19911 13179 19975
rect 13197 19911 13261 19975
rect 13279 19911 13343 19975
rect 13397 19889 13461 19953
rect 12728 19793 12792 19857
rect 12870 19763 12934 19827
rect 12951 19763 13015 19827
rect 13033 19763 13097 19827
rect 13115 19763 13179 19827
rect 13197 19763 13261 19827
rect 13279 19763 13343 19827
rect 12646 19678 12710 19742
rect 12727 19678 12791 19742
rect 12809 19678 12873 19742
rect 12891 19678 12955 19742
rect 12973 19678 13037 19742
rect 13055 19678 13119 19742
rect 13182 19674 13246 19738
rect 12446 19594 12510 19658
rect 12554 19594 12618 19658
rect 12446 19485 12510 19549
rect 12554 19485 12618 19549
rect 12646 19530 12710 19594
rect 12727 19530 12791 19594
rect 12809 19530 12873 19594
rect 12891 19530 12955 19594
rect 12973 19530 13037 19594
rect 13055 19530 13119 19594
rect 12646 19444 12710 19508
rect 12737 19444 12801 19508
rect 12828 19444 12892 19508
rect 12446 19376 12510 19440
rect 12554 19376 12618 19440
rect 12950 19435 13014 19499
rect 12446 19268 12510 19332
rect 12554 19268 12618 19332
rect 12646 19296 12710 19360
rect 12737 19296 12801 19360
rect 12828 19296 12892 19360
rect 12446 19160 12510 19224
rect 12554 19160 12618 19224
rect 5008 8222 5072 8286
rect 5008 8134 5072 8198
rect 5008 8046 5072 8110
rect 5008 7958 5072 8022
rect 5018 4385 5082 4449
rect 5018 4302 5082 4366
rect 5018 4220 5082 4284
rect 5018 4138 5082 4202
rect 5018 4056 5082 4120
rect 5018 3974 5082 4038
rect 5018 3892 5082 3956
rect 5018 3810 5082 3874
rect 5018 3728 5082 3792
rect 5018 3646 5082 3710
rect 5018 3564 5082 3628
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 2393 34197 2567 34198
rect 2219 34137 2370 34158
rect 2219 34073 2220 34137
rect 2284 34073 2305 34137
rect 2369 34073 2370 34137
rect 2219 34052 2370 34073
rect 2393 34133 2394 34197
rect 2458 34133 2502 34197
rect 2566 34133 2567 34197
rect 2393 34089 2567 34133
rect 2122 34051 2349 34052
rect 2122 33987 2123 34051
rect 2187 33987 2204 34051
rect 2268 33987 2284 34051
rect 2348 33987 2349 34051
rect 1997 33915 2098 33936
rect 1997 33851 1998 33915
rect 2062 33851 2098 33915
rect 2122 33933 2349 33987
rect 2122 33869 2123 33933
rect 2187 33869 2204 33933
rect 2268 33869 2284 33933
rect 2348 33869 2349 33933
rect 2122 33868 2349 33869
rect 2393 34025 2394 34089
rect 2458 34025 2502 34089
rect 2566 34025 2567 34089
rect 2393 33981 2567 34025
rect 2393 33917 2394 33981
rect 2458 33917 2502 33981
rect 2566 33917 2567 33981
rect 2393 33872 2567 33917
rect 1997 33830 2098 33851
rect 1892 33818 2367 33819
rect 1892 33754 1893 33818
rect 1957 33754 1975 33818
rect 2039 33754 2057 33818
rect 2121 33754 2139 33818
rect 2203 33754 2221 33818
rect 2285 33754 2302 33818
rect 2366 33754 2367 33818
rect 1765 33683 1866 33704
rect 1765 33619 1766 33683
rect 1830 33619 1866 33683
rect 1765 33598 1866 33619
rect 1892 33670 2367 33754
rect 2393 33808 2394 33872
rect 2458 33808 2502 33872
rect 2566 33808 2567 33872
rect 2393 33763 2567 33808
rect 2393 33699 2394 33763
rect 2458 33699 2502 33763
rect 2566 33699 2567 33763
rect 2393 33698 2567 33699
rect 12445 34197 12619 34198
rect 12445 34133 12446 34197
rect 12510 34133 12554 34197
rect 12618 34133 12619 34197
rect 12445 34089 12619 34133
rect 12445 34025 12446 34089
rect 12510 34025 12554 34089
rect 12618 34025 12619 34089
rect 12445 33981 12619 34025
rect 12445 33917 12446 33981
rect 12510 33917 12554 33981
rect 12618 33917 12619 33981
rect 12445 33872 12619 33917
rect 12445 33808 12446 33872
rect 12510 33808 12554 33872
rect 12618 33808 12619 33872
rect 12645 34045 12893 34046
rect 12645 33981 12646 34045
rect 12710 33981 12737 34045
rect 12801 33981 12828 34045
rect 12892 33981 12893 34045
rect 12645 33897 12893 33981
rect 12645 33833 12646 33897
rect 12710 33833 12737 33897
rect 12801 33833 12828 33897
rect 12892 33833 12893 33897
rect 12645 33832 12893 33833
rect 12914 33915 13015 33936
rect 12914 33851 12950 33915
rect 13014 33851 13015 33915
rect 12914 33830 13015 33851
rect 12445 33763 12619 33808
rect 12445 33699 12446 33763
rect 12510 33699 12554 33763
rect 12618 33699 12619 33763
rect 12445 33698 12619 33699
rect 12647 33800 13099 33801
rect 12647 33736 12648 33800
rect 12712 33736 12777 33800
rect 12841 33736 12906 33800
rect 12970 33736 13034 33800
rect 13098 33736 13099 33800
rect 12647 33698 13099 33736
rect 1892 33606 1893 33670
rect 1957 33606 1975 33670
rect 2039 33606 2057 33670
rect 2121 33606 2139 33670
rect 2203 33606 2221 33670
rect 2285 33606 2302 33670
rect 2366 33606 2367 33670
rect 12647 33634 12648 33698
rect 12712 33634 12777 33698
rect 12841 33634 12906 33698
rect 12970 33634 13034 33698
rect 13098 33634 13099 33698
rect 12647 33633 13099 33634
rect 13146 33683 13247 33704
rect 1892 33605 2367 33606
rect 13146 33619 13182 33683
rect 13246 33619 13247 33683
rect 13146 33598 13247 33619
rect 12869 33594 13344 33595
rect 1683 33572 2140 33573
rect 1683 33508 1684 33572
rect 1748 33508 1782 33572
rect 1846 33508 1880 33572
rect 1944 33508 1978 33572
rect 2042 33508 2075 33572
rect 2139 33508 2140 33572
rect 1550 33468 1651 33489
rect 1550 33404 1551 33468
rect 1615 33404 1651 33468
rect 1550 33383 1651 33404
rect 1683 33448 2140 33508
rect 2184 33564 2285 33585
rect 2184 33500 2220 33564
rect 2284 33500 2285 33564
rect 2184 33479 2285 33500
rect 12727 33564 12828 33585
rect 12727 33500 12728 33564
rect 12792 33500 12828 33564
rect 12727 33479 12828 33500
rect 12869 33530 12870 33594
rect 12934 33530 12951 33594
rect 13015 33530 13033 33594
rect 13097 33530 13115 33594
rect 13179 33530 13197 33594
rect 13261 33530 13279 33594
rect 13343 33530 13344 33594
rect 1683 33384 1684 33448
rect 1748 33384 1782 33448
rect 1846 33384 1880 33448
rect 1944 33384 1978 33448
rect 2042 33384 2075 33448
rect 2139 33384 2140 33448
rect 1683 33383 2140 33384
rect 12869 33446 13344 33530
rect 12869 33382 12870 33446
rect 12934 33382 12951 33446
rect 13015 33382 13033 33446
rect 13097 33382 13115 33446
rect 13179 33382 13197 33446
rect 13261 33382 13279 33446
rect 13343 33382 13344 33446
rect 13361 33468 13462 33489
rect 13361 33404 13397 33468
rect 13461 33404 13462 33468
rect 13361 33383 13462 33404
rect 12869 33381 13344 33382
rect 1470 33366 1945 33367
rect 1470 33302 1471 33366
rect 1535 33302 1553 33366
rect 1617 33302 1635 33366
rect 1699 33302 1717 33366
rect 1781 33302 1799 33366
rect 1863 33302 1880 33366
rect 1944 33302 1945 33366
rect 1311 33229 1412 33250
rect 1311 33165 1312 33229
rect 1376 33165 1412 33229
rect 1311 33144 1412 33165
rect 1470 33218 1945 33302
rect 1969 33349 2070 33370
rect 1969 33285 2005 33349
rect 2069 33285 2070 33349
rect 1969 33264 2070 33285
rect 12942 33349 13043 33370
rect 12942 33285 12943 33349
rect 13007 33285 13043 33349
rect 12942 33264 13043 33285
rect 13067 33366 13542 33367
rect 13067 33302 13068 33366
rect 13132 33302 13149 33366
rect 13213 33302 13231 33366
rect 13295 33302 13313 33366
rect 13377 33302 13395 33366
rect 13459 33302 13477 33366
rect 13541 33302 13542 33366
rect 1470 33154 1471 33218
rect 1535 33154 1553 33218
rect 1617 33154 1635 33218
rect 1699 33154 1717 33218
rect 1781 33154 1799 33218
rect 1863 33154 1880 33218
rect 1944 33154 1945 33218
rect 1470 33153 1945 33154
rect 13067 33218 13542 33302
rect 13067 33154 13068 33218
rect 13132 33154 13149 33218
rect 13213 33154 13231 33218
rect 13295 33154 13313 33218
rect 13377 33154 13395 33218
rect 13459 33154 13477 33218
rect 13541 33154 13542 33218
rect 13067 33153 13542 33154
rect 13600 33229 13701 33250
rect 13600 33165 13636 33229
rect 13700 33165 13701 33229
rect 13600 33144 13701 33165
rect 1214 33138 1689 33139
rect 1214 33074 1215 33138
rect 1279 33074 1297 33138
rect 1361 33074 1379 33138
rect 1443 33074 1461 33138
rect 1525 33074 1543 33138
rect 1607 33074 1624 33138
rect 1688 33074 1689 33138
rect 13323 33138 13798 33139
rect 1088 33006 1189 33027
rect 1088 32942 1089 33006
rect 1153 32942 1189 33006
rect 1088 32921 1189 32942
rect 1214 32990 1689 33074
rect 1730 33110 1831 33131
rect 1730 33046 1766 33110
rect 1830 33046 1831 33110
rect 1730 33025 1831 33046
rect 13181 33110 13282 33131
rect 13181 33046 13182 33110
rect 13246 33046 13282 33110
rect 13181 33025 13282 33046
rect 13323 33074 13324 33138
rect 13388 33074 13405 33138
rect 13469 33074 13487 33138
rect 13551 33074 13569 33138
rect 13633 33074 13651 33138
rect 13715 33074 13733 33138
rect 13797 33074 13798 33138
rect 1214 32926 1215 32990
rect 1279 32926 1297 32990
rect 1361 32926 1379 32990
rect 1443 32926 1461 32990
rect 1525 32926 1543 32990
rect 1607 32926 1624 32990
rect 1688 32926 1689 32990
rect 1214 32925 1689 32926
rect 13323 32990 13798 33074
rect 13323 32926 13324 32990
rect 13388 32926 13405 32990
rect 13469 32926 13487 32990
rect 13551 32926 13569 32990
rect 13633 32926 13651 32990
rect 13715 32926 13733 32990
rect 13797 32926 13798 32990
rect 13323 32925 13798 32926
rect 13823 33006 13924 33027
rect 13823 32942 13859 33006
rect 13923 32942 13924 33006
rect 13823 32921 13924 32942
rect 964 32908 1494 32909
rect 964 32844 967 32908
rect 1031 32844 1059 32908
rect 1123 32844 1151 32908
rect 1215 32844 1243 32908
rect 1307 32844 1335 32908
rect 1399 32844 1427 32908
rect 1491 32844 1494 32908
rect 964 32828 1494 32844
rect 964 32764 967 32828
rect 1031 32764 1059 32828
rect 1123 32764 1151 32828
rect 1215 32764 1243 32828
rect 1307 32764 1335 32828
rect 1399 32764 1427 32828
rect 1491 32764 1494 32828
rect 1507 32887 1608 32908
rect 1507 32823 1543 32887
rect 1607 32823 1608 32887
rect 1507 32802 1608 32823
rect 13404 32887 13505 32908
rect 13404 32823 13405 32887
rect 13469 32870 13505 32887
rect 13469 32869 14033 32870
rect 13469 32823 13506 32869
rect 13404 32805 13506 32823
rect 13570 32805 13598 32869
rect 13662 32805 13690 32869
rect 13754 32805 13782 32869
rect 13846 32805 13874 32869
rect 13938 32805 13966 32869
rect 14030 32805 14033 32869
rect 13404 32802 14033 32805
rect 964 32748 1494 32764
rect 964 32684 967 32748
rect 1031 32684 1059 32748
rect 1123 32684 1151 32748
rect 1215 32684 1243 32748
rect 1307 32684 1335 32748
rect 1399 32684 1427 32748
rect 1491 32684 1494 32748
rect 964 32668 1494 32684
rect 964 32604 967 32668
rect 1031 32604 1059 32668
rect 1123 32604 1151 32668
rect 1215 32604 1243 32668
rect 1307 32604 1335 32668
rect 1399 32604 1427 32668
rect 1491 32604 1494 32668
rect 964 32588 1494 32604
rect 964 32524 967 32588
rect 1031 32524 1059 32588
rect 1123 32524 1151 32588
rect 1215 32524 1243 32588
rect 1307 32524 1335 32588
rect 1399 32524 1427 32588
rect 1491 32524 1494 32588
rect 964 32508 1494 32524
rect 964 32444 967 32508
rect 1031 32444 1059 32508
rect 1123 32444 1151 32508
rect 1215 32444 1243 32508
rect 1307 32444 1335 32508
rect 1399 32444 1427 32508
rect 1491 32444 1494 32508
rect 964 32428 1494 32444
rect 964 32364 967 32428
rect 1031 32364 1059 32428
rect 1123 32364 1151 32428
rect 1215 32364 1243 32428
rect 1307 32364 1335 32428
rect 1399 32364 1427 32428
rect 1491 32364 1494 32428
rect 964 32348 1494 32364
rect 964 32284 967 32348
rect 1031 32284 1059 32348
rect 1123 32284 1151 32348
rect 1215 32284 1243 32348
rect 1307 32284 1335 32348
rect 1399 32284 1427 32348
rect 1491 32284 1494 32348
rect 964 32268 1494 32284
rect 964 32204 967 32268
rect 1031 32204 1059 32268
rect 1123 32204 1151 32268
rect 1215 32204 1243 32268
rect 1307 32204 1335 32268
rect 1399 32204 1427 32268
rect 1491 32204 1494 32268
rect 964 32188 1494 32204
rect 964 32124 967 32188
rect 1031 32124 1059 32188
rect 1123 32124 1151 32188
rect 1215 32124 1243 32188
rect 1307 32124 1335 32188
rect 1399 32124 1427 32188
rect 1491 32124 1494 32188
rect 964 32108 1494 32124
rect 964 32044 967 32108
rect 1031 32044 1059 32108
rect 1123 32044 1151 32108
rect 1215 32044 1243 32108
rect 1307 32044 1335 32108
rect 1399 32044 1427 32108
rect 1491 32044 1494 32108
rect 964 32028 1494 32044
rect 964 31964 967 32028
rect 1031 31964 1059 32028
rect 1123 31964 1151 32028
rect 1215 31964 1243 32028
rect 1307 31964 1335 32028
rect 1399 31964 1427 32028
rect 1491 31964 1494 32028
rect 964 31948 1494 31964
rect 964 31884 967 31948
rect 1031 31884 1059 31948
rect 1123 31884 1151 31948
rect 1215 31884 1243 31948
rect 1307 31884 1335 31948
rect 1399 31884 1427 31948
rect 1491 31884 1494 31948
rect 964 31868 1494 31884
rect 964 31804 967 31868
rect 1031 31804 1059 31868
rect 1123 31804 1151 31868
rect 1215 31804 1243 31868
rect 1307 31804 1335 31868
rect 1399 31804 1427 31868
rect 1491 31804 1494 31868
rect 964 31788 1494 31804
rect 964 31724 967 31788
rect 1031 31724 1059 31788
rect 1123 31724 1151 31788
rect 1215 31724 1243 31788
rect 1307 31724 1335 31788
rect 1399 31724 1427 31788
rect 1491 31724 1494 31788
rect 964 31708 1494 31724
rect 964 31644 967 31708
rect 1031 31644 1059 31708
rect 1123 31644 1151 31708
rect 1215 31644 1243 31708
rect 1307 31644 1335 31708
rect 1399 31644 1427 31708
rect 1491 31644 1494 31708
rect 964 31628 1494 31644
rect 964 31564 967 31628
rect 1031 31564 1059 31628
rect 1123 31564 1151 31628
rect 1215 31564 1243 31628
rect 1307 31564 1335 31628
rect 1399 31564 1427 31628
rect 1491 31564 1494 31628
rect 964 31548 1494 31564
rect 964 31484 967 31548
rect 1031 31484 1059 31548
rect 1123 31484 1151 31548
rect 1215 31484 1243 31548
rect 1307 31484 1335 31548
rect 1399 31484 1427 31548
rect 1491 31484 1494 31548
rect 964 31468 1494 31484
rect 964 31404 967 31468
rect 1031 31404 1059 31468
rect 1123 31404 1151 31468
rect 1215 31404 1243 31468
rect 1307 31404 1335 31468
rect 1399 31404 1427 31468
rect 1491 31404 1494 31468
rect 964 31388 1494 31404
rect 964 31324 967 31388
rect 1031 31324 1059 31388
rect 1123 31324 1151 31388
rect 1215 31324 1243 31388
rect 1307 31324 1335 31388
rect 1399 31324 1427 31388
rect 1491 31324 1494 31388
rect 964 31308 1494 31324
rect 964 31244 967 31308
rect 1031 31244 1059 31308
rect 1123 31244 1151 31308
rect 1215 31244 1243 31308
rect 1307 31244 1335 31308
rect 1399 31244 1427 31308
rect 1491 31244 1494 31308
rect 964 31228 1494 31244
rect 964 31164 967 31228
rect 1031 31164 1059 31228
rect 1123 31164 1151 31228
rect 1215 31164 1243 31228
rect 1307 31164 1335 31228
rect 1399 31164 1427 31228
rect 1491 31164 1494 31228
rect 964 31148 1494 31164
rect 964 31084 967 31148
rect 1031 31084 1059 31148
rect 1123 31084 1151 31148
rect 1215 31084 1243 31148
rect 1307 31084 1335 31148
rect 1399 31084 1427 31148
rect 1491 31084 1494 31148
rect 964 31068 1494 31084
rect 964 31004 967 31068
rect 1031 31004 1059 31068
rect 1123 31004 1151 31068
rect 1215 31004 1243 31068
rect 1307 31004 1335 31068
rect 1399 31004 1427 31068
rect 1491 31004 1494 31068
rect 964 30988 1494 31004
rect 964 30924 967 30988
rect 1031 30924 1059 30988
rect 1123 30924 1151 30988
rect 1215 30924 1243 30988
rect 1307 30924 1335 30988
rect 1399 30924 1427 30988
rect 1491 30924 1494 30988
rect 964 30908 1494 30924
rect 964 30844 967 30908
rect 1031 30844 1059 30908
rect 1123 30844 1151 30908
rect 1215 30844 1243 30908
rect 1307 30844 1335 30908
rect 1399 30844 1427 30908
rect 1491 30844 1494 30908
rect 964 30828 1494 30844
rect 964 30764 967 30828
rect 1031 30764 1059 30828
rect 1123 30764 1151 30828
rect 1215 30764 1243 30828
rect 1307 30764 1335 30828
rect 1399 30764 1427 30828
rect 1491 30764 1494 30828
rect 964 30748 1494 30764
rect 964 30684 967 30748
rect 1031 30684 1059 30748
rect 1123 30684 1151 30748
rect 1215 30684 1243 30748
rect 1307 30684 1335 30748
rect 1399 30684 1427 30748
rect 1491 30684 1494 30748
rect 964 30668 1494 30684
rect 964 30604 967 30668
rect 1031 30604 1059 30668
rect 1123 30604 1151 30668
rect 1215 30604 1243 30668
rect 1307 30604 1335 30668
rect 1399 30604 1427 30668
rect 1491 30604 1494 30668
rect 964 30588 1494 30604
rect 964 30524 967 30588
rect 1031 30524 1059 30588
rect 1123 30524 1151 30588
rect 1215 30524 1243 30588
rect 1307 30524 1335 30588
rect 1399 30524 1427 30588
rect 1491 30524 1494 30588
rect 964 30508 1494 30524
rect 964 30444 967 30508
rect 1031 30444 1059 30508
rect 1123 30444 1151 30508
rect 1215 30444 1243 30508
rect 1307 30444 1335 30508
rect 1399 30444 1427 30508
rect 1491 30444 1494 30508
rect 964 30428 1494 30444
rect 964 30364 967 30428
rect 1031 30364 1059 30428
rect 1123 30364 1151 30428
rect 1215 30364 1243 30428
rect 1307 30364 1335 30428
rect 1399 30364 1427 30428
rect 1491 30364 1494 30428
rect 964 30348 1494 30364
rect 964 30284 967 30348
rect 1031 30284 1059 30348
rect 1123 30284 1151 30348
rect 1215 30284 1243 30348
rect 1307 30284 1335 30348
rect 1399 30284 1427 30348
rect 1491 30284 1494 30348
rect 964 30268 1494 30284
rect 964 30204 967 30268
rect 1031 30204 1059 30268
rect 1123 30204 1151 30268
rect 1215 30204 1243 30268
rect 1307 30204 1335 30268
rect 1399 30204 1427 30268
rect 1491 30204 1494 30268
rect 964 30188 1494 30204
rect 964 30124 967 30188
rect 1031 30124 1059 30188
rect 1123 30124 1151 30188
rect 1215 30124 1243 30188
rect 1307 30124 1335 30188
rect 1399 30124 1427 30188
rect 1491 30124 1494 30188
rect 964 30108 1494 30124
rect 964 30044 967 30108
rect 1031 30044 1059 30108
rect 1123 30044 1151 30108
rect 1215 30044 1243 30108
rect 1307 30044 1335 30108
rect 1399 30044 1427 30108
rect 1491 30044 1494 30108
rect 964 30028 1494 30044
rect 964 29964 967 30028
rect 1031 29964 1059 30028
rect 1123 29964 1151 30028
rect 1215 29964 1243 30028
rect 1307 29964 1335 30028
rect 1399 29964 1427 30028
rect 1491 29964 1494 30028
rect 964 29948 1494 29964
rect 964 29884 967 29948
rect 1031 29884 1059 29948
rect 1123 29884 1151 29948
rect 1215 29884 1243 29948
rect 1307 29884 1335 29948
rect 1399 29884 1427 29948
rect 1491 29884 1494 29948
rect 964 29868 1494 29884
rect 964 29804 967 29868
rect 1031 29804 1059 29868
rect 1123 29804 1151 29868
rect 1215 29804 1243 29868
rect 1307 29804 1335 29868
rect 1399 29804 1427 29868
rect 1491 29804 1494 29868
rect 964 29788 1494 29804
rect 964 29724 967 29788
rect 1031 29724 1059 29788
rect 1123 29724 1151 29788
rect 1215 29724 1243 29788
rect 1307 29724 1335 29788
rect 1399 29724 1427 29788
rect 1491 29724 1494 29788
rect 964 29708 1494 29724
rect 964 29644 967 29708
rect 1031 29644 1059 29708
rect 1123 29644 1151 29708
rect 1215 29644 1243 29708
rect 1307 29644 1335 29708
rect 1399 29644 1427 29708
rect 1491 29644 1494 29708
rect 964 29628 1494 29644
rect 964 29564 967 29628
rect 1031 29564 1059 29628
rect 1123 29564 1151 29628
rect 1215 29564 1243 29628
rect 1307 29564 1335 29628
rect 1399 29564 1427 29628
rect 1491 29564 1494 29628
rect 964 29548 1494 29564
rect 964 29484 967 29548
rect 1031 29484 1059 29548
rect 1123 29484 1151 29548
rect 1215 29484 1243 29548
rect 1307 29484 1335 29548
rect 1399 29484 1427 29548
rect 1491 29484 1494 29548
rect 964 29468 1494 29484
rect 964 29404 967 29468
rect 1031 29404 1059 29468
rect 1123 29404 1151 29468
rect 1215 29404 1243 29468
rect 1307 29404 1335 29468
rect 1399 29404 1427 29468
rect 1491 29404 1494 29468
rect 964 29388 1494 29404
rect 964 29324 967 29388
rect 1031 29324 1059 29388
rect 1123 29324 1151 29388
rect 1215 29324 1243 29388
rect 1307 29324 1335 29388
rect 1399 29324 1427 29388
rect 1491 29324 1494 29388
rect 964 29308 1494 29324
rect 964 29244 967 29308
rect 1031 29244 1059 29308
rect 1123 29244 1151 29308
rect 1215 29244 1243 29308
rect 1307 29244 1335 29308
rect 1399 29244 1427 29308
rect 1491 29244 1494 29308
rect 964 29228 1494 29244
rect 964 29164 967 29228
rect 1031 29164 1059 29228
rect 1123 29164 1151 29228
rect 1215 29164 1243 29228
rect 1307 29164 1335 29228
rect 1399 29164 1427 29228
rect 1491 29164 1494 29228
rect 964 29148 1494 29164
rect 964 29084 967 29148
rect 1031 29084 1059 29148
rect 1123 29084 1151 29148
rect 1215 29084 1243 29148
rect 1307 29084 1335 29148
rect 1399 29084 1427 29148
rect 1491 29084 1494 29148
rect 964 29068 1494 29084
rect 964 29004 967 29068
rect 1031 29004 1059 29068
rect 1123 29004 1151 29068
rect 1215 29004 1243 29068
rect 1307 29004 1335 29068
rect 1399 29004 1427 29068
rect 1491 29004 1494 29068
rect 964 28988 1494 29004
rect 964 28924 967 28988
rect 1031 28924 1059 28988
rect 1123 28924 1151 28988
rect 1215 28924 1243 28988
rect 1307 28924 1335 28988
rect 1399 28924 1427 28988
rect 1491 28924 1494 28988
rect 964 28908 1494 28924
rect 964 28844 967 28908
rect 1031 28844 1059 28908
rect 1123 28844 1151 28908
rect 1215 28844 1243 28908
rect 1307 28844 1335 28908
rect 1399 28844 1427 28908
rect 1491 28844 1494 28908
rect 964 28828 1494 28844
rect 964 28764 967 28828
rect 1031 28764 1059 28828
rect 1123 28764 1151 28828
rect 1215 28764 1243 28828
rect 1307 28764 1335 28828
rect 1399 28764 1427 28828
rect 1491 28764 1494 28828
rect 964 28748 1494 28764
rect 964 28684 967 28748
rect 1031 28684 1059 28748
rect 1123 28684 1151 28748
rect 1215 28684 1243 28748
rect 1307 28684 1335 28748
rect 1399 28684 1427 28748
rect 1491 28684 1494 28748
rect 964 28668 1494 28684
rect 964 28604 967 28668
rect 1031 28604 1059 28668
rect 1123 28604 1151 28668
rect 1215 28604 1243 28668
rect 1307 28604 1335 28668
rect 1399 28604 1427 28668
rect 1491 28604 1494 28668
rect 964 28588 1494 28604
rect 964 28524 967 28588
rect 1031 28524 1059 28588
rect 1123 28524 1151 28588
rect 1215 28524 1243 28588
rect 1307 28524 1335 28588
rect 1399 28524 1427 28588
rect 1491 28524 1494 28588
rect 964 28508 1494 28524
rect 964 28444 967 28508
rect 1031 28444 1059 28508
rect 1123 28444 1151 28508
rect 1215 28444 1243 28508
rect 1307 28444 1335 28508
rect 1399 28444 1427 28508
rect 1491 28444 1494 28508
rect 964 28428 1494 28444
rect 964 28364 967 28428
rect 1031 28364 1059 28428
rect 1123 28364 1151 28428
rect 1215 28364 1243 28428
rect 1307 28364 1335 28428
rect 1399 28364 1427 28428
rect 1491 28364 1494 28428
rect 964 28348 1494 28364
rect 964 28284 967 28348
rect 1031 28284 1059 28348
rect 1123 28284 1151 28348
rect 1215 28284 1243 28348
rect 1307 28284 1335 28348
rect 1399 28284 1427 28348
rect 1491 28284 1494 28348
rect 964 28268 1494 28284
rect 964 28204 967 28268
rect 1031 28204 1059 28268
rect 1123 28204 1151 28268
rect 1215 28204 1243 28268
rect 1307 28204 1335 28268
rect 1399 28204 1427 28268
rect 1491 28204 1494 28268
rect 964 28188 1494 28204
rect 964 28124 967 28188
rect 1031 28124 1059 28188
rect 1123 28124 1151 28188
rect 1215 28124 1243 28188
rect 1307 28124 1335 28188
rect 1399 28124 1427 28188
rect 1491 28124 1494 28188
rect 964 28108 1494 28124
rect 964 28044 967 28108
rect 1031 28044 1059 28108
rect 1123 28044 1151 28108
rect 1215 28044 1243 28108
rect 1307 28044 1335 28108
rect 1399 28044 1427 28108
rect 1491 28044 1494 28108
rect 964 28028 1494 28044
rect 964 27964 967 28028
rect 1031 27964 1059 28028
rect 1123 27964 1151 28028
rect 1215 27964 1243 28028
rect 1307 27964 1335 28028
rect 1399 27964 1427 28028
rect 1491 27964 1494 28028
rect 964 27948 1494 27964
rect 964 27884 967 27948
rect 1031 27884 1059 27948
rect 1123 27884 1151 27948
rect 1215 27884 1243 27948
rect 1307 27884 1335 27948
rect 1399 27884 1427 27948
rect 1491 27884 1494 27948
rect 964 27868 1494 27884
rect 964 27804 967 27868
rect 1031 27804 1059 27868
rect 1123 27804 1151 27868
rect 1215 27804 1243 27868
rect 1307 27804 1335 27868
rect 1399 27804 1427 27868
rect 1491 27804 1494 27868
rect 964 27788 1494 27804
rect 964 27724 967 27788
rect 1031 27724 1059 27788
rect 1123 27724 1151 27788
rect 1215 27724 1243 27788
rect 1307 27724 1335 27788
rect 1399 27724 1427 27788
rect 1491 27724 1494 27788
rect 964 27708 1494 27724
rect 964 27644 967 27708
rect 1031 27644 1059 27708
rect 1123 27644 1151 27708
rect 1215 27644 1243 27708
rect 1307 27644 1335 27708
rect 1399 27644 1427 27708
rect 1491 27644 1494 27708
rect 964 27628 1494 27644
rect 964 27564 967 27628
rect 1031 27564 1059 27628
rect 1123 27564 1151 27628
rect 1215 27564 1243 27628
rect 1307 27564 1335 27628
rect 1399 27564 1427 27628
rect 1491 27564 1494 27628
rect 964 27548 1494 27564
rect 964 27484 967 27548
rect 1031 27484 1059 27548
rect 1123 27484 1151 27548
rect 1215 27484 1243 27548
rect 1307 27484 1335 27548
rect 1399 27484 1427 27548
rect 1491 27484 1494 27548
rect 964 27468 1494 27484
rect 964 27404 967 27468
rect 1031 27404 1059 27468
rect 1123 27404 1151 27468
rect 1215 27404 1243 27468
rect 1307 27404 1335 27468
rect 1399 27404 1427 27468
rect 1491 27404 1494 27468
rect 964 27388 1494 27404
rect 964 27324 967 27388
rect 1031 27324 1059 27388
rect 1123 27324 1151 27388
rect 1215 27324 1243 27388
rect 1307 27324 1335 27388
rect 1399 27324 1427 27388
rect 1491 27324 1494 27388
rect 964 27308 1494 27324
rect 964 27244 967 27308
rect 1031 27244 1059 27308
rect 1123 27244 1151 27308
rect 1215 27244 1243 27308
rect 1307 27244 1335 27308
rect 1399 27244 1427 27308
rect 1491 27244 1494 27308
rect 964 27228 1494 27244
rect 964 27164 967 27228
rect 1031 27164 1059 27228
rect 1123 27164 1151 27228
rect 1215 27164 1243 27228
rect 1307 27164 1335 27228
rect 1399 27164 1427 27228
rect 1491 27164 1494 27228
rect 964 27148 1494 27164
rect 964 27084 967 27148
rect 1031 27084 1059 27148
rect 1123 27084 1151 27148
rect 1215 27084 1243 27148
rect 1307 27084 1335 27148
rect 1399 27084 1427 27148
rect 1491 27084 1494 27148
rect 964 27068 1494 27084
rect 964 27004 967 27068
rect 1031 27004 1059 27068
rect 1123 27004 1151 27068
rect 1215 27004 1243 27068
rect 1307 27004 1335 27068
rect 1399 27004 1427 27068
rect 1491 27004 1494 27068
rect 964 26988 1494 27004
rect 964 26924 967 26988
rect 1031 26924 1059 26988
rect 1123 26924 1151 26988
rect 1215 26924 1243 26988
rect 1307 26924 1335 26988
rect 1399 26924 1427 26988
rect 1491 26924 1494 26988
rect 964 26908 1494 26924
rect 964 26844 967 26908
rect 1031 26844 1059 26908
rect 1123 26844 1151 26908
rect 1215 26844 1243 26908
rect 1307 26844 1335 26908
rect 1399 26844 1427 26908
rect 1491 26844 1494 26908
rect 964 26828 1494 26844
rect 964 26764 967 26828
rect 1031 26764 1059 26828
rect 1123 26764 1151 26828
rect 1215 26764 1243 26828
rect 1307 26764 1335 26828
rect 1399 26764 1427 26828
rect 1491 26764 1494 26828
rect 964 26748 1494 26764
rect 964 26684 967 26748
rect 1031 26684 1059 26748
rect 1123 26684 1151 26748
rect 1215 26684 1243 26748
rect 1307 26684 1335 26748
rect 1399 26684 1427 26748
rect 1491 26684 1494 26748
rect 964 26668 1494 26684
rect 964 26604 967 26668
rect 1031 26604 1059 26668
rect 1123 26604 1151 26668
rect 1215 26604 1243 26668
rect 1307 26604 1335 26668
rect 1399 26604 1427 26668
rect 1491 26604 1494 26668
rect 964 26588 1494 26604
rect 964 26524 967 26588
rect 1031 26524 1059 26588
rect 1123 26524 1151 26588
rect 1215 26524 1243 26588
rect 1307 26524 1335 26588
rect 1399 26524 1427 26588
rect 1491 26524 1494 26588
rect 964 26508 1494 26524
rect 964 26444 967 26508
rect 1031 26444 1059 26508
rect 1123 26444 1151 26508
rect 1215 26444 1243 26508
rect 1307 26444 1335 26508
rect 1399 26444 1427 26508
rect 1491 26444 1494 26508
rect 964 26428 1494 26444
rect 964 26364 967 26428
rect 1031 26364 1059 26428
rect 1123 26364 1151 26428
rect 1215 26364 1243 26428
rect 1307 26364 1335 26428
rect 1399 26364 1427 26428
rect 1491 26364 1494 26428
rect 964 26348 1494 26364
rect 964 26284 967 26348
rect 1031 26284 1059 26348
rect 1123 26284 1151 26348
rect 1215 26284 1243 26348
rect 1307 26284 1335 26348
rect 1399 26284 1427 26348
rect 1491 26284 1494 26348
rect 964 26268 1494 26284
rect 964 26204 967 26268
rect 1031 26204 1059 26268
rect 1123 26204 1151 26268
rect 1215 26204 1243 26268
rect 1307 26204 1335 26268
rect 1399 26204 1427 26268
rect 1491 26204 1494 26268
rect 964 26188 1494 26204
rect 964 26124 967 26188
rect 1031 26124 1059 26188
rect 1123 26124 1151 26188
rect 1215 26124 1243 26188
rect 1307 26124 1335 26188
rect 1399 26124 1427 26188
rect 1491 26124 1494 26188
rect 964 26108 1494 26124
rect 964 26044 967 26108
rect 1031 26044 1059 26108
rect 1123 26044 1151 26108
rect 1215 26044 1243 26108
rect 1307 26044 1335 26108
rect 1399 26044 1427 26108
rect 1491 26044 1494 26108
rect 964 26028 1494 26044
rect 964 25964 967 26028
rect 1031 25964 1059 26028
rect 1123 25964 1151 26028
rect 1215 25964 1243 26028
rect 1307 25964 1335 26028
rect 1399 25964 1427 26028
rect 1491 25964 1494 26028
rect 964 25948 1494 25964
rect 964 25884 967 25948
rect 1031 25884 1059 25948
rect 1123 25884 1151 25948
rect 1215 25884 1243 25948
rect 1307 25884 1335 25948
rect 1399 25884 1427 25948
rect 1491 25884 1494 25948
rect 964 25868 1494 25884
rect 964 25804 967 25868
rect 1031 25804 1059 25868
rect 1123 25804 1151 25868
rect 1215 25804 1243 25868
rect 1307 25804 1335 25868
rect 1399 25804 1427 25868
rect 1491 25804 1494 25868
rect 964 25788 1494 25804
rect 964 25724 967 25788
rect 1031 25724 1059 25788
rect 1123 25724 1151 25788
rect 1215 25724 1243 25788
rect 1307 25724 1335 25788
rect 1399 25724 1427 25788
rect 1491 25724 1494 25788
rect 964 25708 1494 25724
rect 964 25644 967 25708
rect 1031 25644 1059 25708
rect 1123 25644 1151 25708
rect 1215 25644 1243 25708
rect 1307 25644 1335 25708
rect 1399 25644 1427 25708
rect 1491 25644 1494 25708
rect 964 25628 1494 25644
rect 964 25564 967 25628
rect 1031 25564 1059 25628
rect 1123 25564 1151 25628
rect 1215 25564 1243 25628
rect 1307 25564 1335 25628
rect 1399 25564 1427 25628
rect 1491 25564 1494 25628
rect 964 25547 1494 25564
rect 964 25483 967 25547
rect 1031 25483 1059 25547
rect 1123 25483 1151 25547
rect 1215 25483 1243 25547
rect 1307 25483 1335 25547
rect 1399 25483 1427 25547
rect 1491 25483 1494 25547
rect 964 25466 1494 25483
rect 964 25402 967 25466
rect 1031 25402 1059 25466
rect 1123 25402 1151 25466
rect 1215 25402 1243 25466
rect 1307 25402 1335 25466
rect 1399 25402 1427 25466
rect 1491 25402 1494 25466
rect 964 25385 1494 25402
rect 964 25321 967 25385
rect 1031 25321 1059 25385
rect 1123 25321 1151 25385
rect 1215 25321 1243 25385
rect 1307 25321 1335 25385
rect 1399 25321 1427 25385
rect 1491 25321 1494 25385
rect 964 25304 1494 25321
rect 964 25240 967 25304
rect 1031 25240 1059 25304
rect 1123 25240 1151 25304
rect 1215 25240 1243 25304
rect 1307 25240 1335 25304
rect 1399 25240 1427 25304
rect 1491 25240 1494 25304
rect 964 25223 1494 25240
rect 964 25159 967 25223
rect 1031 25159 1059 25223
rect 1123 25159 1151 25223
rect 1215 25159 1243 25223
rect 1307 25159 1335 25223
rect 1399 25159 1427 25223
rect 1491 25159 1494 25223
rect 964 25142 1494 25159
rect 964 25078 967 25142
rect 1031 25078 1059 25142
rect 1123 25078 1151 25142
rect 1215 25078 1243 25142
rect 1307 25078 1335 25142
rect 1399 25078 1427 25142
rect 1491 25078 1494 25142
rect 964 25061 1494 25078
rect 964 24997 967 25061
rect 1031 24997 1059 25061
rect 1123 24997 1151 25061
rect 1215 24997 1243 25061
rect 1307 24997 1335 25061
rect 1399 24997 1427 25061
rect 1491 24997 1494 25061
rect 964 24980 1494 24997
rect 964 24916 967 24980
rect 1031 24916 1059 24980
rect 1123 24916 1151 24980
rect 1215 24916 1243 24980
rect 1307 24916 1335 24980
rect 1399 24916 1427 24980
rect 1491 24916 1494 24980
rect 964 24899 1494 24916
rect 964 24835 967 24899
rect 1031 24835 1059 24899
rect 1123 24835 1151 24899
rect 1215 24835 1243 24899
rect 1307 24835 1335 24899
rect 1399 24835 1427 24899
rect 1491 24835 1494 24899
rect 964 24818 1494 24835
rect 964 24754 967 24818
rect 1031 24754 1059 24818
rect 1123 24754 1151 24818
rect 1215 24754 1243 24818
rect 1307 24754 1335 24818
rect 1399 24754 1427 24818
rect 1491 24754 1494 24818
rect 964 24737 1494 24754
rect 964 24673 967 24737
rect 1031 24673 1059 24737
rect 1123 24673 1151 24737
rect 1215 24673 1243 24737
rect 1307 24673 1335 24737
rect 1399 24673 1427 24737
rect 1491 24673 1494 24737
rect 964 24656 1494 24673
rect 964 24592 967 24656
rect 1031 24592 1059 24656
rect 1123 24592 1151 24656
rect 1215 24592 1243 24656
rect 1307 24592 1335 24656
rect 1399 24592 1427 24656
rect 1491 24592 1494 24656
rect 964 24575 1494 24592
rect 964 24511 967 24575
rect 1031 24511 1059 24575
rect 1123 24511 1151 24575
rect 1215 24511 1243 24575
rect 1307 24511 1335 24575
rect 1399 24511 1427 24575
rect 1491 24511 1494 24575
rect 964 24494 1494 24511
rect 964 24430 967 24494
rect 1031 24430 1059 24494
rect 1123 24430 1151 24494
rect 1215 24430 1243 24494
rect 1307 24430 1335 24494
rect 1399 24430 1427 24494
rect 1491 24430 1494 24494
rect 964 24413 1494 24430
rect 964 24349 967 24413
rect 1031 24349 1059 24413
rect 1123 24349 1151 24413
rect 1215 24349 1243 24413
rect 1307 24349 1335 24413
rect 1399 24349 1427 24413
rect 1491 24349 1494 24413
rect 964 24332 1494 24349
rect 964 24268 967 24332
rect 1031 24268 1059 24332
rect 1123 24268 1151 24332
rect 1215 24268 1243 24332
rect 1307 24268 1335 24332
rect 1399 24268 1427 24332
rect 1491 24268 1494 24332
rect 964 24251 1494 24268
rect 964 24187 967 24251
rect 1031 24187 1059 24251
rect 1123 24187 1151 24251
rect 1215 24187 1243 24251
rect 1307 24187 1335 24251
rect 1399 24187 1427 24251
rect 1491 24187 1494 24251
rect 964 24170 1494 24187
rect 964 24106 967 24170
rect 1031 24106 1059 24170
rect 1123 24106 1151 24170
rect 1215 24106 1243 24170
rect 1307 24106 1335 24170
rect 1399 24106 1427 24170
rect 1491 24106 1494 24170
rect 964 24089 1494 24106
rect 964 24025 967 24089
rect 1031 24025 1059 24089
rect 1123 24025 1151 24089
rect 1215 24025 1243 24089
rect 1307 24025 1335 24089
rect 1399 24025 1427 24089
rect 1491 24025 1494 24089
rect 964 24008 1494 24025
rect 964 23944 967 24008
rect 1031 23944 1059 24008
rect 1123 23944 1151 24008
rect 1215 23944 1243 24008
rect 1307 23944 1335 24008
rect 1399 23944 1427 24008
rect 1491 23944 1494 24008
rect 964 23927 1494 23944
rect 964 23863 967 23927
rect 1031 23863 1059 23927
rect 1123 23863 1151 23927
rect 1215 23863 1243 23927
rect 1307 23863 1335 23927
rect 1399 23863 1427 23927
rect 1491 23863 1494 23927
rect 964 23846 1494 23863
rect 964 23782 967 23846
rect 1031 23782 1059 23846
rect 1123 23782 1151 23846
rect 1215 23782 1243 23846
rect 1307 23782 1335 23846
rect 1399 23782 1427 23846
rect 1491 23782 1494 23846
rect 964 23765 1494 23782
rect 964 23701 967 23765
rect 1031 23701 1059 23765
rect 1123 23701 1151 23765
rect 1215 23701 1243 23765
rect 1307 23701 1335 23765
rect 1399 23701 1427 23765
rect 1491 23701 1494 23765
rect 964 23684 1494 23701
rect 964 23620 967 23684
rect 1031 23620 1059 23684
rect 1123 23620 1151 23684
rect 1215 23620 1243 23684
rect 1307 23620 1335 23684
rect 1399 23620 1427 23684
rect 1491 23620 1494 23684
rect 964 23603 1494 23620
rect 964 23539 967 23603
rect 1031 23539 1059 23603
rect 1123 23539 1151 23603
rect 1215 23539 1243 23603
rect 1307 23539 1335 23603
rect 1399 23539 1427 23603
rect 1491 23539 1494 23603
rect 964 23522 1494 23539
rect 964 23458 967 23522
rect 1031 23458 1059 23522
rect 1123 23458 1151 23522
rect 1215 23458 1243 23522
rect 1307 23458 1335 23522
rect 1399 23458 1427 23522
rect 1491 23458 1494 23522
rect 964 23441 1494 23458
rect 964 23377 967 23441
rect 1031 23377 1059 23441
rect 1123 23377 1151 23441
rect 1215 23377 1243 23441
rect 1307 23377 1335 23441
rect 1399 23377 1427 23441
rect 1491 23377 1494 23441
rect 964 23360 1494 23377
rect 964 23296 967 23360
rect 1031 23296 1059 23360
rect 1123 23296 1151 23360
rect 1215 23296 1243 23360
rect 1307 23296 1335 23360
rect 1399 23296 1427 23360
rect 1491 23296 1494 23360
rect 964 23279 1494 23296
rect 964 23215 967 23279
rect 1031 23215 1059 23279
rect 1123 23215 1151 23279
rect 1215 23215 1243 23279
rect 1307 23215 1335 23279
rect 1399 23215 1427 23279
rect 1491 23215 1494 23279
rect 964 23198 1494 23215
rect 964 23134 967 23198
rect 1031 23134 1059 23198
rect 1123 23134 1151 23198
rect 1215 23134 1243 23198
rect 1307 23134 1335 23198
rect 1399 23134 1427 23198
rect 1491 23134 1494 23198
rect 964 23117 1494 23134
rect 964 23053 967 23117
rect 1031 23053 1059 23117
rect 1123 23053 1151 23117
rect 1215 23053 1243 23117
rect 1307 23053 1335 23117
rect 1399 23053 1427 23117
rect 1491 23053 1494 23117
rect 964 23036 1494 23053
rect 964 22972 967 23036
rect 1031 22972 1059 23036
rect 1123 22972 1151 23036
rect 1215 22972 1243 23036
rect 1307 22972 1335 23036
rect 1399 22972 1427 23036
rect 1491 22972 1494 23036
rect 964 22955 1494 22972
rect 964 22891 967 22955
rect 1031 22891 1059 22955
rect 1123 22891 1151 22955
rect 1215 22891 1243 22955
rect 1307 22891 1335 22955
rect 1399 22891 1427 22955
rect 1491 22891 1494 22955
rect 964 22874 1494 22891
rect 964 22810 967 22874
rect 1031 22810 1059 22874
rect 1123 22810 1151 22874
rect 1215 22810 1243 22874
rect 1307 22810 1335 22874
rect 1399 22810 1427 22874
rect 1491 22810 1494 22874
rect 964 22793 1494 22810
rect 964 22729 967 22793
rect 1031 22729 1059 22793
rect 1123 22729 1151 22793
rect 1215 22729 1243 22793
rect 1307 22729 1335 22793
rect 1399 22729 1427 22793
rect 1491 22729 1494 22793
rect 964 22712 1494 22729
rect 964 22648 967 22712
rect 1031 22648 1059 22712
rect 1123 22648 1151 22712
rect 1215 22648 1243 22712
rect 1307 22648 1335 22712
rect 1399 22648 1427 22712
rect 1491 22648 1494 22712
rect 964 22631 1494 22648
rect 964 22567 967 22631
rect 1031 22567 1059 22631
rect 1123 22567 1151 22631
rect 1215 22567 1243 22631
rect 1307 22567 1335 22631
rect 1399 22567 1427 22631
rect 1491 22567 1494 22631
rect 964 22550 1494 22567
rect 964 22486 967 22550
rect 1031 22486 1059 22550
rect 1123 22486 1151 22550
rect 1215 22486 1243 22550
rect 1307 22486 1335 22550
rect 1399 22486 1427 22550
rect 1491 22486 1494 22550
rect 964 22469 1494 22486
rect 964 22405 967 22469
rect 1031 22405 1059 22469
rect 1123 22405 1151 22469
rect 1215 22405 1243 22469
rect 1307 22405 1335 22469
rect 1399 22405 1427 22469
rect 1491 22405 1494 22469
rect 964 22388 1494 22405
rect 964 22324 967 22388
rect 1031 22324 1059 22388
rect 1123 22324 1151 22388
rect 1215 22324 1243 22388
rect 1307 22324 1335 22388
rect 1399 22324 1427 22388
rect 1491 22324 1494 22388
rect 964 22307 1494 22324
rect 964 22243 967 22307
rect 1031 22243 1059 22307
rect 1123 22243 1151 22307
rect 1215 22243 1243 22307
rect 1307 22243 1335 22307
rect 1399 22243 1427 22307
rect 1491 22243 1494 22307
rect 964 22226 1494 22243
rect 964 22162 967 22226
rect 1031 22162 1059 22226
rect 1123 22162 1151 22226
rect 1215 22162 1243 22226
rect 1307 22162 1335 22226
rect 1399 22162 1427 22226
rect 1491 22162 1494 22226
rect 964 22145 1494 22162
rect 964 22081 967 22145
rect 1031 22081 1059 22145
rect 1123 22081 1151 22145
rect 1215 22081 1243 22145
rect 1307 22081 1335 22145
rect 1399 22081 1427 22145
rect 1491 22081 1494 22145
rect 964 22064 1494 22081
rect 964 22000 967 22064
rect 1031 22000 1059 22064
rect 1123 22000 1151 22064
rect 1215 22000 1243 22064
rect 1307 22000 1335 22064
rect 1399 22000 1427 22064
rect 1491 22000 1494 22064
rect 964 21983 1494 22000
rect 964 21919 967 21983
rect 1031 21919 1059 21983
rect 1123 21919 1151 21983
rect 1215 21919 1243 21983
rect 1307 21919 1335 21983
rect 1399 21919 1427 21983
rect 1491 21919 1494 21983
rect 964 21902 1494 21919
rect 964 21838 967 21902
rect 1031 21838 1059 21902
rect 1123 21838 1151 21902
rect 1215 21838 1243 21902
rect 1307 21838 1335 21902
rect 1399 21838 1427 21902
rect 1491 21838 1494 21902
rect 964 21821 1494 21838
rect 964 21757 967 21821
rect 1031 21757 1059 21821
rect 1123 21757 1151 21821
rect 1215 21757 1243 21821
rect 1307 21757 1335 21821
rect 1399 21757 1427 21821
rect 1491 21757 1494 21821
rect 964 21740 1494 21757
rect 964 21676 967 21740
rect 1031 21676 1059 21740
rect 1123 21676 1151 21740
rect 1215 21676 1243 21740
rect 1307 21676 1335 21740
rect 1399 21676 1427 21740
rect 1491 21676 1494 21740
rect 964 21659 1494 21676
rect 964 21595 967 21659
rect 1031 21595 1059 21659
rect 1123 21595 1151 21659
rect 1215 21595 1243 21659
rect 1307 21595 1335 21659
rect 1399 21595 1427 21659
rect 1491 21595 1494 21659
rect 964 21578 1494 21595
rect 964 21514 967 21578
rect 1031 21514 1059 21578
rect 1123 21514 1151 21578
rect 1215 21514 1243 21578
rect 1307 21514 1335 21578
rect 1399 21514 1427 21578
rect 1491 21514 1494 21578
rect 964 21497 1494 21514
rect 964 21433 967 21497
rect 1031 21433 1059 21497
rect 1123 21433 1151 21497
rect 1215 21433 1243 21497
rect 1307 21433 1335 21497
rect 1399 21433 1427 21497
rect 1491 21433 1494 21497
rect 964 21416 1494 21433
rect 964 21352 967 21416
rect 1031 21352 1059 21416
rect 1123 21352 1151 21416
rect 1215 21352 1243 21416
rect 1307 21352 1335 21416
rect 1399 21352 1427 21416
rect 1491 21352 1494 21416
rect 964 21335 1494 21352
rect 964 21271 967 21335
rect 1031 21271 1059 21335
rect 1123 21271 1151 21335
rect 1215 21271 1243 21335
rect 1307 21271 1335 21335
rect 1399 21271 1427 21335
rect 1491 21271 1494 21335
rect 964 21254 1494 21271
rect 964 21190 967 21254
rect 1031 21190 1059 21254
rect 1123 21190 1151 21254
rect 1215 21190 1243 21254
rect 1307 21190 1335 21254
rect 1399 21190 1427 21254
rect 1491 21190 1494 21254
rect 964 21173 1494 21190
rect 964 21109 967 21173
rect 1031 21109 1059 21173
rect 1123 21109 1151 21173
rect 1215 21109 1243 21173
rect 1307 21109 1335 21173
rect 1399 21109 1427 21173
rect 1491 21109 1494 21173
rect 964 21092 1494 21109
rect 964 21028 967 21092
rect 1031 21028 1059 21092
rect 1123 21028 1151 21092
rect 1215 21028 1243 21092
rect 1307 21028 1335 21092
rect 1399 21028 1427 21092
rect 1491 21028 1494 21092
rect 964 21011 1494 21028
rect 964 20947 967 21011
rect 1031 20947 1059 21011
rect 1123 20947 1151 21011
rect 1215 20947 1243 21011
rect 1307 20947 1335 21011
rect 1399 20947 1427 21011
rect 1491 20947 1494 21011
rect 964 20930 1494 20947
rect 964 20866 967 20930
rect 1031 20866 1059 20930
rect 1123 20866 1151 20930
rect 1215 20866 1243 20930
rect 1307 20866 1335 20930
rect 1399 20866 1427 20930
rect 1491 20866 1494 20930
rect 964 20849 1494 20866
rect 964 20785 967 20849
rect 1031 20785 1059 20849
rect 1123 20785 1151 20849
rect 1215 20785 1243 20849
rect 1307 20785 1335 20849
rect 1399 20785 1427 20849
rect 1491 20785 1494 20849
rect 964 20768 1494 20785
rect 964 20704 967 20768
rect 1031 20704 1059 20768
rect 1123 20704 1151 20768
rect 1215 20704 1243 20768
rect 1307 20704 1335 20768
rect 1399 20704 1427 20768
rect 1491 20704 1494 20768
rect 964 20687 1494 20704
rect 964 20623 967 20687
rect 1031 20623 1059 20687
rect 1123 20623 1151 20687
rect 1215 20623 1243 20687
rect 1307 20623 1335 20687
rect 1399 20623 1427 20687
rect 1491 20623 1494 20687
rect 964 20606 1494 20623
rect 964 20542 967 20606
rect 1031 20542 1059 20606
rect 1123 20542 1151 20606
rect 1215 20542 1243 20606
rect 1307 20542 1335 20606
rect 1399 20542 1427 20606
rect 1491 20542 1494 20606
rect 13503 32789 14033 32802
rect 13503 32725 13506 32789
rect 13570 32725 13598 32789
rect 13662 32725 13690 32789
rect 13754 32725 13782 32789
rect 13846 32725 13874 32789
rect 13938 32725 13966 32789
rect 14030 32725 14033 32789
rect 13503 32709 14033 32725
rect 13503 32645 13506 32709
rect 13570 32645 13598 32709
rect 13662 32645 13690 32709
rect 13754 32645 13782 32709
rect 13846 32645 13874 32709
rect 13938 32645 13966 32709
rect 14030 32645 14033 32709
rect 13503 32629 14033 32645
rect 13503 32565 13506 32629
rect 13570 32565 13598 32629
rect 13662 32565 13690 32629
rect 13754 32565 13782 32629
rect 13846 32565 13874 32629
rect 13938 32565 13966 32629
rect 14030 32565 14033 32629
rect 13503 32549 14033 32565
rect 13503 32485 13506 32549
rect 13570 32485 13598 32549
rect 13662 32485 13690 32549
rect 13754 32485 13782 32549
rect 13846 32485 13874 32549
rect 13938 32485 13966 32549
rect 14030 32485 14033 32549
rect 13503 32469 14033 32485
rect 13503 32405 13506 32469
rect 13570 32405 13598 32469
rect 13662 32405 13690 32469
rect 13754 32405 13782 32469
rect 13846 32405 13874 32469
rect 13938 32405 13966 32469
rect 14030 32405 14033 32469
rect 13503 32389 14033 32405
rect 13503 32325 13506 32389
rect 13570 32325 13598 32389
rect 13662 32325 13690 32389
rect 13754 32325 13782 32389
rect 13846 32325 13874 32389
rect 13938 32325 13966 32389
rect 14030 32325 14033 32389
rect 13503 32309 14033 32325
rect 13503 32245 13506 32309
rect 13570 32245 13598 32309
rect 13662 32245 13690 32309
rect 13754 32245 13782 32309
rect 13846 32245 13874 32309
rect 13938 32245 13966 32309
rect 14030 32245 14033 32309
rect 13503 32229 14033 32245
rect 13503 32165 13506 32229
rect 13570 32165 13598 32229
rect 13662 32165 13690 32229
rect 13754 32165 13782 32229
rect 13846 32165 13874 32229
rect 13938 32165 13966 32229
rect 14030 32165 14033 32229
rect 13503 32149 14033 32165
rect 13503 32085 13506 32149
rect 13570 32085 13598 32149
rect 13662 32085 13690 32149
rect 13754 32085 13782 32149
rect 13846 32085 13874 32149
rect 13938 32085 13966 32149
rect 14030 32085 14033 32149
rect 13503 32069 14033 32085
rect 13503 32005 13506 32069
rect 13570 32005 13598 32069
rect 13662 32005 13690 32069
rect 13754 32005 13782 32069
rect 13846 32005 13874 32069
rect 13938 32005 13966 32069
rect 14030 32005 14033 32069
rect 13503 31989 14033 32005
rect 13503 31925 13506 31989
rect 13570 31925 13598 31989
rect 13662 31925 13690 31989
rect 13754 31925 13782 31989
rect 13846 31925 13874 31989
rect 13938 31925 13966 31989
rect 14030 31925 14033 31989
rect 13503 31909 14033 31925
rect 13503 31845 13506 31909
rect 13570 31845 13598 31909
rect 13662 31845 13690 31909
rect 13754 31845 13782 31909
rect 13846 31845 13874 31909
rect 13938 31845 13966 31909
rect 14030 31845 14033 31909
rect 13503 31829 14033 31845
rect 13503 31765 13506 31829
rect 13570 31765 13598 31829
rect 13662 31765 13690 31829
rect 13754 31765 13782 31829
rect 13846 31765 13874 31829
rect 13938 31765 13966 31829
rect 14030 31765 14033 31829
rect 13503 31749 14033 31765
rect 13503 31685 13506 31749
rect 13570 31685 13598 31749
rect 13662 31685 13690 31749
rect 13754 31685 13782 31749
rect 13846 31685 13874 31749
rect 13938 31685 13966 31749
rect 14030 31685 14033 31749
rect 13503 31669 14033 31685
rect 13503 31605 13506 31669
rect 13570 31605 13598 31669
rect 13662 31605 13690 31669
rect 13754 31605 13782 31669
rect 13846 31605 13874 31669
rect 13938 31605 13966 31669
rect 14030 31605 14033 31669
rect 13503 31589 14033 31605
rect 13503 31525 13506 31589
rect 13570 31525 13598 31589
rect 13662 31525 13690 31589
rect 13754 31525 13782 31589
rect 13846 31525 13874 31589
rect 13938 31525 13966 31589
rect 14030 31525 14033 31589
rect 13503 31509 14033 31525
rect 13503 31445 13506 31509
rect 13570 31445 13598 31509
rect 13662 31445 13690 31509
rect 13754 31445 13782 31509
rect 13846 31445 13874 31509
rect 13938 31445 13966 31509
rect 14030 31445 14033 31509
rect 13503 31429 14033 31445
rect 13503 31365 13506 31429
rect 13570 31365 13598 31429
rect 13662 31365 13690 31429
rect 13754 31365 13782 31429
rect 13846 31365 13874 31429
rect 13938 31365 13966 31429
rect 14030 31365 14033 31429
rect 13503 31349 14033 31365
rect 13503 31285 13506 31349
rect 13570 31285 13598 31349
rect 13662 31285 13690 31349
rect 13754 31285 13782 31349
rect 13846 31285 13874 31349
rect 13938 31285 13966 31349
rect 14030 31285 14033 31349
rect 13503 31269 14033 31285
rect 13503 31205 13506 31269
rect 13570 31205 13598 31269
rect 13662 31205 13690 31269
rect 13754 31205 13782 31269
rect 13846 31205 13874 31269
rect 13938 31205 13966 31269
rect 14030 31205 14033 31269
rect 13503 31189 14033 31205
rect 13503 31125 13506 31189
rect 13570 31125 13598 31189
rect 13662 31125 13690 31189
rect 13754 31125 13782 31189
rect 13846 31125 13874 31189
rect 13938 31125 13966 31189
rect 14030 31125 14033 31189
rect 13503 31109 14033 31125
rect 13503 31045 13506 31109
rect 13570 31045 13598 31109
rect 13662 31045 13690 31109
rect 13754 31045 13782 31109
rect 13846 31045 13874 31109
rect 13938 31045 13966 31109
rect 14030 31045 14033 31109
rect 13503 31029 14033 31045
rect 13503 30965 13506 31029
rect 13570 30965 13598 31029
rect 13662 30965 13690 31029
rect 13754 30965 13782 31029
rect 13846 30965 13874 31029
rect 13938 30965 13966 31029
rect 14030 30965 14033 31029
rect 13503 30949 14033 30965
rect 13503 30885 13506 30949
rect 13570 30885 13598 30949
rect 13662 30885 13690 30949
rect 13754 30885 13782 30949
rect 13846 30885 13874 30949
rect 13938 30885 13966 30949
rect 14030 30885 14033 30949
rect 13503 30869 14033 30885
rect 13503 30805 13506 30869
rect 13570 30805 13598 30869
rect 13662 30805 13690 30869
rect 13754 30805 13782 30869
rect 13846 30805 13874 30869
rect 13938 30805 13966 30869
rect 14030 30805 14033 30869
rect 13503 30789 14033 30805
rect 13503 30725 13506 30789
rect 13570 30725 13598 30789
rect 13662 30725 13690 30789
rect 13754 30725 13782 30789
rect 13846 30725 13874 30789
rect 13938 30725 13966 30789
rect 14030 30725 14033 30789
rect 13503 30709 14033 30725
rect 13503 30645 13506 30709
rect 13570 30645 13598 30709
rect 13662 30645 13690 30709
rect 13754 30645 13782 30709
rect 13846 30645 13874 30709
rect 13938 30645 13966 30709
rect 14030 30645 14033 30709
rect 13503 30629 14033 30645
rect 13503 30565 13506 30629
rect 13570 30565 13598 30629
rect 13662 30565 13690 30629
rect 13754 30565 13782 30629
rect 13846 30565 13874 30629
rect 13938 30565 13966 30629
rect 14030 30565 14033 30629
rect 13503 30549 14033 30565
rect 13503 30485 13506 30549
rect 13570 30485 13598 30549
rect 13662 30485 13690 30549
rect 13754 30485 13782 30549
rect 13846 30485 13874 30549
rect 13938 30485 13966 30549
rect 14030 30485 14033 30549
rect 13503 30469 14033 30485
rect 13503 30405 13506 30469
rect 13570 30405 13598 30469
rect 13662 30405 13690 30469
rect 13754 30405 13782 30469
rect 13846 30405 13874 30469
rect 13938 30405 13966 30469
rect 14030 30405 14033 30469
rect 13503 30389 14033 30405
rect 13503 30325 13506 30389
rect 13570 30325 13598 30389
rect 13662 30325 13690 30389
rect 13754 30325 13782 30389
rect 13846 30325 13874 30389
rect 13938 30325 13966 30389
rect 14030 30325 14033 30389
rect 13503 30309 14033 30325
rect 13503 30245 13506 30309
rect 13570 30245 13598 30309
rect 13662 30245 13690 30309
rect 13754 30245 13782 30309
rect 13846 30245 13874 30309
rect 13938 30245 13966 30309
rect 14030 30245 14033 30309
rect 13503 30229 14033 30245
rect 13503 30165 13506 30229
rect 13570 30165 13598 30229
rect 13662 30165 13690 30229
rect 13754 30165 13782 30229
rect 13846 30165 13874 30229
rect 13938 30165 13966 30229
rect 14030 30165 14033 30229
rect 13503 30149 14033 30165
rect 13503 30085 13506 30149
rect 13570 30085 13598 30149
rect 13662 30085 13690 30149
rect 13754 30085 13782 30149
rect 13846 30085 13874 30149
rect 13938 30085 13966 30149
rect 14030 30085 14033 30149
rect 13503 30069 14033 30085
rect 13503 30005 13506 30069
rect 13570 30005 13598 30069
rect 13662 30005 13690 30069
rect 13754 30005 13782 30069
rect 13846 30005 13874 30069
rect 13938 30005 13966 30069
rect 14030 30005 14033 30069
rect 13503 29989 14033 30005
rect 13503 29925 13506 29989
rect 13570 29925 13598 29989
rect 13662 29925 13690 29989
rect 13754 29925 13782 29989
rect 13846 29925 13874 29989
rect 13938 29925 13966 29989
rect 14030 29925 14033 29989
rect 13503 29909 14033 29925
rect 13503 29845 13506 29909
rect 13570 29845 13598 29909
rect 13662 29845 13690 29909
rect 13754 29845 13782 29909
rect 13846 29845 13874 29909
rect 13938 29845 13966 29909
rect 14030 29845 14033 29909
rect 13503 29829 14033 29845
rect 13503 29765 13506 29829
rect 13570 29765 13598 29829
rect 13662 29765 13690 29829
rect 13754 29765 13782 29829
rect 13846 29765 13874 29829
rect 13938 29765 13966 29829
rect 14030 29765 14033 29829
rect 13503 29749 14033 29765
rect 13503 29685 13506 29749
rect 13570 29685 13598 29749
rect 13662 29685 13690 29749
rect 13754 29685 13782 29749
rect 13846 29685 13874 29749
rect 13938 29685 13966 29749
rect 14030 29685 14033 29749
rect 13503 29669 14033 29685
rect 13503 29605 13506 29669
rect 13570 29605 13598 29669
rect 13662 29605 13690 29669
rect 13754 29605 13782 29669
rect 13846 29605 13874 29669
rect 13938 29605 13966 29669
rect 14030 29605 14033 29669
rect 13503 29589 14033 29605
rect 13503 29525 13506 29589
rect 13570 29525 13598 29589
rect 13662 29525 13690 29589
rect 13754 29525 13782 29589
rect 13846 29525 13874 29589
rect 13938 29525 13966 29589
rect 14030 29525 14033 29589
rect 13503 29509 14033 29525
rect 13503 29445 13506 29509
rect 13570 29445 13598 29509
rect 13662 29445 13690 29509
rect 13754 29445 13782 29509
rect 13846 29445 13874 29509
rect 13938 29445 13966 29509
rect 14030 29445 14033 29509
rect 13503 29429 14033 29445
rect 13503 29365 13506 29429
rect 13570 29365 13598 29429
rect 13662 29365 13690 29429
rect 13754 29365 13782 29429
rect 13846 29365 13874 29429
rect 13938 29365 13966 29429
rect 14030 29365 14033 29429
rect 13503 29349 14033 29365
rect 13503 29285 13506 29349
rect 13570 29285 13598 29349
rect 13662 29285 13690 29349
rect 13754 29285 13782 29349
rect 13846 29285 13874 29349
rect 13938 29285 13966 29349
rect 14030 29285 14033 29349
rect 13503 29269 14033 29285
rect 13503 29205 13506 29269
rect 13570 29205 13598 29269
rect 13662 29205 13690 29269
rect 13754 29205 13782 29269
rect 13846 29205 13874 29269
rect 13938 29205 13966 29269
rect 14030 29205 14033 29269
rect 13503 29189 14033 29205
rect 13503 29125 13506 29189
rect 13570 29125 13598 29189
rect 13662 29125 13690 29189
rect 13754 29125 13782 29189
rect 13846 29125 13874 29189
rect 13938 29125 13966 29189
rect 14030 29125 14033 29189
rect 13503 29109 14033 29125
rect 13503 29045 13506 29109
rect 13570 29045 13598 29109
rect 13662 29045 13690 29109
rect 13754 29045 13782 29109
rect 13846 29045 13874 29109
rect 13938 29045 13966 29109
rect 14030 29045 14033 29109
rect 13503 29029 14033 29045
rect 13503 28965 13506 29029
rect 13570 28965 13598 29029
rect 13662 28965 13690 29029
rect 13754 28965 13782 29029
rect 13846 28965 13874 29029
rect 13938 28965 13966 29029
rect 14030 28965 14033 29029
rect 13503 28949 14033 28965
rect 13503 28885 13506 28949
rect 13570 28885 13598 28949
rect 13662 28885 13690 28949
rect 13754 28885 13782 28949
rect 13846 28885 13874 28949
rect 13938 28885 13966 28949
rect 14030 28885 14033 28949
rect 13503 28869 14033 28885
rect 13503 28805 13506 28869
rect 13570 28805 13598 28869
rect 13662 28805 13690 28869
rect 13754 28805 13782 28869
rect 13846 28805 13874 28869
rect 13938 28805 13966 28869
rect 14030 28805 14033 28869
rect 13503 28789 14033 28805
rect 13503 28725 13506 28789
rect 13570 28725 13598 28789
rect 13662 28725 13690 28789
rect 13754 28725 13782 28789
rect 13846 28725 13874 28789
rect 13938 28725 13966 28789
rect 14030 28725 14033 28789
rect 13503 28709 14033 28725
rect 13503 28645 13506 28709
rect 13570 28645 13598 28709
rect 13662 28645 13690 28709
rect 13754 28645 13782 28709
rect 13846 28645 13874 28709
rect 13938 28645 13966 28709
rect 14030 28645 14033 28709
rect 13503 28629 14033 28645
rect 13503 28565 13506 28629
rect 13570 28565 13598 28629
rect 13662 28565 13690 28629
rect 13754 28565 13782 28629
rect 13846 28565 13874 28629
rect 13938 28565 13966 28629
rect 14030 28565 14033 28629
rect 13503 28549 14033 28565
rect 13503 28485 13506 28549
rect 13570 28485 13598 28549
rect 13662 28485 13690 28549
rect 13754 28485 13782 28549
rect 13846 28485 13874 28549
rect 13938 28485 13966 28549
rect 14030 28485 14033 28549
rect 13503 28469 14033 28485
rect 13503 28405 13506 28469
rect 13570 28405 13598 28469
rect 13662 28405 13690 28469
rect 13754 28405 13782 28469
rect 13846 28405 13874 28469
rect 13938 28405 13966 28469
rect 14030 28405 14033 28469
rect 13503 28389 14033 28405
rect 13503 28325 13506 28389
rect 13570 28325 13598 28389
rect 13662 28325 13690 28389
rect 13754 28325 13782 28389
rect 13846 28325 13874 28389
rect 13938 28325 13966 28389
rect 14030 28325 14033 28389
rect 13503 28309 14033 28325
rect 13503 28245 13506 28309
rect 13570 28245 13598 28309
rect 13662 28245 13690 28309
rect 13754 28245 13782 28309
rect 13846 28245 13874 28309
rect 13938 28245 13966 28309
rect 14030 28245 14033 28309
rect 13503 28229 14033 28245
rect 13503 28165 13506 28229
rect 13570 28165 13598 28229
rect 13662 28165 13690 28229
rect 13754 28165 13782 28229
rect 13846 28165 13874 28229
rect 13938 28165 13966 28229
rect 14030 28165 14033 28229
rect 13503 28149 14033 28165
rect 13503 28085 13506 28149
rect 13570 28085 13598 28149
rect 13662 28085 13690 28149
rect 13754 28085 13782 28149
rect 13846 28085 13874 28149
rect 13938 28085 13966 28149
rect 14030 28085 14033 28149
rect 13503 28069 14033 28085
rect 13503 28005 13506 28069
rect 13570 28005 13598 28069
rect 13662 28005 13690 28069
rect 13754 28005 13782 28069
rect 13846 28005 13874 28069
rect 13938 28005 13966 28069
rect 14030 28005 14033 28069
rect 13503 27989 14033 28005
rect 13503 27925 13506 27989
rect 13570 27925 13598 27989
rect 13662 27925 13690 27989
rect 13754 27925 13782 27989
rect 13846 27925 13874 27989
rect 13938 27925 13966 27989
rect 14030 27925 14033 27989
rect 13503 27909 14033 27925
rect 13503 27845 13506 27909
rect 13570 27845 13598 27909
rect 13662 27845 13690 27909
rect 13754 27845 13782 27909
rect 13846 27845 13874 27909
rect 13938 27845 13966 27909
rect 14030 27845 14033 27909
rect 13503 27829 14033 27845
rect 13503 27765 13506 27829
rect 13570 27765 13598 27829
rect 13662 27765 13690 27829
rect 13754 27765 13782 27829
rect 13846 27765 13874 27829
rect 13938 27765 13966 27829
rect 14030 27765 14033 27829
rect 13503 27749 14033 27765
rect 13503 27685 13506 27749
rect 13570 27685 13598 27749
rect 13662 27685 13690 27749
rect 13754 27685 13782 27749
rect 13846 27685 13874 27749
rect 13938 27685 13966 27749
rect 14030 27685 14033 27749
rect 13503 27669 14033 27685
rect 13503 27605 13506 27669
rect 13570 27605 13598 27669
rect 13662 27605 13690 27669
rect 13754 27605 13782 27669
rect 13846 27605 13874 27669
rect 13938 27605 13966 27669
rect 14030 27605 14033 27669
rect 13503 27589 14033 27605
rect 13503 27525 13506 27589
rect 13570 27525 13598 27589
rect 13662 27525 13690 27589
rect 13754 27525 13782 27589
rect 13846 27525 13874 27589
rect 13938 27525 13966 27589
rect 14030 27525 14033 27589
rect 13503 27509 14033 27525
rect 13503 27445 13506 27509
rect 13570 27445 13598 27509
rect 13662 27445 13690 27509
rect 13754 27445 13782 27509
rect 13846 27445 13874 27509
rect 13938 27445 13966 27509
rect 14030 27445 14033 27509
rect 13503 27429 14033 27445
rect 13503 27365 13506 27429
rect 13570 27365 13598 27429
rect 13662 27365 13690 27429
rect 13754 27365 13782 27429
rect 13846 27365 13874 27429
rect 13938 27365 13966 27429
rect 14030 27365 14033 27429
rect 13503 27349 14033 27365
rect 13503 27285 13506 27349
rect 13570 27285 13598 27349
rect 13662 27285 13690 27349
rect 13754 27285 13782 27349
rect 13846 27285 13874 27349
rect 13938 27285 13966 27349
rect 14030 27285 14033 27349
rect 13503 27269 14033 27285
rect 13503 27205 13506 27269
rect 13570 27205 13598 27269
rect 13662 27205 13690 27269
rect 13754 27205 13782 27269
rect 13846 27205 13874 27269
rect 13938 27205 13966 27269
rect 14030 27205 14033 27269
rect 13503 27189 14033 27205
rect 13503 27125 13506 27189
rect 13570 27125 13598 27189
rect 13662 27125 13690 27189
rect 13754 27125 13782 27189
rect 13846 27125 13874 27189
rect 13938 27125 13966 27189
rect 14030 27125 14033 27189
rect 13503 27109 14033 27125
rect 13503 27045 13506 27109
rect 13570 27045 13598 27109
rect 13662 27045 13690 27109
rect 13754 27045 13782 27109
rect 13846 27045 13874 27109
rect 13938 27045 13966 27109
rect 14030 27045 14033 27109
rect 13503 27029 14033 27045
rect 13503 26965 13506 27029
rect 13570 26965 13598 27029
rect 13662 26965 13690 27029
rect 13754 26965 13782 27029
rect 13846 26965 13874 27029
rect 13938 26965 13966 27029
rect 14030 26965 14033 27029
rect 13503 26949 14033 26965
rect 13503 26885 13506 26949
rect 13570 26885 13598 26949
rect 13662 26885 13690 26949
rect 13754 26885 13782 26949
rect 13846 26885 13874 26949
rect 13938 26885 13966 26949
rect 14030 26885 14033 26949
rect 13503 26869 14033 26885
rect 13503 26805 13506 26869
rect 13570 26805 13598 26869
rect 13662 26805 13690 26869
rect 13754 26805 13782 26869
rect 13846 26805 13874 26869
rect 13938 26805 13966 26869
rect 14030 26805 14033 26869
rect 13503 26789 14033 26805
rect 13503 26725 13506 26789
rect 13570 26725 13598 26789
rect 13662 26725 13690 26789
rect 13754 26725 13782 26789
rect 13846 26725 13874 26789
rect 13938 26725 13966 26789
rect 14030 26725 14033 26789
rect 13503 26709 14033 26725
rect 13503 26645 13506 26709
rect 13570 26645 13598 26709
rect 13662 26645 13690 26709
rect 13754 26645 13782 26709
rect 13846 26645 13874 26709
rect 13938 26645 13966 26709
rect 14030 26645 14033 26709
rect 13503 26629 14033 26645
rect 13503 26565 13506 26629
rect 13570 26565 13598 26629
rect 13662 26565 13690 26629
rect 13754 26565 13782 26629
rect 13846 26565 13874 26629
rect 13938 26565 13966 26629
rect 14030 26565 14033 26629
rect 13503 26549 14033 26565
rect 13503 26485 13506 26549
rect 13570 26485 13598 26549
rect 13662 26485 13690 26549
rect 13754 26485 13782 26549
rect 13846 26485 13874 26549
rect 13938 26485 13966 26549
rect 14030 26485 14033 26549
rect 13503 26469 14033 26485
rect 13503 26405 13506 26469
rect 13570 26405 13598 26469
rect 13662 26405 13690 26469
rect 13754 26405 13782 26469
rect 13846 26405 13874 26469
rect 13938 26405 13966 26469
rect 14030 26405 14033 26469
rect 13503 26389 14033 26405
rect 13503 26325 13506 26389
rect 13570 26325 13598 26389
rect 13662 26325 13690 26389
rect 13754 26325 13782 26389
rect 13846 26325 13874 26389
rect 13938 26325 13966 26389
rect 14030 26325 14033 26389
rect 13503 26309 14033 26325
rect 13503 26245 13506 26309
rect 13570 26245 13598 26309
rect 13662 26245 13690 26309
rect 13754 26245 13782 26309
rect 13846 26245 13874 26309
rect 13938 26245 13966 26309
rect 14030 26245 14033 26309
rect 13503 26229 14033 26245
rect 13503 26165 13506 26229
rect 13570 26165 13598 26229
rect 13662 26165 13690 26229
rect 13754 26165 13782 26229
rect 13846 26165 13874 26229
rect 13938 26165 13966 26229
rect 14030 26165 14033 26229
rect 13503 26149 14033 26165
rect 13503 26085 13506 26149
rect 13570 26085 13598 26149
rect 13662 26085 13690 26149
rect 13754 26085 13782 26149
rect 13846 26085 13874 26149
rect 13938 26085 13966 26149
rect 14030 26085 14033 26149
rect 13503 26069 14033 26085
rect 13503 26005 13506 26069
rect 13570 26005 13598 26069
rect 13662 26005 13690 26069
rect 13754 26005 13782 26069
rect 13846 26005 13874 26069
rect 13938 26005 13966 26069
rect 14030 26005 14033 26069
rect 13503 25989 14033 26005
rect 13503 25925 13506 25989
rect 13570 25925 13598 25989
rect 13662 25925 13690 25989
rect 13754 25925 13782 25989
rect 13846 25925 13874 25989
rect 13938 25925 13966 25989
rect 14030 25925 14033 25989
rect 13503 25909 14033 25925
rect 13503 25845 13506 25909
rect 13570 25845 13598 25909
rect 13662 25845 13690 25909
rect 13754 25845 13782 25909
rect 13846 25845 13874 25909
rect 13938 25845 13966 25909
rect 14030 25845 14033 25909
rect 13503 25829 14033 25845
rect 13503 25765 13506 25829
rect 13570 25765 13598 25829
rect 13662 25765 13690 25829
rect 13754 25765 13782 25829
rect 13846 25765 13874 25829
rect 13938 25765 13966 25829
rect 14030 25765 14033 25829
rect 13503 25749 14033 25765
rect 13503 25685 13506 25749
rect 13570 25685 13598 25749
rect 13662 25685 13690 25749
rect 13754 25685 13782 25749
rect 13846 25685 13874 25749
rect 13938 25685 13966 25749
rect 14030 25685 14033 25749
rect 13503 25669 14033 25685
rect 13503 25605 13506 25669
rect 13570 25605 13598 25669
rect 13662 25605 13690 25669
rect 13754 25605 13782 25669
rect 13846 25605 13874 25669
rect 13938 25605 13966 25669
rect 14030 25605 14033 25669
rect 13503 25589 14033 25605
rect 13503 25525 13506 25589
rect 13570 25525 13598 25589
rect 13662 25525 13690 25589
rect 13754 25525 13782 25589
rect 13846 25525 13874 25589
rect 13938 25525 13966 25589
rect 14030 25525 14033 25589
rect 13503 25509 14033 25525
rect 13503 25445 13506 25509
rect 13570 25445 13598 25509
rect 13662 25445 13690 25509
rect 13754 25445 13782 25509
rect 13846 25445 13874 25509
rect 13938 25445 13966 25509
rect 14030 25445 14033 25509
rect 13503 25429 14033 25445
rect 13503 25365 13506 25429
rect 13570 25365 13598 25429
rect 13662 25365 13690 25429
rect 13754 25365 13782 25429
rect 13846 25365 13874 25429
rect 13938 25365 13966 25429
rect 14030 25365 14033 25429
rect 13503 25349 14033 25365
rect 13503 25285 13506 25349
rect 13570 25285 13598 25349
rect 13662 25285 13690 25349
rect 13754 25285 13782 25349
rect 13846 25285 13874 25349
rect 13938 25285 13966 25349
rect 14030 25285 14033 25349
rect 13503 25269 14033 25285
rect 13503 25205 13506 25269
rect 13570 25205 13598 25269
rect 13662 25205 13690 25269
rect 13754 25205 13782 25269
rect 13846 25205 13874 25269
rect 13938 25205 13966 25269
rect 14030 25205 14033 25269
rect 13503 25189 14033 25205
rect 13503 25125 13506 25189
rect 13570 25125 13598 25189
rect 13662 25125 13690 25189
rect 13754 25125 13782 25189
rect 13846 25125 13874 25189
rect 13938 25125 13966 25189
rect 14030 25125 14033 25189
rect 13503 25109 14033 25125
rect 13503 25045 13506 25109
rect 13570 25045 13598 25109
rect 13662 25045 13690 25109
rect 13754 25045 13782 25109
rect 13846 25045 13874 25109
rect 13938 25045 13966 25109
rect 14030 25045 14033 25109
rect 13503 25029 14033 25045
rect 13503 24965 13506 25029
rect 13570 24965 13598 25029
rect 13662 24965 13690 25029
rect 13754 24965 13782 25029
rect 13846 24965 13874 25029
rect 13938 24965 13966 25029
rect 14030 24965 14033 25029
rect 13503 24949 14033 24965
rect 13503 24885 13506 24949
rect 13570 24885 13598 24949
rect 13662 24885 13690 24949
rect 13754 24885 13782 24949
rect 13846 24885 13874 24949
rect 13938 24885 13966 24949
rect 14030 24885 14033 24949
rect 13503 24869 14033 24885
rect 13503 24805 13506 24869
rect 13570 24805 13598 24869
rect 13662 24805 13690 24869
rect 13754 24805 13782 24869
rect 13846 24805 13874 24869
rect 13938 24805 13966 24869
rect 14030 24805 14033 24869
rect 13503 24789 14033 24805
rect 13503 24725 13506 24789
rect 13570 24725 13598 24789
rect 13662 24725 13690 24789
rect 13754 24725 13782 24789
rect 13846 24725 13874 24789
rect 13938 24725 13966 24789
rect 14030 24725 14033 24789
rect 13503 24709 14033 24725
rect 13503 24645 13506 24709
rect 13570 24645 13598 24709
rect 13662 24645 13690 24709
rect 13754 24645 13782 24709
rect 13846 24645 13874 24709
rect 13938 24645 13966 24709
rect 14030 24645 14033 24709
rect 13503 24629 14033 24645
rect 13503 24565 13506 24629
rect 13570 24565 13598 24629
rect 13662 24565 13690 24629
rect 13754 24565 13782 24629
rect 13846 24565 13874 24629
rect 13938 24565 13966 24629
rect 14030 24565 14033 24629
rect 13503 24549 14033 24565
rect 13503 24485 13506 24549
rect 13570 24485 13598 24549
rect 13662 24485 13690 24549
rect 13754 24485 13782 24549
rect 13846 24485 13874 24549
rect 13938 24485 13966 24549
rect 14030 24485 14033 24549
rect 13503 24469 14033 24485
rect 13503 24405 13506 24469
rect 13570 24405 13598 24469
rect 13662 24405 13690 24469
rect 13754 24405 13782 24469
rect 13846 24405 13874 24469
rect 13938 24405 13966 24469
rect 14030 24405 14033 24469
rect 13503 24389 14033 24405
rect 13503 24325 13506 24389
rect 13570 24325 13598 24389
rect 13662 24325 13690 24389
rect 13754 24325 13782 24389
rect 13846 24325 13874 24389
rect 13938 24325 13966 24389
rect 14030 24325 14033 24389
rect 13503 24309 14033 24325
rect 13503 24245 13506 24309
rect 13570 24245 13598 24309
rect 13662 24245 13690 24309
rect 13754 24245 13782 24309
rect 13846 24245 13874 24309
rect 13938 24245 13966 24309
rect 14030 24245 14033 24309
rect 13503 24229 14033 24245
rect 13503 24165 13506 24229
rect 13570 24165 13598 24229
rect 13662 24165 13690 24229
rect 13754 24165 13782 24229
rect 13846 24165 13874 24229
rect 13938 24165 13966 24229
rect 14030 24165 14033 24229
rect 13503 24148 14033 24165
rect 13503 24084 13506 24148
rect 13570 24084 13598 24148
rect 13662 24084 13690 24148
rect 13754 24084 13782 24148
rect 13846 24084 13874 24148
rect 13938 24084 13966 24148
rect 14030 24084 14033 24148
rect 13503 24067 14033 24084
rect 13503 24003 13506 24067
rect 13570 24003 13598 24067
rect 13662 24003 13690 24067
rect 13754 24003 13782 24067
rect 13846 24003 13874 24067
rect 13938 24003 13966 24067
rect 14030 24003 14033 24067
rect 13503 23986 14033 24003
rect 13503 23922 13506 23986
rect 13570 23922 13598 23986
rect 13662 23922 13690 23986
rect 13754 23922 13782 23986
rect 13846 23922 13874 23986
rect 13938 23922 13966 23986
rect 14030 23922 14033 23986
rect 13503 23905 14033 23922
rect 13503 23841 13506 23905
rect 13570 23841 13598 23905
rect 13662 23841 13690 23905
rect 13754 23841 13782 23905
rect 13846 23841 13874 23905
rect 13938 23841 13966 23905
rect 14030 23841 14033 23905
rect 13503 23824 14033 23841
rect 13503 23760 13506 23824
rect 13570 23760 13598 23824
rect 13662 23760 13690 23824
rect 13754 23760 13782 23824
rect 13846 23760 13874 23824
rect 13938 23760 13966 23824
rect 14030 23760 14033 23824
rect 13503 23743 14033 23760
rect 13503 23679 13506 23743
rect 13570 23679 13598 23743
rect 13662 23679 13690 23743
rect 13754 23679 13782 23743
rect 13846 23679 13874 23743
rect 13938 23679 13966 23743
rect 14030 23679 14033 23743
rect 13503 23662 14033 23679
rect 13503 23598 13506 23662
rect 13570 23598 13598 23662
rect 13662 23598 13690 23662
rect 13754 23598 13782 23662
rect 13846 23598 13874 23662
rect 13938 23598 13966 23662
rect 14030 23598 14033 23662
rect 13503 23581 14033 23598
rect 13503 23517 13506 23581
rect 13570 23517 13598 23581
rect 13662 23517 13690 23581
rect 13754 23517 13782 23581
rect 13846 23517 13874 23581
rect 13938 23517 13966 23581
rect 14030 23517 14033 23581
rect 13503 23500 14033 23517
rect 13503 23436 13506 23500
rect 13570 23436 13598 23500
rect 13662 23436 13690 23500
rect 13754 23436 13782 23500
rect 13846 23436 13874 23500
rect 13938 23436 13966 23500
rect 14030 23436 14033 23500
rect 13503 23419 14033 23436
rect 13503 23355 13506 23419
rect 13570 23355 13598 23419
rect 13662 23355 13690 23419
rect 13754 23355 13782 23419
rect 13846 23355 13874 23419
rect 13938 23355 13966 23419
rect 14030 23355 14033 23419
rect 13503 23338 14033 23355
rect 13503 23274 13506 23338
rect 13570 23274 13598 23338
rect 13662 23274 13690 23338
rect 13754 23274 13782 23338
rect 13846 23274 13874 23338
rect 13938 23274 13966 23338
rect 14030 23274 14033 23338
rect 13503 23257 14033 23274
rect 13503 23193 13506 23257
rect 13570 23193 13598 23257
rect 13662 23193 13690 23257
rect 13754 23193 13782 23257
rect 13846 23193 13874 23257
rect 13938 23193 13966 23257
rect 14030 23193 14033 23257
rect 13503 23176 14033 23193
rect 13503 23112 13506 23176
rect 13570 23112 13598 23176
rect 13662 23112 13690 23176
rect 13754 23112 13782 23176
rect 13846 23112 13874 23176
rect 13938 23112 13966 23176
rect 14030 23112 14033 23176
rect 13503 23095 14033 23112
rect 13503 23031 13506 23095
rect 13570 23031 13598 23095
rect 13662 23031 13690 23095
rect 13754 23031 13782 23095
rect 13846 23031 13874 23095
rect 13938 23031 13966 23095
rect 14030 23031 14033 23095
rect 13503 23014 14033 23031
rect 13503 22950 13506 23014
rect 13570 22950 13598 23014
rect 13662 22950 13690 23014
rect 13754 22950 13782 23014
rect 13846 22950 13874 23014
rect 13938 22950 13966 23014
rect 14030 22950 14033 23014
rect 13503 22933 14033 22950
rect 13503 22869 13506 22933
rect 13570 22869 13598 22933
rect 13662 22869 13690 22933
rect 13754 22869 13782 22933
rect 13846 22869 13874 22933
rect 13938 22869 13966 22933
rect 14030 22869 14033 22933
rect 13503 22852 14033 22869
rect 13503 22788 13506 22852
rect 13570 22788 13598 22852
rect 13662 22788 13690 22852
rect 13754 22788 13782 22852
rect 13846 22788 13874 22852
rect 13938 22788 13966 22852
rect 14030 22788 14033 22852
rect 13503 22771 14033 22788
rect 13503 22707 13506 22771
rect 13570 22707 13598 22771
rect 13662 22707 13690 22771
rect 13754 22707 13782 22771
rect 13846 22707 13874 22771
rect 13938 22707 13966 22771
rect 14030 22707 14033 22771
rect 13503 22690 14033 22707
rect 13503 22626 13506 22690
rect 13570 22626 13598 22690
rect 13662 22626 13690 22690
rect 13754 22626 13782 22690
rect 13846 22626 13874 22690
rect 13938 22626 13966 22690
rect 14030 22626 14033 22690
rect 13503 22609 14033 22626
rect 13503 22545 13506 22609
rect 13570 22545 13598 22609
rect 13662 22545 13690 22609
rect 13754 22545 13782 22609
rect 13846 22545 13874 22609
rect 13938 22545 13966 22609
rect 14030 22545 14033 22609
rect 13503 22528 14033 22545
rect 13503 22464 13506 22528
rect 13570 22464 13598 22528
rect 13662 22464 13690 22528
rect 13754 22464 13782 22528
rect 13846 22464 13874 22528
rect 13938 22464 13966 22528
rect 14030 22464 14033 22528
rect 13503 22447 14033 22464
rect 13503 22383 13506 22447
rect 13570 22383 13598 22447
rect 13662 22383 13690 22447
rect 13754 22383 13782 22447
rect 13846 22383 13874 22447
rect 13938 22383 13966 22447
rect 14030 22383 14033 22447
rect 13503 22366 14033 22383
rect 13503 22302 13506 22366
rect 13570 22302 13598 22366
rect 13662 22302 13690 22366
rect 13754 22302 13782 22366
rect 13846 22302 13874 22366
rect 13938 22302 13966 22366
rect 14030 22302 14033 22366
rect 13503 22285 14033 22302
rect 13503 22221 13506 22285
rect 13570 22221 13598 22285
rect 13662 22221 13690 22285
rect 13754 22221 13782 22285
rect 13846 22221 13874 22285
rect 13938 22221 13966 22285
rect 14030 22221 14033 22285
rect 13503 22204 14033 22221
rect 13503 22140 13506 22204
rect 13570 22140 13598 22204
rect 13662 22140 13690 22204
rect 13754 22140 13782 22204
rect 13846 22140 13874 22204
rect 13938 22140 13966 22204
rect 14030 22140 14033 22204
rect 13503 22123 14033 22140
rect 13503 22059 13506 22123
rect 13570 22059 13598 22123
rect 13662 22059 13690 22123
rect 13754 22059 13782 22123
rect 13846 22059 13874 22123
rect 13938 22059 13966 22123
rect 14030 22059 14033 22123
rect 13503 22042 14033 22059
rect 13503 21978 13506 22042
rect 13570 21978 13598 22042
rect 13662 21978 13690 22042
rect 13754 21978 13782 22042
rect 13846 21978 13874 22042
rect 13938 21978 13966 22042
rect 14030 21978 14033 22042
rect 13503 21961 14033 21978
rect 13503 21897 13506 21961
rect 13570 21897 13598 21961
rect 13662 21897 13690 21961
rect 13754 21897 13782 21961
rect 13846 21897 13874 21961
rect 13938 21897 13966 21961
rect 14030 21897 14033 21961
rect 13503 21880 14033 21897
rect 13503 21816 13506 21880
rect 13570 21816 13598 21880
rect 13662 21816 13690 21880
rect 13754 21816 13782 21880
rect 13846 21816 13874 21880
rect 13938 21816 13966 21880
rect 14030 21816 14033 21880
rect 13503 21799 14033 21816
rect 13503 21735 13506 21799
rect 13570 21735 13598 21799
rect 13662 21735 13690 21799
rect 13754 21735 13782 21799
rect 13846 21735 13874 21799
rect 13938 21735 13966 21799
rect 14030 21735 14033 21799
rect 13503 21718 14033 21735
rect 13503 21654 13506 21718
rect 13570 21654 13598 21718
rect 13662 21654 13690 21718
rect 13754 21654 13782 21718
rect 13846 21654 13874 21718
rect 13938 21654 13966 21718
rect 14030 21654 14033 21718
rect 13503 21637 14033 21654
rect 13503 21573 13506 21637
rect 13570 21573 13598 21637
rect 13662 21573 13690 21637
rect 13754 21573 13782 21637
rect 13846 21573 13874 21637
rect 13938 21573 13966 21637
rect 14030 21573 14033 21637
rect 13503 21556 14033 21573
rect 13503 21492 13506 21556
rect 13570 21492 13598 21556
rect 13662 21492 13690 21556
rect 13754 21492 13782 21556
rect 13846 21492 13874 21556
rect 13938 21492 13966 21556
rect 14030 21492 14033 21556
rect 13503 21475 14033 21492
rect 13503 21411 13506 21475
rect 13570 21411 13598 21475
rect 13662 21411 13690 21475
rect 13754 21411 13782 21475
rect 13846 21411 13874 21475
rect 13938 21411 13966 21475
rect 14030 21411 14033 21475
rect 13503 21394 14033 21411
rect 13503 21330 13506 21394
rect 13570 21330 13598 21394
rect 13662 21330 13690 21394
rect 13754 21330 13782 21394
rect 13846 21330 13874 21394
rect 13938 21330 13966 21394
rect 14030 21330 14033 21394
rect 13503 21313 14033 21330
rect 13503 21249 13506 21313
rect 13570 21249 13598 21313
rect 13662 21249 13690 21313
rect 13754 21249 13782 21313
rect 13846 21249 13874 21313
rect 13938 21249 13966 21313
rect 14030 21249 14033 21313
rect 13503 21232 14033 21249
rect 13503 21168 13506 21232
rect 13570 21168 13598 21232
rect 13662 21168 13690 21232
rect 13754 21168 13782 21232
rect 13846 21168 13874 21232
rect 13938 21168 13966 21232
rect 14030 21168 14033 21232
rect 13503 21151 14033 21168
rect 13503 21087 13506 21151
rect 13570 21087 13598 21151
rect 13662 21087 13690 21151
rect 13754 21087 13782 21151
rect 13846 21087 13874 21151
rect 13938 21087 13966 21151
rect 14030 21087 14033 21151
rect 13503 21070 14033 21087
rect 13503 21006 13506 21070
rect 13570 21006 13598 21070
rect 13662 21006 13690 21070
rect 13754 21006 13782 21070
rect 13846 21006 13874 21070
rect 13938 21006 13966 21070
rect 14030 21006 14033 21070
rect 13503 20989 14033 21006
rect 13503 20925 13506 20989
rect 13570 20925 13598 20989
rect 13662 20925 13690 20989
rect 13754 20925 13782 20989
rect 13846 20925 13874 20989
rect 13938 20925 13966 20989
rect 14030 20925 14033 20989
rect 13503 20908 14033 20925
rect 13503 20844 13506 20908
rect 13570 20844 13598 20908
rect 13662 20844 13690 20908
rect 13754 20844 13782 20908
rect 13846 20844 13874 20908
rect 13938 20844 13966 20908
rect 14030 20844 14033 20908
rect 13503 20827 14033 20844
rect 13503 20763 13506 20827
rect 13570 20763 13598 20827
rect 13662 20763 13690 20827
rect 13754 20763 13782 20827
rect 13846 20763 13874 20827
rect 13938 20763 13966 20827
rect 14030 20763 14033 20827
rect 13503 20746 14033 20763
rect 13503 20682 13506 20746
rect 13570 20682 13598 20746
rect 13662 20682 13690 20746
rect 13754 20682 13782 20746
rect 13846 20682 13874 20746
rect 13938 20682 13966 20746
rect 14030 20682 14033 20746
rect 13503 20665 14033 20682
rect 13503 20601 13506 20665
rect 13570 20601 13598 20665
rect 13662 20601 13690 20665
rect 13754 20601 13782 20665
rect 13846 20601 13874 20665
rect 13938 20601 13966 20665
rect 14030 20601 14033 20665
rect 13503 20600 14033 20601
rect 964 20525 1494 20542
rect 964 20461 967 20525
rect 1031 20461 1059 20525
rect 1123 20461 1151 20525
rect 1215 20461 1243 20525
rect 1307 20461 1335 20525
rect 1399 20461 1427 20525
rect 1491 20461 1494 20525
rect 964 20460 1494 20461
rect 1507 20534 1608 20555
rect 1507 20470 1543 20534
rect 1607 20470 1608 20534
rect 1507 20449 1608 20470
rect 13404 20534 14022 20555
rect 13404 20470 13405 20534
rect 13469 20470 13497 20534
rect 13561 20470 13589 20534
rect 13653 20470 13681 20534
rect 13745 20470 13773 20534
rect 13837 20470 13865 20534
rect 13929 20470 13957 20534
rect 14021 20470 14022 20534
rect 13404 20449 14022 20470
rect 1088 20415 1189 20436
rect 1088 20351 1089 20415
rect 1153 20351 1189 20415
rect 1088 20330 1189 20351
rect 1214 20431 1689 20432
rect 1214 20367 1215 20431
rect 1279 20367 1297 20431
rect 1361 20367 1379 20431
rect 1443 20367 1461 20431
rect 1525 20367 1543 20431
rect 1607 20367 1624 20431
rect 1688 20367 1689 20431
rect 1214 20283 1689 20367
rect 13323 20431 13798 20432
rect 13323 20367 13324 20431
rect 13388 20367 13405 20431
rect 13469 20367 13487 20431
rect 13551 20367 13569 20431
rect 13633 20367 13651 20431
rect 13715 20367 13733 20431
rect 13797 20367 13798 20431
rect 1214 20219 1215 20283
rect 1279 20219 1297 20283
rect 1361 20219 1379 20283
rect 1443 20219 1461 20283
rect 1525 20219 1543 20283
rect 1607 20219 1624 20283
rect 1688 20219 1689 20283
rect 1730 20311 1831 20332
rect 1730 20247 1766 20311
rect 1830 20247 1831 20311
rect 1730 20226 1831 20247
rect 13181 20311 13282 20332
rect 13181 20247 13182 20311
rect 13246 20247 13282 20311
rect 13181 20226 13282 20247
rect 13323 20283 13798 20367
rect 13823 20415 13924 20436
rect 13823 20351 13859 20415
rect 13923 20351 13924 20415
rect 13823 20330 13924 20351
rect 1214 20218 1689 20219
rect 13323 20219 13324 20283
rect 13388 20219 13405 20283
rect 13469 20219 13487 20283
rect 13551 20219 13569 20283
rect 13633 20219 13651 20283
rect 13715 20219 13733 20283
rect 13797 20219 13798 20283
rect 13323 20218 13798 20219
rect 1311 20192 1412 20213
rect 1311 20128 1312 20192
rect 1376 20128 1412 20192
rect 1311 20107 1412 20128
rect 1470 20203 1945 20204
rect 1470 20139 1471 20203
rect 1535 20139 1553 20203
rect 1617 20139 1635 20203
rect 1699 20139 1717 20203
rect 1781 20139 1799 20203
rect 1863 20139 1880 20203
rect 1944 20139 1945 20203
rect 1470 20055 1945 20139
rect 13067 20203 13542 20204
rect 13067 20139 13068 20203
rect 13132 20139 13149 20203
rect 13213 20139 13231 20203
rect 13295 20139 13313 20203
rect 13377 20139 13395 20203
rect 13459 20139 13477 20203
rect 13541 20139 13542 20203
rect 1470 19991 1471 20055
rect 1535 19991 1553 20055
rect 1617 19991 1635 20055
rect 1699 19991 1717 20055
rect 1781 19991 1799 20055
rect 1863 19991 1880 20055
rect 1944 19991 1945 20055
rect 1470 19990 1945 19991
rect 1969 20072 2070 20093
rect 1969 20008 2005 20072
rect 2069 20008 2070 20072
rect 1969 19987 2070 20008
rect 12942 20072 13043 20093
rect 12942 20008 12943 20072
rect 13007 20008 13043 20072
rect 12942 19987 13043 20008
rect 13067 20055 13542 20139
rect 13600 20192 13701 20213
rect 13600 20128 13636 20192
rect 13700 20128 13701 20192
rect 13600 20107 13701 20128
rect 13067 19991 13068 20055
rect 13132 19991 13149 20055
rect 13213 19991 13231 20055
rect 13295 19991 13313 20055
rect 13377 19991 13395 20055
rect 13459 19991 13477 20055
rect 13541 19991 13542 20055
rect 13067 19990 13542 19991
rect 1668 19975 2143 19976
rect 1550 19953 1651 19974
rect 1550 19889 1551 19953
rect 1615 19889 1651 19953
rect 1550 19868 1651 19889
rect 1668 19911 1669 19975
rect 1733 19911 1751 19975
rect 1815 19911 1833 19975
rect 1897 19911 1915 19975
rect 1979 19911 1997 19975
rect 2061 19911 2078 19975
rect 2142 19911 2143 19975
rect 1668 19827 2143 19911
rect 12869 19975 13344 19976
rect 12869 19911 12870 19975
rect 12934 19911 12951 19975
rect 13015 19911 13033 19975
rect 13097 19911 13115 19975
rect 13179 19911 13197 19975
rect 13261 19911 13279 19975
rect 13343 19911 13344 19975
rect 1668 19763 1669 19827
rect 1733 19763 1751 19827
rect 1815 19763 1833 19827
rect 1897 19763 1915 19827
rect 1979 19763 1997 19827
rect 2061 19763 2078 19827
rect 2142 19763 2143 19827
rect 2184 19857 2285 19878
rect 2184 19793 2220 19857
rect 2284 19793 2285 19857
rect 2184 19772 2285 19793
rect 12727 19857 12828 19878
rect 12727 19793 12728 19857
rect 12792 19793 12828 19857
rect 12727 19772 12828 19793
rect 12869 19827 13344 19911
rect 13361 19953 13462 19974
rect 13361 19889 13397 19953
rect 13461 19889 13462 19953
rect 13361 19868 13462 19889
rect 1668 19762 2143 19763
rect 12869 19763 12870 19827
rect 12934 19763 12951 19827
rect 13015 19763 13033 19827
rect 13097 19763 13115 19827
rect 13179 19763 13197 19827
rect 13261 19763 13279 19827
rect 13343 19763 13344 19827
rect 12869 19762 13344 19763
rect 1765 19738 1866 19759
rect 1765 19674 1766 19738
rect 1830 19674 1866 19738
rect 1765 19653 1866 19674
rect 1892 19742 2367 19743
rect 1892 19678 1893 19742
rect 1957 19678 1975 19742
rect 2039 19678 2057 19742
rect 2121 19678 2139 19742
rect 2203 19678 2221 19742
rect 2285 19678 2302 19742
rect 2366 19678 2367 19742
rect 1892 19594 2367 19678
rect 12645 19742 13120 19743
rect 12645 19678 12646 19742
rect 12710 19678 12727 19742
rect 12791 19678 12809 19742
rect 12873 19678 12891 19742
rect 12955 19678 12973 19742
rect 13037 19678 13055 19742
rect 13119 19678 13120 19742
rect 1892 19530 1893 19594
rect 1957 19530 1975 19594
rect 2039 19530 2057 19594
rect 2121 19530 2139 19594
rect 2203 19530 2221 19594
rect 2285 19530 2302 19594
rect 2366 19530 2367 19594
rect 1892 19529 2367 19530
rect 2393 19658 2567 19659
rect 2393 19594 2394 19658
rect 2458 19594 2502 19658
rect 2566 19594 2567 19658
rect 2393 19549 2567 19594
rect 1997 19499 2098 19520
rect 1997 19435 1998 19499
rect 2062 19435 2098 19499
rect 1997 19414 2098 19435
rect 2119 19508 2367 19509
rect 2119 19444 2120 19508
rect 2184 19444 2211 19508
rect 2275 19444 2302 19508
rect 2366 19444 2367 19508
rect 2119 19360 2367 19444
rect 2119 19296 2120 19360
rect 2184 19296 2211 19360
rect 2275 19296 2302 19360
rect 2366 19296 2367 19360
rect 2393 19485 2394 19549
rect 2458 19485 2502 19549
rect 2566 19485 2567 19549
rect 2393 19440 2567 19485
rect 2393 19376 2394 19440
rect 2458 19376 2502 19440
rect 2566 19376 2567 19440
rect 2393 19332 2567 19376
rect 2119 19295 2370 19296
rect 2219 19275 2370 19295
rect 2219 19211 2220 19275
rect 2284 19211 2305 19275
rect 2369 19211 2370 19275
rect 2219 19190 2370 19211
rect 2393 19268 2394 19332
rect 2458 19268 2502 19332
rect 2566 19268 2567 19332
rect 2393 19224 2567 19268
rect 2393 19160 2394 19224
rect 2458 19160 2502 19224
rect 2566 19160 2567 19224
rect 2393 19159 2567 19160
rect 12445 19658 12619 19659
rect 12445 19594 12446 19658
rect 12510 19594 12554 19658
rect 12618 19594 12619 19658
rect 12445 19549 12619 19594
rect 12445 19485 12446 19549
rect 12510 19485 12554 19549
rect 12618 19485 12619 19549
rect 12645 19594 13120 19678
rect 13146 19738 13247 19759
rect 13146 19674 13182 19738
rect 13246 19674 13247 19738
rect 13146 19653 13247 19674
rect 12645 19530 12646 19594
rect 12710 19530 12727 19594
rect 12791 19530 12809 19594
rect 12873 19530 12891 19594
rect 12955 19530 12973 19594
rect 13037 19530 13055 19594
rect 13119 19530 13120 19594
rect 12645 19529 13120 19530
rect 12445 19440 12619 19485
rect 12445 19376 12446 19440
rect 12510 19376 12554 19440
rect 12618 19376 12619 19440
rect 12445 19332 12619 19376
rect 12445 19268 12446 19332
rect 12510 19268 12554 19332
rect 12618 19268 12619 19332
rect 12645 19508 12893 19509
rect 12645 19444 12646 19508
rect 12710 19444 12737 19508
rect 12801 19444 12828 19508
rect 12892 19444 12893 19508
rect 12645 19360 12893 19444
rect 12914 19499 13015 19520
rect 12914 19435 12950 19499
rect 13014 19435 13015 19499
rect 12914 19414 13015 19435
rect 12645 19296 12646 19360
rect 12710 19296 12737 19360
rect 12801 19296 12828 19360
rect 12892 19296 12893 19360
rect 12645 19295 12893 19296
rect 12445 19224 12619 19268
rect 12445 19160 12446 19224
rect 12510 19160 12554 19224
rect 12618 19160 12619 19224
rect 12445 19159 12619 19160
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 7917 254 8847
rect 5007 8286 5073 8287
rect 5007 8222 5008 8286
rect 5072 8222 5073 8286
rect 5007 8198 5073 8222
rect 5007 8134 5008 8198
rect 5072 8134 5073 8198
rect 5007 8110 5073 8134
rect 5007 8046 5008 8110
rect 5072 8046 5073 8110
rect 5007 8022 5073 8046
rect 5007 7958 5008 8022
rect 5072 7958 5073 8022
rect 5007 7957 5073 7958
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 5007 4449 5093 4450
rect 5007 4385 5018 4449
rect 5082 4385 5093 4449
rect 5007 4366 5093 4385
rect 5007 4302 5018 4366
rect 5082 4302 5093 4366
rect 5007 4284 5093 4302
rect 5007 4220 5018 4284
rect 5082 4220 5093 4284
rect 5007 4202 5093 4220
rect 5007 4138 5018 4202
rect 5082 4138 5093 4202
rect 5007 4120 5093 4138
rect 5007 4056 5018 4120
rect 5082 4056 5093 4120
rect 5007 4038 5093 4056
rect 5007 3974 5018 4038
rect 5082 3974 5093 4038
rect 5007 3956 5093 3974
rect 5007 3892 5018 3956
rect 5082 3892 5093 3956
rect 5007 3874 5093 3892
rect 5007 3810 5018 3874
rect 5082 3810 5093 3874
rect 5007 3792 5093 3810
rect 5007 3728 5018 3792
rect 5082 3728 5093 3792
rect 5007 3710 5093 3728
rect 5007 3646 5018 3710
rect 5082 3646 5093 3710
rect 5007 3628 5093 3646
rect 5007 3564 5018 3628
rect 5082 3564 5093 3628
rect 5007 3563 5093 3564
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 6339 32553 10468 33424
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_0
timestamp 1606744421
transform 1 0 6274 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_1
timestamp 1606744421
transform 1 0 5720 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_2
timestamp 1606744421
transform 1 0 5234 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_3
timestamp 1606744421
transform 1 0 5166 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_4
timestamp 1606744421
transform 1 0 4680 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_5
timestamp 1606744421
transform 1 0 4612 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_6
timestamp 1606744421
transform 1 0 4126 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_7
timestamp 1606744421
transform 1 0 4058 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_8
timestamp 1606744421
transform 1 0 3572 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_9
timestamp 1606744421
transform 1 0 3504 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_10
timestamp 1606744421
transform 1 0 12922 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_11
timestamp 1606744421
transform 1 0 12990 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_12
timestamp 1606744421
transform 1 0 7450 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_13
timestamp 1606744421
transform 1 0 8004 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_14
timestamp 1606744421
transform 1 0 12922 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_15
timestamp 1606744421
transform 1 0 12990 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_16
timestamp 1606744421
transform 1 0 8490 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_17
timestamp 1606744421
transform 1 0 9044 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_18
timestamp 1606744421
transform 1 0 9598 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_19
timestamp 1606744421
transform 1 0 10152 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_20
timestamp 1606744421
transform 1 0 10706 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_21
timestamp 1606744421
transform 1 0 8558 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_22
timestamp 1606744421
transform 1 0 9112 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_23
timestamp 1606744421
transform 1 0 9666 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_24
timestamp 1606744421
transform 1 0 10220 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_25
timestamp 1606744421
transform 1 0 10774 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_26
timestamp 1606744421
transform 1 0 11260 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_27
timestamp 1606744421
transform 1 0 11814 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_28
timestamp 1606744421
transform 1 0 12368 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_29
timestamp 1606744421
transform 1 0 11328 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_30
timestamp 1606744421
transform 1 0 11882 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_31
timestamp 1606744421
transform 1 0 12436 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_32
timestamp 1606744421
transform 1 0 2950 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_33
timestamp 1606744421
transform 1 0 3018 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_34
timestamp 1606744421
transform 1 0 3504 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_35
timestamp 1606744421
transform 1 0 3572 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_36
timestamp 1606744421
transform 1 0 4058 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_37
timestamp 1606744421
transform 1 0 4126 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_38
timestamp 1606744421
transform 1 0 4612 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_39
timestamp 1606744421
transform 1 0 4680 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_40
timestamp 1606744421
transform 1 0 5166 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_41
timestamp 1606744421
transform 1 0 5234 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_42
timestamp 1606744421
transform 1 0 5720 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_43
timestamp 1606744421
transform 1 0 6274 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_44
timestamp 1606744421
transform 1 0 6828 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_45
timestamp 1606744421
transform 1 0 7382 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_46
timestamp 1606744421
transform 1 0 7936 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_47
timestamp 1606744421
transform 1 0 5788 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_48
timestamp 1606744421
transform 1 0 6342 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_49
timestamp 1606744421
transform 1 0 6896 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_50
timestamp 1606744421
transform 1 0 7450 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_51
timestamp 1606744421
transform 1 0 8004 0 -1 10722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_52
timestamp 1606744421
transform 1 0 12922 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_53
timestamp 1606744421
transform 1 0 12990 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_54
timestamp 1606744421
transform 1 0 8490 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_55
timestamp 1606744421
transform 1 0 9044 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_56
timestamp 1606744421
transform 1 0 9598 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_57
timestamp 1606744421
transform 1 0 10152 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_58
timestamp 1606744421
transform 1 0 10706 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_59
timestamp 1606744421
transform 1 0 8558 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_60
timestamp 1606744421
transform 1 0 9112 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_61
timestamp 1606744421
transform 1 0 9666 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_62
timestamp 1606744421
transform 1 0 10220 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_63
timestamp 1606744421
transform 1 0 10774 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_64
timestamp 1606744421
transform 1 0 11260 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_65
timestamp 1606744421
transform 1 0 11814 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_66
timestamp 1606744421
transform 1 0 12368 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_67
timestamp 1606744421
transform 1 0 11328 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_68
timestamp 1606744421
transform 1 0 11882 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_69
timestamp 1606744421
transform 1 0 12436 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_70
timestamp 1606744421
transform 1 0 2950 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_71
timestamp 1606744421
transform 1 0 3018 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_72
timestamp 1606744421
transform 1 0 3504 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_73
timestamp 1606744421
transform 1 0 3572 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_74
timestamp 1606744421
transform 1 0 4058 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_75
timestamp 1606744421
transform 1 0 4126 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_76
timestamp 1606744421
transform 1 0 4612 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_77
timestamp 1606744421
transform 1 0 4680 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_78
timestamp 1606744421
transform 1 0 5166 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_79
timestamp 1606744421
transform 1 0 5234 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_80
timestamp 1606744421
transform 1 0 5720 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_81
timestamp 1606744421
transform 1 0 6274 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_82
timestamp 1606744421
transform 1 0 6828 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_83
timestamp 1606744421
transform 1 0 7382 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_84
timestamp 1606744421
transform 1 0 7936 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_85
timestamp 1606744421
transform 1 0 5788 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_86
timestamp 1606744421
transform 1 0 6342 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_87
timestamp 1606744421
transform 1 0 8558 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_88
timestamp 1606744421
transform 1 0 9112 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_89
timestamp 1606744421
transform 1 0 9666 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_90
timestamp 1606744421
transform 1 0 10220 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_91
timestamp 1606744421
transform 1 0 12922 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_92
timestamp 1606744421
transform 1 0 12990 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_93
timestamp 1606744421
transform 1 0 12436 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_94
timestamp 1606744421
transform 1 0 11882 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_95
timestamp 1606744421
transform 1 0 11328 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_96
timestamp 1606744421
transform 1 0 12368 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_97
timestamp 1606744421
transform 1 0 11814 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_98
timestamp 1606744421
transform 1 0 11260 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_99
timestamp 1606744421
transform 1 0 10774 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_100
timestamp 1606744421
transform 1 0 10220 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_101
timestamp 1606744421
transform 1 0 9666 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_102
timestamp 1606744421
transform 1 0 9112 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_103
timestamp 1606744421
transform 1 0 8558 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_104
timestamp 1606744421
transform 1 0 8004 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_105
timestamp 1606744421
transform 1 0 7450 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_106
timestamp 1606744421
transform 1 0 6896 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_107
timestamp 1606744421
transform 1 0 6342 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_108
timestamp 1606744421
transform 1 0 5788 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_109
timestamp 1606744421
transform 1 0 10706 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_110
timestamp 1606744421
transform 1 0 10152 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_111
timestamp 1606744421
transform 1 0 9598 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_112
timestamp 1606744421
transform 1 0 9044 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_113
timestamp 1606744421
transform 1 0 8490 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_114
timestamp 1606744421
transform 1 0 7936 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_115
timestamp 1606744421
transform 1 0 7382 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_116
timestamp 1606744421
transform 1 0 6828 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_117
timestamp 1606744421
transform 1 0 6274 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_118
timestamp 1606744421
transform 1 0 5720 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_119
timestamp 1606744421
transform 1 0 5234 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_120
timestamp 1606744421
transform 1 0 5166 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_121
timestamp 1606744421
transform 1 0 4680 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_122
timestamp 1606744421
transform 1 0 4612 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_123
timestamp 1606744421
transform 1 0 4126 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_124
timestamp 1606744421
transform 1 0 4058 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_125
timestamp 1606744421
transform 1 0 3572 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_126
timestamp 1606744421
transform 1 0 3504 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_127
timestamp 1606744421
transform 1 0 3018 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_128
timestamp 1606744421
transform 1 0 2950 0 -1 38722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_129
timestamp 1606744421
transform 1 0 7382 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_130
timestamp 1606744421
transform 1 0 7936 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_131
timestamp 1606744421
transform 1 0 8490 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_132
timestamp 1606744421
transform 1 0 10774 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_133
timestamp 1606744421
transform 1 0 7450 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_134
timestamp 1606744421
transform 1 0 2950 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_135
timestamp 1606744421
transform 1 0 3018 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_136
timestamp 1606744421
transform 1 0 3504 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_137
timestamp 1606744421
transform 1 0 3572 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_138
timestamp 1606744421
transform 1 0 4058 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_139
timestamp 1606744421
transform 1 0 4126 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_140
timestamp 1606744421
transform 1 0 4612 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_141
timestamp 1606744421
transform 1 0 4680 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_142
timestamp 1606744421
transform 1 0 5166 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_143
timestamp 1606744421
transform 1 0 5234 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_144
timestamp 1606744421
transform 1 0 5720 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_145
timestamp 1606744421
transform 1 0 6274 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_146
timestamp 1606744421
transform 1 0 6828 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_147
timestamp 1606744421
transform 1 0 7382 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_148
timestamp 1606744421
transform 1 0 5788 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_149
timestamp 1606744421
transform 1 0 6342 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_150
timestamp 1606744421
transform 1 0 6896 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_151
timestamp 1606744421
transform 1 0 12922 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_152
timestamp 1606744421
transform 1 0 12990 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_153
timestamp 1606744421
transform 1 0 8490 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_154
timestamp 1606744421
transform 1 0 9044 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_155
timestamp 1606744421
transform 1 0 9598 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_156
timestamp 1606744421
transform 1 0 10152 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_157
timestamp 1606744421
transform 1 0 10706 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_158
timestamp 1606744421
transform 1 0 8558 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_159
timestamp 1606744421
transform 1 0 9112 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_160
timestamp 1606744421
transform 1 0 9666 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_161
timestamp 1606744421
transform 1 0 10220 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_162
timestamp 1606744421
transform 1 0 10774 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_163
timestamp 1606744421
transform 1 0 11260 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_164
timestamp 1606744421
transform 1 0 11814 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_165
timestamp 1606744421
transform 1 0 12368 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_166
timestamp 1606744421
transform 1 0 11328 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_167
timestamp 1606744421
transform 1 0 11882 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_168
timestamp 1606744421
transform 1 0 12436 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_169
timestamp 1606744421
transform 1 0 7936 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_170
timestamp 1606744421
transform 1 0 8004 0 -1 8722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_171
timestamp 1606744421
transform 1 0 7450 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_172
timestamp 1606744421
transform 1 0 2950 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_173
timestamp 1606744421
transform 1 0 3018 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_174
timestamp 1606744421
transform 1 0 3504 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_175
timestamp 1606744421
transform 1 0 3572 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_176
timestamp 1606744421
transform 1 0 4058 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_177
timestamp 1606744421
transform 1 0 4126 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_178
timestamp 1606744421
transform 1 0 4612 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_179
timestamp 1606744421
transform 1 0 4680 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_180
timestamp 1606744421
transform 1 0 5166 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_181
timestamp 1606744421
transform 1 0 5234 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_182
timestamp 1606744421
transform 1 0 5720 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_183
timestamp 1606744421
transform 1 0 6274 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_184
timestamp 1606744421
transform 1 0 6828 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_185
timestamp 1606744421
transform 1 0 7382 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_186
timestamp 1606744421
transform 1 0 5788 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_187
timestamp 1606744421
transform 1 0 6342 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_188
timestamp 1606744421
transform 1 0 6896 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_189
timestamp 1606744421
transform 1 0 12922 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_190
timestamp 1606744421
transform 1 0 12990 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_191
timestamp 1606744421
transform 1 0 8490 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_192
timestamp 1606744421
transform 1 0 9044 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_193
timestamp 1606744421
transform 1 0 9598 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_194
timestamp 1606744421
transform 1 0 10152 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_195
timestamp 1606744421
transform 1 0 10706 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_196
timestamp 1606744421
transform 1 0 8558 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_197
timestamp 1606744421
transform 1 0 9112 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_198
timestamp 1606744421
transform 1 0 9666 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_199
timestamp 1606744421
transform 1 0 10220 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_200
timestamp 1606744421
transform 1 0 10774 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_201
timestamp 1606744421
transform 1 0 11260 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_202
timestamp 1606744421
transform 1 0 11814 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_203
timestamp 1606744421
transform 1 0 12368 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_204
timestamp 1606744421
transform 1 0 11328 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_205
timestamp 1606744421
transform 1 0 11882 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_206
timestamp 1606744421
transform 1 0 12436 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_207
timestamp 1606744421
transform 1 0 7936 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_208
timestamp 1606744421
transform 1 0 8004 0 -1 6722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_209
timestamp 1606744421
transform 1 0 9044 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_210
timestamp 1606744421
transform 1 0 9598 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_211
timestamp 1606744421
transform 1 0 12849 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_212
timestamp 1606744421
transform 1 0 12013 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_213
timestamp 1606744421
transform 1 0 11177 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_214
timestamp 1606744421
transform 1 0 10341 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_215
timestamp 1606744421
transform 1 0 9505 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_216
timestamp 1606744421
transform 1 0 8669 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_217
timestamp 1606744421
transform 1 0 7833 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_218
timestamp 1606744421
transform 1 0 6997 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_219
timestamp 1606744421
transform 1 0 6161 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_220
timestamp 1606744421
transform 1 0 5325 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_221
timestamp 1606744421
transform 1 0 4489 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_222
timestamp 1606744421
transform 1 0 12781 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_223
timestamp 1606744421
transform 1 0 11945 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_224
timestamp 1606744421
transform 1 0 11109 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_225
timestamp 1606744421
transform 1 0 10273 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_226
timestamp 1606744421
transform 1 0 9437 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_227
timestamp 1606744421
transform 1 0 8601 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_228
timestamp 1606744421
transform 1 0 7765 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_229
timestamp 1606744421
transform 1 0 6929 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_230
timestamp 1606744421
transform 1 0 6093 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_231
timestamp 1606744421
transform 1 0 5257 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_232
timestamp 1606744421
transform 1 0 4421 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_233
timestamp 1606744421
transform 1 0 11260 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_234
timestamp 1606744421
transform 1 0 10152 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_235
timestamp 1606744421
transform 1 0 10706 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_236
timestamp 1606744421
transform 1 0 12849 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_237
timestamp 1606744421
transform 1 0 12013 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_238
timestamp 1606744421
transform 1 0 11177 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_239
timestamp 1606744421
transform 1 0 10341 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_240
timestamp 1606744421
transform 1 0 9505 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_241
timestamp 1606744421
transform 1 0 8669 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_242
timestamp 1606744421
transform 1 0 7833 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_243
timestamp 1606744421
transform 1 0 12781 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_244
timestamp 1606744421
transform 1 0 11945 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_245
timestamp 1606744421
transform 1 0 11109 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_246
timestamp 1606744421
transform 1 0 10273 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_247
timestamp 1606744421
transform 1 0 9437 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_248
timestamp 1606744421
transform 1 0 8601 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_249
timestamp 1606744421
transform 1 0 7765 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_250
timestamp 1606744421
transform 1 0 6929 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_251
timestamp 1606744421
transform 1 0 6093 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_252
timestamp 1606744421
transform 1 0 5257 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_253
timestamp 1606744421
transform 1 0 4421 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_254
timestamp 1606744421
transform 1 0 9505 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_255
timestamp 1606744421
transform 1 0 8669 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_256
timestamp 1606744421
transform 1 0 7833 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_257
timestamp 1606744421
transform 1 0 6997 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_258
timestamp 1606744421
transform 1 0 6161 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_259
timestamp 1606744421
transform 1 0 5325 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_260
timestamp 1606744421
transform 1 0 4489 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_261
timestamp 1606744421
transform 1 0 9437 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_262
timestamp 1606744421
transform 1 0 8601 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_263
timestamp 1606744421
transform 1 0 7765 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_264
timestamp 1606744421
transform 1 0 6929 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_265
timestamp 1606744421
transform 1 0 6093 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_266
timestamp 1606744421
transform 1 0 5257 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_267
timestamp 1606744421
transform 1 0 4421 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_268
timestamp 1606744421
transform 1 0 3653 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_269
timestamp 1606744421
transform 1 0 3585 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_270
timestamp 1606744421
transform 1 0 3653 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_271
timestamp 1606744421
transform 1 0 3585 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_272
timestamp 1606744421
transform 1 0 12849 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_273
timestamp 1606744421
transform 1 0 12013 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_274
timestamp 1606744421
transform 1 0 11177 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_275
timestamp 1606744421
transform 1 0 10341 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_276
timestamp 1606744421
transform 1 0 12781 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_277
timestamp 1606744421
transform 1 0 11945 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_278
timestamp 1606744421
transform 1 0 11109 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_279
timestamp 1606744421
transform 1 0 10273 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_280
timestamp 1606744421
transform 1 0 12849 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_281
timestamp 1606744421
transform 1 0 12013 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_282
timestamp 1606744421
transform 1 0 11177 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_283
timestamp 1606744421
transform 1 0 10341 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_284
timestamp 1606744421
transform 1 0 4489 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_285
timestamp 1606744421
transform 1 0 9437 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_286
timestamp 1606744421
transform 1 0 11945 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_287
timestamp 1606744421
transform 1 0 11109 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_288
timestamp 1606744421
transform 1 0 10273 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_289
timestamp 1606744421
transform 1 0 9505 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_290
timestamp 1606744421
transform 1 0 8669 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_291
timestamp 1606744421
transform 1 0 7833 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_292
timestamp 1606744421
transform 1 0 6997 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_293
timestamp 1606744421
transform 1 0 6161 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_294
timestamp 1606744421
transform 1 0 11814 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_295
timestamp 1606744421
transform 1 0 12368 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_296
timestamp 1606744421
transform 1 0 5788 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_297
timestamp 1606744421
transform 1 0 6342 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_298
timestamp 1606744421
transform 1 0 6896 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_299
timestamp 1606744421
transform 1 0 11328 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_300
timestamp 1606744421
transform 1 0 6828 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_301
timestamp 1606744421
transform 1 0 5325 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_302
timestamp 1606744421
transform 1 0 12781 0 1 31372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_303
timestamp 1606744421
transform 1 0 8601 0 1 29372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_304
timestamp 1606744421
transform 1 0 3653 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_305
timestamp 1606744421
transform 1 0 3585 0 1 33372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_306
timestamp 1606744421
transform 1 0 6896 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_307
timestamp 1606744421
transform 1 0 7450 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_308
timestamp 1606744421
transform 1 0 8004 0 -1 12722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_309
timestamp 1606744421
transform 1 0 6997 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_310
timestamp 1606744421
transform 1 0 6929 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_311
timestamp 1606744421
transform 1 0 6161 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_312
timestamp 1606744421
transform 1 0 6093 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_313
timestamp 1606744421
transform 1 0 5325 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_314
timestamp 1606744421
transform 1 0 5257 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_315
timestamp 1606744421
transform 1 0 7765 0 1 27372
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_316
timestamp 1606744421
transform 1 0 11882 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808682  sky130_fd_pr__dfl1__example_55959141808682_317
timestamp 1606744421
transform 1 0 12436 0 -1 36722
box 0 -4 50 1354
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_0
timestamp 1606744421
transform 1 0 12922 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_1
timestamp 1606744421
transform 1 0 12990 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_2
timestamp 1606744421
transform 1 0 2950 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_3
timestamp 1606744421
transform 1 0 3018 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_4
timestamp 1606744421
transform 1 0 3504 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_5
timestamp 1606744421
transform 1 0 3572 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_6
timestamp 1606744421
transform 1 0 4058 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_7
timestamp 1606744421
transform 1 0 4126 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_8
timestamp 1606744421
transform 1 0 4612 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_9
timestamp 1606744421
transform 1 0 4680 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_10
timestamp 1606744421
transform 1 0 5166 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_11
timestamp 1606744421
transform 1 0 5234 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_12
timestamp 1606744421
transform 1 0 5720 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_13
timestamp 1606744421
transform 1 0 6274 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_14
timestamp 1606744421
transform 1 0 6828 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_15
timestamp 1606744421
transform 1 0 7382 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_16
timestamp 1606744421
transform 1 0 7936 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_17
timestamp 1606744421
transform 1 0 8490 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_18
timestamp 1606744421
transform 1 0 9044 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_19
timestamp 1606744421
transform 1 0 9598 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_20
timestamp 1606744421
transform 1 0 10152 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_21
timestamp 1606744421
transform 1 0 10706 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_22
timestamp 1606744421
transform 1 0 5788 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_23
timestamp 1606744421
transform 1 0 6342 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_24
timestamp 1606744421
transform 1 0 6896 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_25
timestamp 1606744421
transform 1 0 7450 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_26
timestamp 1606744421
transform 1 0 8004 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_27
timestamp 1606744421
transform 1 0 8558 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_28
timestamp 1606744421
transform 1 0 9112 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_29
timestamp 1606744421
transform 1 0 9666 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_30
timestamp 1606744421
transform 1 0 10220 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_31
timestamp 1606744421
transform 1 0 10774 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_32
timestamp 1606744421
transform 1 0 11260 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_33
timestamp 1606744421
transform 1 0 11814 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_34
timestamp 1606744421
transform 1 0 12368 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_35
timestamp 1606744421
transform 1 0 11328 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_36
timestamp 1606744421
transform 1 0 11882 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_37
timestamp 1606744421
transform 1 0 12436 0 -1 14341
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_38
timestamp 1606744421
transform 1 0 12849 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_39
timestamp 1606744421
transform 1 0 12013 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_40
timestamp 1606744421
transform 1 0 11177 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_41
timestamp 1606744421
transform 1 0 10341 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_42
timestamp 1606744421
transform 1 0 9505 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_43
timestamp 1606744421
transform 1 0 8669 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_44
timestamp 1606744421
transform 1 0 7833 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_45
timestamp 1606744421
transform 1 0 12781 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_46
timestamp 1606744421
transform 1 0 11945 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_47
timestamp 1606744421
transform 1 0 11109 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_48
timestamp 1606744421
transform 1 0 10273 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_49
timestamp 1606744421
transform 1 0 9437 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_50
timestamp 1606744421
transform 1 0 8601 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_51
timestamp 1606744421
transform 1 0 6997 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_52
timestamp 1606744421
transform 1 0 6929 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_53
timestamp 1606744421
transform 1 0 6161 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_54
timestamp 1606744421
transform 1 0 6093 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_55
timestamp 1606744421
transform 1 0 5325 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_56
timestamp 1606744421
transform 1 0 5257 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__dfl1__example_55959141808681  sky130_fd_pr__dfl1__example_55959141808681_57
timestamp 1606744421
transform 1 0 7765 0 1 25780
box 0 -4 50 946
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1606744421
transform 0 -1 114 1 0 3722
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1606744421
transform 0 -1 1734 1 0 39154
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808705  sky130_fd_pr__nfet_01v8__example_55959141808705_0
timestamp 1606744421
transform 1 0 2872 0 1 5372
box -240 -32 10486 1432
use sky130_fd_pr__nfet_01v8__example_55959141808705  sky130_fd_pr__nfet_01v8__example_55959141808705_1
timestamp 1606744421
transform 1 0 2872 0 1 9372
box -240 -32 10486 1432
use sky130_fd_pr__nfet_01v8__example_55959141808705  sky130_fd_pr__nfet_01v8__example_55959141808705_2
timestamp 1606744421
transform 1 0 2872 0 1 11372
box -240 -32 10486 1432
use sky130_fd_pr__nfet_01v8__example_55959141808705  sky130_fd_pr__nfet_01v8__example_55959141808705_3
timestamp 1606744421
transform 1 0 2872 0 1 37372
box -240 -32 10486 1432
use sky130_fd_pr__nfet_01v8__example_55959141808705  sky130_fd_pr__nfet_01v8__example_55959141808705_4
timestamp 1606744421
transform 1 0 2872 0 1 7372
box -240 -32 10486 1432
use sky130_fd_pr__nfet_01v8__example_55959141808704  sky130_fd_pr__nfet_01v8__example_55959141808704_0
timestamp 1606744421
transform 1 0 5163 0 1 27372
box -365 -32 8195 1432
use sky130_fd_pr__nfet_01v8__example_55959141808703  sky130_fd_pr__nfet_01v8__example_55959141808703_0
timestamp 1606744421
transform 1 0 3491 0 1 29372
box -365 -32 9867 1432
use sky130_fd_pr__nfet_01v8__example_55959141808703  sky130_fd_pr__nfet_01v8__example_55959141808703_1
timestamp 1606744421
transform 1 0 3491 0 1 31372
box -365 -32 9867 1432
use sky130_fd_pr__nfet_01v8__example_55959141808703  sky130_fd_pr__nfet_01v8__example_55959141808703_2
timestamp 1606744421
transform 1 0 3491 0 1 33372
box -365 -32 9867 1432
use sky130_fd_pr__nfet_01v8__example_55959141808701  sky130_fd_pr__nfet_01v8__example_55959141808701_0
timestamp 1606744421
transform 1 0 3426 0 1 35372
box -240 -32 9932 1432
use sky130_fd_pr__nfet_01v8__example_55959141808699  sky130_fd_pr__nfet_01v8__example_55959141808699_0
timestamp 1606744421
transform 1 0 5107 0 1 21980
box -53 -32 8277 1432
use sky130_fd_pr__nfet_01v8__example_55959141808699  sky130_fd_pr__nfet_01v8__example_55959141808699_1
timestamp 1606744421
transform 1 0 5107 0 1 18260
box -53 -32 8277 1432
use sky130_fd_pr__nfet_01v8__example_55959141808699  sky130_fd_pr__nfet_01v8__example_55959141808699_2
timestamp 1606744421
transform 1 0 5107 0 -1 25145
box -53 -32 8277 1432
use sky130_fd_pr__nfet_01v8__example_55959141808699  sky130_fd_pr__nfet_01v8__example_55959141808699_3
timestamp 1606744421
transform 1 0 5107 0 1 20281
box -53 -32 8277 1432
use sky130_fd_pr__nfet_01v8__example_55959141808699  sky130_fd_pr__nfet_01v8__example_55959141808699_4
timestamp 1606744421
transform 1 0 5107 0 1 16561
box -53 -32 8277 1432
use sky130_fd_pr__nfet_01v8__example_55959141808698  sky130_fd_pr__nfet_01v8__example_55959141808698_0
timestamp 1606744421
transform 1 0 3451 0 1 15161
box -53 -32 9933 1032
use sky130_fd_pr__nfet_01v8__example_55959141808697  sky130_fd_pr__nfet_01v8__example_55959141808697_0
timestamp 1606744421
transform -1 0 3395 0 1 15161
box -53 -32 853 1032
use sky130_fd_pr__nfet_01v8__example_55959141808696  sky130_fd_pr__nfet_01v8__example_55959141808696_0
timestamp 1606744421
transform 1 0 4934 0 -1 25145
box -136 -32 173 1432
use sky130_fd_pr__nfet_01v8__example_55959141808696  sky130_fd_pr__nfet_01v8__example_55959141808696_1
timestamp 1606744421
transform 1 0 4934 0 1 21980
box -136 -32 173 1432
use sky130_fd_pr__nfet_01v8__example_55959141808696  sky130_fd_pr__nfet_01v8__example_55959141808696_2
timestamp 1606744421
transform 1 0 4934 0 1 16561
box -136 -32 173 1432
use sky130_fd_pr__nfet_01v8__example_55959141808696  sky130_fd_pr__nfet_01v8__example_55959141808696_3
timestamp 1606744421
transform 1 0 4934 0 1 20281
box -136 -32 173 1432
use sky130_fd_pr__nfet_01v8__example_55959141808696  sky130_fd_pr__nfet_01v8__example_55959141808696_4
timestamp 1606744421
transform 1 0 4934 0 1 18260
box -136 -32 173 1432
use sky130_fd_pr__nfet_01v8__example_55959141808695  sky130_fd_pr__nfet_01v8__example_55959141808695_0
timestamp 1606744421
transform 1 0 5163 0 1 25751
box -365 -32 8195 1032
use sky130_fd_pr__nfet_01v8__example_55959141808693  sky130_fd_pr__nfet_01v8__example_55959141808693_0
timestamp 1606744421
transform 1 0 2872 0 1 13372
box -240 -32 10486 1032
use sky130_fd_pr__res_bent_po__example_55959141808692  sky130_fd_pr__res_bent_po__example_55959141808692_0
timestamp 1606744421
transform 0 -1 14193 1 0 3626
box -50 -648 35946 66
use sky130_fd_pr__res_bent_po__example_55959141808691  sky130_fd_pr__res_bent_po__example_55959141808691_0
timestamp 1606744421
transform 0 1 13357 1 0 349
box -50 -1944 3007 66
use sky130_fd_pr__res_bent_po__example_55959141808690  sky130_fd_pr__res_bent_po__example_55959141808690_0
timestamp 1606744421
transform -1 0 13955 0 -1 3902
box -50 -648 11946 66
use sky130_fd_pr__res_bent_po__example_55959141808689  sky130_fd_pr__res_bent_po__example_55959141808689_0
timestamp 1606744421
transform 0 -1 114 1 0 3840
box -50 -1620 35387 66
use sky130_fd_pr__res_bent_po__example_55959141808688  sky130_fd_pr__res_bent_po__example_55959141808688_0
timestamp 1606744421
transform 0 -1 2249 1 0 16866
box -50 -1782 11931 66
use sky130_fd_pr__pfet_01v8__example_55959141808687  sky130_fd_pr__pfet_01v8__example_55959141808687_0
timestamp 1606744421
transform 1 0 13667 0 1 416
box -92 -36 956 1436
use sky130_fd_pr__pfet_01v8__example_55959141808687  sky130_fd_pr__pfet_01v8__example_55959141808687_1
timestamp 1606744421
transform 1 0 13667 0 1 1946
box -92 -36 956 1436
use sky130_fd_pr__pfet_01v8__example_55959141808687  sky130_fd_pr__pfet_01v8__example_55959141808687_2
timestamp 1606744421
transform 1 0 414 0 1 1934
box -92 -36 956 1436
use sky130_fd_pr__pfet_01v8__example_55959141808687  sky130_fd_pr__pfet_01v8__example_55959141808687_3
timestamp 1606744421
transform 1 0 414 0 1 404
box -92 -36 956 1436
use sky130_fd_io__gnd2gnd_120x2_lv_isosub  sky130_fd_io__gnd2gnd_120x2_lv_isosub_0
timestamp 1606744421
transform 1 0 3305 0 -1 3696
box 26 26 8008 3632
use sky130_fd_io__com_busses_esd  sky130_fd_io__com_busses_esd_0
timestamp 1606744421
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal4 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal4 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal4 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 4 nsew power bidirectional
flabel metal4 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 5 nsew power bidirectional
flabel metal4 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 4 nsew power bidirectional
flabel metal4 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 5 nsew power bidirectional
flabel metal4 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal4 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal4 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 9 nsew power bidirectional
flabel metal4 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 10 nsew signal bidirectional
flabel metal4 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 9 nsew power bidirectional
flabel metal4 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 10 nsew signal bidirectional
flabel metal4 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 12 nsew ground bidirectional
flabel metal4 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 12 nsew ground bidirectional
flabel metal4 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal4 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal5 6339 32553 10468 33424 0 FreeSans 2000 0 0 0 G_PAD
port 13 nsew signal bidirectional
flabel metal5 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal5 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal5 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal5 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal5 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal5 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 12 nsew ground bidirectional
flabel metal5 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 9 nsew power bidirectional
flabel metal5 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 5 nsew power bidirectional
flabel metal5 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 7 nsew ground bidirectional
flabel metal5 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 12 nsew ground bidirectional
flabel metal5 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 9 nsew power bidirectional
flabel metal5 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 5 nsew power bidirectional
flabel metal5 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel comment s 8128 39216 8128 39216 0 FreeSans 600 0 0 0 CONDIODE
flabel comment s 8037 22958 8037 22958 0 FreeSans 600 0 0 0 CONDIODE
flabel comment s 8121 6986 8121 6986 0 FreeSans 600 0 0 0 CONDIODE
flabel metal2 100 0 4099 294 0 FreeSans 2000 0 0 0 SRC_BDY_LVC1
port 14 nsew ground bidirectional
flabel metal2 10953 0 14940 722 0 FreeSans 2000 0 0 0 SRC_BDY_LVC2
port 15 nsew ground bidirectional
flabel metal2 6888 0 8888 65 0 FreeSans 400 0 0 0 BDY2_B2B
port 16 nsew ground bidirectional
flabel metal3 7676 0 9850 925 0 FreeSans 2000 0 0 0 DRN_LVC2
port 17 nsew power bidirectional
flabel metal3 5200 0 7374 925 0 FreeSans 2000 0 0 0 DRN_LVC1
port 18 nsew power bidirectional
flabel metal1 5242 0 5540 28 0 FreeSans 200 0 0 0 OGC_LVC
port 20 nsew power bidirectional
rlabel metal3 s 12409 19151 14940 34447 1 G_CORE
port 19 nsew ground bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string GDS_FILE /home/roshan/Desktop/pdks/sky130A/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 35304112
string GDS_START 31685712
<< end >>
