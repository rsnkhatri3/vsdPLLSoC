# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# High density, double height
SITE unithddbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 0.34 ;
  OFFSET 0.23 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.2 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.34 ;
  OFFSET 0.17 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 ;
  OFFSET 0.23 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;

  EDGECAPACITANCE 37.759E-6 ;
  CAPACITANCE CPERSQDIST 16.9423E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.68 ;
  OFFSET 0.34 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 40.989E-6 ;
  CAPACITANCE CPERSQDIST 12.3729E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.92 ;
  OFFSET 0.46 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;            # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 36.676E-6 ;
  CAPACITANCE CPERSQDIST 8.41537E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.4 ;
  OFFSET 1.7 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 38.851E-6 ;
  CAPACITANCE CPERSQDIST 6.32063E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###



MACRO sky130_fd_sc_hd__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 1.075 1.39 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.67 1.445 ;
        RECT 0.425 1.445 1.73 1.615 ;
        RECT 1.56 1.075 1.935 1.245 ;
        RECT 1.56 1.245 1.73 1.445 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.800500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.72 0.315 2.675 0.485 ;
        RECT 2.505 0.485 2.675 1.365 ;
        RECT 2.505 1.365 3.135 1.535 ;
        RECT 2.815 1.535 3.135 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.655 2.335 0.825 ;
      RECT 0.085 0.825 0.255 1.785 ;
      RECT 0.085 1.785 0.465 2.465 ;
      RECT 0.135 0.085 0.465 0.475 ;
      RECT 0.635 0.335 0.805 0.655 ;
      RECT 0.975 0.085 1.305 0.475 ;
      RECT 1.055 1.785 1.225 2.635 ;
      RECT 1.395 1.785 2.635 1.955 ;
      RECT 1.395 1.955 1.725 2.465 ;
      RECT 1.895 2.125 2.065 2.635 ;
      RECT 2.105 0.825 2.335 1.325 ;
      RECT 2.235 1.955 2.635 2.465 ;
      RECT 2.845 0.085 3.135 0.92 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__xor2_1
MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 0.875 1.275 ;
        RECT 0.705 1.275 0.875 1.445 ;
        RECT 0.705 1.445 1.88 1.615 ;
        RECT 1.71 1.075 3.23 1.275 ;
        RECT 1.71 1.275 1.88 1.445 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.54 1.275 ;
      LAYER mcon ;
        RECT 1.065 1.105 1.235 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.42 1.075 4.09 1.275 ;
      LAYER mcon ;
        RECT 3.825 1.105 3.995 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.005 1.075 1.295 1.12 ;
        RECT 1.005 1.12 4.055 1.26 ;
        RECT 1.005 1.26 1.295 1.305 ;
        RECT 3.765 1.075 4.055 1.12 ;
        RECT 3.765 1.26 4.055 1.305 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.656750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.625 0.645 3.955 0.725 ;
        RECT 3.625 0.725 5.895 0.905 ;
        RECT 4.985 0.645 5.315 0.725 ;
        RECT 5.025 1.415 5.895 1.625 ;
        RECT 5.025 1.625 5.275 2.125 ;
        RECT 5.485 0.905 5.895 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.12 0.725 1.7 0.905 ;
      RECT 0.12 0.905 0.29 1.785 ;
      RECT 0.12 1.785 2.22 1.955 ;
      RECT 0.12 2.135 0.4 2.465 ;
      RECT 0.145 2.125 0.315 2.135 ;
      RECT 0.19 0.085 0.36 0.555 ;
      RECT 0.53 0.255 0.86 0.725 ;
      RECT 0.57 2.135 0.82 2.635 ;
      RECT 0.99 2.135 1.24 2.295 ;
      RECT 0.99 2.295 2.08 2.465 ;
      RECT 1.03 0.085 1.2 0.555 ;
      RECT 1.065 2.125 1.235 2.135 ;
      RECT 1.37 0.255 1.7 0.725 ;
      RECT 1.41 1.955 1.66 2.125 ;
      RECT 1.83 2.135 2.08 2.295 ;
      RECT 1.87 0.085 2.04 0.555 ;
      RECT 2.05 1.445 4.785 1.615 ;
      RECT 2.05 1.615 2.22 1.785 ;
      RECT 2.285 2.125 2.6 2.465 ;
      RECT 2.31 0.255 2.64 0.725 ;
      RECT 2.31 0.725 3.4 0.905 ;
      RECT 2.39 1.785 4.855 1.955 ;
      RECT 2.39 1.955 2.6 2.125 ;
      RECT 2.77 2.135 3.02 2.635 ;
      RECT 2.81 0.085 2.98 0.555 ;
      RECT 3.15 0.255 4.38 0.475 ;
      RECT 3.15 0.475 3.4 0.725 ;
      RECT 3.19 1.955 3.44 2.465 ;
      RECT 3.61 2.135 3.915 2.635 ;
      RECT 4.085 1.955 4.855 2.295 ;
      RECT 4.085 2.295 5.695 2.465 ;
      RECT 4.615 1.075 5.275 1.245 ;
      RECT 4.615 1.245 4.785 1.445 ;
      RECT 4.645 0.085 4.815 0.555 ;
      RECT 5.445 1.795 5.695 2.295 ;
      RECT 5.485 0.085 5.655 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 0.085 2.095 0.375 2.14 ;
      RECT 0.085 2.14 1.295 2.28 ;
      RECT 0.085 2.28 0.375 2.325 ;
      RECT 1.005 2.095 1.295 2.14 ;
      RECT 1.005 2.28 1.295 2.325 ;
  END
END sky130_fd_sc_hd__xor2_2
MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 2.8 1.275 ;
        RECT 2.63 1.275 2.8 1.445 ;
        RECT 2.63 1.445 6.165 1.615 ;
        RECT 5.995 1.075 7.37 1.275 ;
        RECT 5.995 1.275 6.165 1.445 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.075 5 1.105 ;
        RECT 2.97 1.105 5.74 1.275 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.524450 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 0.645 5.58 0.905 ;
        RECT 5.15 0.905 5.58 0.935 ;
      LAYER mcon ;
        RECT 5.205 0.765 5.375 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.85 0.725 8.63 0.735 ;
        RECT 7.85 0.735 10.035 0.905 ;
        RECT 7.85 0.905 8.305 0.935 ;
        RECT 7.88 1.445 10.035 1.625 ;
        RECT 7.88 1.625 9.01 1.665 ;
        RECT 7.88 1.665 8.17 2.125 ;
        RECT 8.3 0.255 8.63 0.725 ;
        RECT 8.76 1.665 9.01 2.125 ;
        RECT 9.14 0.255 9.47 0.735 ;
        RECT 9.6 1.625 10.035 2.465 ;
        RECT 9.735 0.905 10.035 1.445 ;
      LAYER mcon ;
        RECT 7.965 0.765 8.135 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.145 0.735 5.435 0.78 ;
        RECT 5.145 0.78 8.195 0.92 ;
        RECT 5.145 0.92 5.435 0.965 ;
        RECT 7.905 0.735 8.195 0.78 ;
        RECT 7.905 0.92 8.195 0.965 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.085 0.085 0.36 0.565 ;
      RECT 0.085 0.735 3.38 0.905 ;
      RECT 0.085 0.905 0.255 1.445 ;
      RECT 0.085 1.445 2.42 1.615 ;
      RECT 0.085 1.785 2.08 2.005 ;
      RECT 0.085 2.005 0.4 2.465 ;
      RECT 0.53 0.255 0.86 0.725 ;
      RECT 0.53 0.725 3.38 0.735 ;
      RECT 0.57 2.175 0.82 2.635 ;
      RECT 0.99 2.005 1.24 2.465 ;
      RECT 1.03 0.085 1.2 0.555 ;
      RECT 1.37 0.255 1.7 0.725 ;
      RECT 1.41 2.175 1.66 2.635 ;
      RECT 1.83 2.005 2.08 2.295 ;
      RECT 1.83 2.295 3.76 2.465 ;
      RECT 1.87 0.085 2.04 0.555 ;
      RECT 2.21 0.255 2.54 0.725 ;
      RECT 2.25 1.615 2.42 1.785 ;
      RECT 2.25 1.785 3.34 1.955 ;
      RECT 2.25 1.955 2.5 2.125 ;
      RECT 2.67 2.125 2.92 2.295 ;
      RECT 2.71 0.085 2.88 0.555 ;
      RECT 3.05 0.255 3.38 0.725 ;
      RECT 3.09 1.955 3.34 2.125 ;
      RECT 3.51 1.795 3.76 2.295 ;
      RECT 3.55 0.085 3.82 0.895 ;
      RECT 3.99 0.255 6 0.475 ;
      RECT 4.03 1.785 7.64 2.005 ;
      RECT 4.03 2.005 4.28 2.465 ;
      RECT 4.45 2.175 4.7 2.635 ;
      RECT 4.87 2.005 5.12 2.465 ;
      RECT 5.29 2.175 5.54 2.635 ;
      RECT 5.71 2.005 5.96 2.465 ;
      RECT 5.75 0.475 6 0.725 ;
      RECT 5.75 0.725 7.68 0.905 ;
      RECT 6.13 2.175 6.38 2.635 ;
      RECT 6.17 0.085 6.34 0.555 ;
      RECT 6.51 0.255 6.84 0.725 ;
      RECT 6.55 1.455 6.8 1.785 ;
      RECT 6.55 2.005 6.8 2.465 ;
      RECT 6.97 2.175 7.22 2.635 ;
      RECT 7.01 0.085 7.18 0.555 ;
      RECT 7.26 1.445 7.71 1.615 ;
      RECT 7.35 0.255 7.68 0.725 ;
      RECT 7.39 2.005 7.64 2.295 ;
      RECT 7.39 2.295 9.43 2.465 ;
      RECT 7.54 1.105 9.565 1.275 ;
      RECT 7.54 1.275 7.71 1.445 ;
      RECT 7.96 0.085 8.13 0.555 ;
      RECT 8.34 1.835 8.59 2.295 ;
      RECT 8.54 1.075 9.565 1.105 ;
      RECT 8.8 0.085 8.97 0.555 ;
      RECT 9.18 1.795 9.43 2.295 ;
      RECT 9.64 0.085 9.81 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 1.445 2.155 1.615 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 1.445 7.675 1.615 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
    LAYER met1 ;
      RECT 1.925 1.415 2.215 1.46 ;
      RECT 1.925 1.46 7.735 1.6 ;
      RECT 1.925 1.6 2.215 1.645 ;
      RECT 7.445 1.415 7.735 1.46 ;
      RECT 7.445 1.6 7.735 1.645 ;
  END
END sky130_fd_sc_hd__xor2_4
MACRO sky130_fd_sc_hd__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.28 1.68 0.735 ;
        RECT 1.42 0.735 4.73 0.905 ;
        RECT 1.42 1.495 4.73 1.735 ;
        RECT 1.42 1.735 1.68 2.46 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 3.76 0.905 4.73 1.495 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.095 1.525 0.39 2.635 ;
      RECT 0.145 0.085 0.39 0.545 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 3.59 1.325 ;
      RECT 0.57 1.325 0.82 2.46 ;
      RECT 0.99 0.085 1.25 0.61 ;
      RECT 0.99 1.525 1.25 2.635 ;
      RECT 1.85 0.085 2.11 0.565 ;
      RECT 1.85 1.905 2.11 2.635 ;
      RECT 2.71 0.085 2.97 0.565 ;
      RECT 2.71 1.905 2.97 2.635 ;
      RECT 3.57 0.085 3.83 0.565 ;
      RECT 3.57 1.905 3.83 2.635 ;
      RECT 4.43 0.085 4.73 0.565 ;
      RECT 4.43 1.905 4.725 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__clkbuf_8
MACRO sky130_fd_sc_hd__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 0.735 9.025 0.905 ;
        RECT 2.28 1.495 9.025 1.72 ;
        RECT 2.28 1.72 7.685 1.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
        RECT 4.845 0.28 5.12 0.735 ;
        RECT 4.86 1.735 5.12 2.46 ;
        RECT 5.705 0.28 5.965 0.735 ;
        RECT 5.705 1.735 5.965 2.46 ;
        RECT 6.565 0.28 6.825 0.735 ;
        RECT 6.565 1.735 6.825 2.46 ;
        RECT 7.425 0.28 7.685 0.735 ;
        RECT 7.425 1.735 7.685 2.46 ;
        RECT 7.86 0.905 9.025 1.495 ;
        RECT 8.295 0.28 8.555 0.735 ;
        RECT 8.295 1.72 8.585 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.085 0.085 0.39 0.595 ;
      RECT 0.095 1.825 0.39 2.635 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 7.69 1.325 ;
      RECT 0.57 1.325 0.815 2.465 ;
      RECT 0.99 0.085 1.25 0.61 ;
      RECT 0.99 1.825 1.25 2.635 ;
      RECT 1.43 0.265 1.68 1.075 ;
      RECT 1.43 1.325 1.68 2.46 ;
      RECT 1.85 0.085 2.11 0.645 ;
      RECT 1.85 1.835 2.11 2.63 ;
      RECT 1.85 2.63 8.125 2.635 ;
      RECT 2.71 0.085 2.97 0.565 ;
      RECT 2.71 1.905 2.97 2.63 ;
      RECT 3.57 0.085 3.83 0.565 ;
      RECT 3.57 1.905 3.83 2.63 ;
      RECT 4.43 0.085 4.675 0.565 ;
      RECT 4.43 1.905 4.69 2.63 ;
      RECT 5.29 0.085 5.535 0.565 ;
      RECT 5.29 1.905 5.535 2.63 ;
      RECT 6.145 0.085 6.395 0.565 ;
      RECT 6.15 1.905 6.395 2.63 ;
      RECT 7.005 0.085 7.255 0.565 ;
      RECT 7.01 1.905 7.255 2.63 ;
      RECT 7.865 0.085 8.125 0.565 ;
      RECT 7.87 1.905 8.125 2.63 ;
      RECT 8.725 0.085 9.025 0.565 ;
      RECT 8.755 1.89 9.025 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
  END
END sky130_fd_sc_hd__clkbuf_16
MACRO sky130_fd_sc_hd__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.345 1.305 0.735 ;
        RECT 1.01 0.735 2.66 0.905 ;
        RECT 1.045 1.835 2.165 2.005 ;
        RECT 1.045 2.005 1.305 2.465 ;
        RECT 1.905 0.345 2.165 0.735 ;
        RECT 1.905 1.415 2.66 1.585 ;
        RECT 1.905 1.585 2.165 1.835 ;
        RECT 1.905 2.005 2.165 2.465 ;
        RECT 2.255 0.905 2.66 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.255 0.385 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.115 1.665 ;
      RECT 0.085 1.665 0.395 2.465 ;
      RECT 0.555 0.085 0.83 0.565 ;
      RECT 0.565 1.835 0.875 2.635 ;
      RECT 0.945 1.075 2.085 1.245 ;
      RECT 0.945 1.245 1.115 1.495 ;
      RECT 1.475 0.085 1.73 0.565 ;
      RECT 1.475 2.175 1.73 2.635 ;
      RECT 2.335 0.085 2.615 0.565 ;
      RECT 2.335 1.765 2.62 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__clkbuf_4
MACRO sky130_fd_sc_hd__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.255 1.245 0.655 ;
        RECT 1.04 0.655 1.725 0.825 ;
        RECT 1.06 1.855 1.725 2.03 ;
        RECT 1.06 2.03 1.245 2.435 ;
        RECT 1.385 0.825 1.725 1.855 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.215 1.665 ;
      RECT 0.085 1.665 0.355 2.435 ;
      RECT 0.525 1.855 0.855 2.635 ;
      RECT 0.555 0.085 0.83 0.565 ;
      RECT 0.965 0.995 1.215 1.495 ;
      RECT 1.415 0.085 1.75 0.485 ;
      RECT 1.415 2.21 1.75 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__clkbuf_2
MACRO sky130_fd_sc_hd__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.76 ;
        RECT 0.085 0.76 0.255 1.56 ;
        RECT 0.085 1.56 0.355 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065 -0.085 1.235 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.425 1.06 0.71 1.39 ;
      RECT 0.525 0.085 0.855 0.465 ;
      RECT 0.525 1.875 0.855 2.635 ;
      RECT 0.54 0.635 1.205 0.805 ;
      RECT 0.54 0.805 0.71 1.06 ;
      RECT 0.54 1.39 0.71 1.535 ;
      RECT 0.54 1.535 1.205 1.705 ;
      RECT 1.035 0.255 1.205 0.635 ;
      RECT 1.035 1.705 1.205 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__clkbuf_1
MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 1.005 2.17 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.115 0.255 12.345 0.825 ;
        RECT 12.115 1.445 12.345 2.465 ;
        RECT 12.16 0.825 12.345 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.24 0.255 10.5 0.715 ;
        RECT 10.24 1.63 10.5 2.465 ;
        RECT 10.32 0.715 10.5 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.25 1.095 9.73 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.6 0.735 4.01 0.965 ;
        RECT 3.6 0.965 3.93 1.065 ;
      LAYER mcon ;
        RECT 3.84 0.765 4.01 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.47 0.735 7.845 1.065 ;
      LAYER mcon ;
        RECT 7.52 0.765 7.69 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.78 0.735 4.07 0.78 ;
        RECT 3.78 0.78 7.75 0.92 ;
        RECT 3.78 0.92 4.07 0.965 ;
        RECT 7.46 0.735 7.75 0.78 ;
        RECT 7.46 0.92 7.75 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.44 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 13.07 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.88 0.085 ;
      RECT 0 2.635 12.88 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.84 0.805 ;
      RECT 0.085 1.795 0.84 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.42 0.635 2.125 0.825 ;
      RECT 1.42 0.825 1.59 1.795 ;
      RECT 1.42 1.795 2.125 1.965 ;
      RECT 1.445 0.085 1.785 0.465 ;
      RECT 1.445 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.34 0.705 2.56 1.575 ;
      RECT 2.34 1.575 2.84 1.955 ;
      RECT 2.35 2.25 3.18 2.42 ;
      RECT 2.415 0.265 3.41 0.465 ;
      RECT 2.74 0.645 3.07 1.015 ;
      RECT 3.01 1.195 3.41 1.235 ;
      RECT 3.01 1.235 4.36 1.405 ;
      RECT 3.01 1.405 3.18 2.25 ;
      RECT 3.24 0.465 3.41 1.195 ;
      RECT 3.35 1.575 3.6 1.785 ;
      RECT 3.35 1.785 4.7 2.035 ;
      RECT 3.42 2.205 3.8 2.635 ;
      RECT 3.58 0.085 3.75 0.525 ;
      RECT 3.92 0.255 5.17 0.425 ;
      RECT 3.92 0.425 4.25 0.545 ;
      RECT 4.1 2.035 4.27 2.375 ;
      RECT 4.11 1.405 4.36 1.485 ;
      RECT 4.14 1.155 4.36 1.235 ;
      RECT 4.42 0.595 4.75 0.765 ;
      RECT 4.53 0.765 4.75 0.895 ;
      RECT 4.53 0.895 5.84 1.065 ;
      RECT 4.53 1.065 4.7 1.785 ;
      RECT 4.87 1.235 5.2 1.415 ;
      RECT 4.87 1.415 5.875 1.655 ;
      RECT 4.89 1.915 5.22 2.635 ;
      RECT 4.92 0.425 5.17 0.715 ;
      RECT 5.36 0.085 5.69 0.465 ;
      RECT 5.51 1.065 5.84 1.235 ;
      RECT 6.075 1.575 6.31 1.985 ;
      RECT 6.135 0.705 6.42 1.125 ;
      RECT 6.135 1.125 6.755 1.305 ;
      RECT 6.265 2.25 7.095 2.42 ;
      RECT 6.33 0.265 7.095 0.465 ;
      RECT 6.55 1.305 6.755 1.905 ;
      RECT 6.925 0.465 7.095 1.235 ;
      RECT 6.925 1.235 8.275 1.405 ;
      RECT 6.925 1.405 7.095 2.25 ;
      RECT 7.265 1.575 7.515 1.915 ;
      RECT 7.265 1.915 10.07 2.085 ;
      RECT 7.275 0.085 7.535 0.525 ;
      RECT 7.335 2.255 7.715 2.635 ;
      RECT 7.795 0.255 8.965 0.425 ;
      RECT 7.795 0.425 8.125 0.545 ;
      RECT 7.955 2.085 8.125 2.375 ;
      RECT 8.055 1.075 8.275 1.235 ;
      RECT 8.295 0.595 8.625 0.78 ;
      RECT 8.445 0.78 8.625 1.915 ;
      RECT 8.655 2.255 10.07 2.635 ;
      RECT 8.795 0.425 8.965 0.585 ;
      RECT 8.795 0.755 9.5 0.925 ;
      RECT 8.795 0.925 9.07 1.575 ;
      RECT 8.795 1.575 9.57 1.745 ;
      RECT 9.28 0.265 9.5 0.755 ;
      RECT 9.74 0.085 10.07 0.805 ;
      RECT 9.9 0.995 10.14 1.325 ;
      RECT 9.9 1.325 10.07 1.915 ;
      RECT 10.68 0.085 10.91 0.885 ;
      RECT 10.68 1.465 10.91 2.635 ;
      RECT 11.215 0.255 11.47 0.995 ;
      RECT 11.215 0.995 11.99 1.325 ;
      RECT 11.215 1.325 11.47 2.415 ;
      RECT 11.65 0.085 11.945 0.545 ;
      RECT 11.65 1.765 11.945 2.635 ;
      RECT 12.515 0.085 12.795 0.885 ;
      RECT 12.515 1.465 12.795 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 0.765 0.78 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.46 1.785 2.63 1.955 ;
      RECT 2.9 0.765 3.07 0.935 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.68 1.445 5.85 1.615 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.14 1.105 6.31 1.275 ;
      RECT 6.14 1.785 6.31 1.955 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.9 1.445 9.07 1.615 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
    LAYER met1 ;
      RECT 0.55 0.735 0.84 0.78 ;
      RECT 0.55 0.78 3.13 0.92 ;
      RECT 0.55 0.92 0.84 0.965 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 6.37 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.4 1.755 2.69 1.8 ;
      RECT 2.4 1.94 2.69 1.985 ;
      RECT 2.84 0.735 3.13 0.78 ;
      RECT 2.84 0.92 3.13 0.965 ;
      RECT 2.935 0.965 3.13 1.12 ;
      RECT 2.935 1.12 6.37 1.26 ;
      RECT 5.62 1.415 5.91 1.46 ;
      RECT 5.62 1.46 9.13 1.6 ;
      RECT 5.62 1.6 5.91 1.645 ;
      RECT 6.08 1.075 6.37 1.12 ;
      RECT 6.08 1.26 6.37 1.305 ;
      RECT 6.08 1.755 6.37 1.8 ;
      RECT 6.08 1.94 6.37 1.985 ;
      RECT 8.84 1.415 9.13 1.46 ;
      RECT 8.84 1.6 9.13 1.645 ;
  END
END sky130_fd_sc_hd__dfbbn_2
MACRO sky130_fd_sc_hd__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.745 1.005 2.155 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615 0.255 11.875 0.825 ;
        RECT 11.615 1.455 11.875 2.465 ;
        RECT 11.665 0.825 11.875 1.455 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.2 0.255 10.485 0.715 ;
        RECT 10.2 1.63 10.485 2.465 ;
        RECT 10.305 0.715 10.485 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.235 1.095 9.69 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.585 0.735 3.995 0.965 ;
        RECT 3.585 0.965 3.915 1.065 ;
      LAYER mcon ;
        RECT 3.825 0.765 3.995 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.28 0.735 7.825 1.065 ;
      LAYER mcon ;
        RECT 7.575 0.765 7.745 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.805 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 7.515 0.735 7.805 0.78 ;
        RECT 7.515 0.92 7.805 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.15 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 1.405 0.635 2.125 0.825 ;
      RECT 1.405 0.825 1.575 1.795 ;
      RECT 1.405 1.795 2.125 1.965 ;
      RECT 1.43 0.085 1.785 0.465 ;
      RECT 1.43 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.325 0.705 2.545 1.575 ;
      RECT 2.325 1.575 2.825 1.955 ;
      RECT 2.335 2.25 3.165 2.42 ;
      RECT 2.4 0.265 3.415 0.465 ;
      RECT 2.725 0.645 3.075 1.015 ;
      RECT 2.995 1.195 3.415 1.235 ;
      RECT 2.995 1.235 4.345 1.405 ;
      RECT 2.995 1.405 3.165 2.25 ;
      RECT 3.245 0.465 3.415 1.195 ;
      RECT 3.335 1.575 3.585 1.785 ;
      RECT 3.335 1.785 4.685 2.035 ;
      RECT 3.405 2.205 3.785 2.635 ;
      RECT 3.585 0.085 3.755 0.525 ;
      RECT 3.925 0.255 5.075 0.425 ;
      RECT 3.925 0.425 4.255 0.505 ;
      RECT 4.085 2.035 4.255 2.375 ;
      RECT 4.095 1.405 4.345 1.485 ;
      RECT 4.125 1.155 4.345 1.235 ;
      RECT 4.405 0.595 4.735 0.765 ;
      RECT 4.515 0.765 4.735 0.895 ;
      RECT 4.515 0.895 5.825 1.065 ;
      RECT 4.515 1.065 4.685 1.785 ;
      RECT 4.855 1.235 5.185 1.415 ;
      RECT 4.855 1.415 5.86 1.655 ;
      RECT 4.875 1.915 5.205 2.635 ;
      RECT 4.905 0.425 5.075 0.715 ;
      RECT 5.325 0.085 5.675 0.465 ;
      RECT 5.495 1.065 5.825 1.235 ;
      RECT 6.06 1.575 6.295 1.985 ;
      RECT 6.065 1.06 6.405 1.125 ;
      RECT 6.065 1.125 6.74 1.305 ;
      RECT 6.185 0.705 6.405 1.06 ;
      RECT 6.25 2.25 7.08 2.42 ;
      RECT 6.3 0.265 7.08 0.465 ;
      RECT 6.535 1.305 6.74 1.905 ;
      RECT 6.91 0.465 7.08 1.235 ;
      RECT 6.91 1.235 8.26 1.405 ;
      RECT 6.91 1.405 7.08 2.25 ;
      RECT 7.25 0.085 7.575 0.525 ;
      RECT 7.25 1.575 7.5 1.915 ;
      RECT 7.25 1.915 10.03 2.085 ;
      RECT 7.32 2.255 7.7 2.635 ;
      RECT 7.745 0.255 8.955 0.425 ;
      RECT 7.745 0.425 8.075 0.545 ;
      RECT 7.94 2.085 8.11 2.375 ;
      RECT 8.04 1.075 8.26 1.235 ;
      RECT 8.215 0.665 8.615 0.835 ;
      RECT 8.43 0.835 8.615 0.84 ;
      RECT 8.43 0.84 8.6 1.915 ;
      RECT 8.64 2.255 10.03 2.635 ;
      RECT 8.77 1.11 9.055 1.575 ;
      RECT 8.77 1.575 9.555 1.745 ;
      RECT 8.785 0.425 8.955 0.585 ;
      RECT 8.835 0.755 9.475 0.925 ;
      RECT 8.835 0.925 9.055 1.11 ;
      RECT 9.265 0.265 9.475 0.755 ;
      RECT 9.725 0.085 10.03 0.805 ;
      RECT 9.86 0.995 10.125 1.325 ;
      RECT 9.86 1.325 10.03 1.915 ;
      RECT 10.66 0.255 10.975 0.995 ;
      RECT 10.66 0.995 11.495 1.325 ;
      RECT 10.66 1.325 10.975 2.415 ;
      RECT 11.15 0.085 11.445 0.545 ;
      RECT 11.155 1.765 11.445 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 0.765 0.78 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 1.105 6.295 1.275 ;
      RECT 6.125 1.785 6.295 1.955 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.855 1.445 9.025 1.615 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
    LAYER met1 ;
      RECT 0.55 0.735 0.84 0.78 ;
      RECT 0.55 0.78 3.135 0.92 ;
      RECT 0.55 0.92 0.84 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 6.355 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 6.355 1.26 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.46 9.085 1.6 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.065 1.075 6.355 1.12 ;
      RECT 6.065 1.26 6.355 1.305 ;
      RECT 6.065 1.755 6.355 1.8 ;
      RECT 6.065 1.94 6.355 1.985 ;
      RECT 8.795 1.415 9.085 1.46 ;
      RECT 8.795 1.6 9.085 1.645 ;
  END
END sky130_fd_sc_hd__dfbbn_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.615 1.32 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.075 4.7 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.34 0.28 7.6 0.735 ;
        RECT 7.34 0.735 14.085 0.905 ;
        RECT 7.375 1.495 14.085 1.72 ;
        RECT 7.375 1.72 12.745 1.735 ;
        RECT 7.375 1.735 7.6 2.46 ;
        RECT 8.2 0.28 8.46 0.735 ;
        RECT 8.2 1.735 8.46 2.46 ;
        RECT 9.06 0.28 9.32 0.735 ;
        RECT 9.06 1.735 9.32 2.46 ;
        RECT 9.905 0.28 10.18 0.735 ;
        RECT 9.92 1.735 10.18 2.46 ;
        RECT 10.765 0.28 11.025 0.735 ;
        RECT 10.765 1.735 11.025 2.46 ;
        RECT 11.625 0.28 11.885 0.735 ;
        RECT 11.625 1.735 11.885 2.46 ;
        RECT 12.485 0.28 12.745 0.735 ;
        RECT 12.485 1.735 12.745 2.46 ;
        RECT 12.92 0.905 14.085 1.495 ;
        RECT 13.355 0.28 13.615 0.735 ;
        RECT 13.355 1.72 13.645 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 10.35 1.905 10.595 2.465 ;
      LAYER mcon ;
        RECT 10.395 2.125 10.565 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.21 1.905 11.455 2.465 ;
      LAYER mcon ;
        RECT 11.255 2.125 11.425 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.07 1.905 12.315 2.465 ;
      LAYER mcon ;
        RECT 12.11 2.125 12.28 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.93 1.905 13.185 2.465 ;
      LAYER mcon ;
        RECT 12.96 2.125 13.13 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.815 1.89 14.085 2.465 ;
      LAYER mcon ;
        RECT 13.84 2.125 14.01 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.155 1.495 5.485 2.465 ;
      LAYER mcon ;
        RECT 5.235 2.125 5.405 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.015 1.495 6.345 2.465 ;
      LAYER mcon ;
        RECT 6.095 2.125 6.265 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.875 1.495 7.205 2.465 ;
      LAYER mcon ;
        RECT 6.95 2.125 7.12 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.77 1.905 8.03 2.465 ;
      LAYER mcon ;
        RECT 7.8 2.125 7.97 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.63 1.905 8.89 2.465 ;
      LAYER mcon ;
        RECT 8.68 2.125 8.85 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.49 1.905 9.75 2.465 ;
      LAYER mcon ;
        RECT 9.54 2.125 9.71 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 14.19 2.34 ;
        RECT 5.175 2.08 5.465 2.14 ;
        RECT 6.035 2.08 6.325 2.14 ;
        RECT 6.89 2.08 7.18 2.14 ;
        RECT 7.74 2.08 8.03 2.14 ;
        RECT 8.62 2.08 8.91 2.14 ;
        RECT 9.48 2.08 9.77 2.14 ;
        RECT 10.335 2.08 10.625 2.14 ;
        RECT 11.195 2.08 11.485 2.14 ;
        RECT 12.05 2.08 12.34 2.14 ;
        RECT 12.9 2.08 13.19 2.14 ;
        RECT 13.78 2.08 14.07 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
    PORT
      LAYER pwell ;
        RECT 5.205 -0.085 5.375 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 14.45 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.26 0.085 ;
      RECT 0 2.635 14.26 2.805 ;
      RECT 0.13 1.495 0.535 2.635 ;
      RECT 0.245 0.085 0.535 0.905 ;
      RECT 0.705 0.255 1.035 0.815 ;
      RECT 0.705 1.575 1.035 2.465 ;
      RECT 0.785 0.815 1.035 1.075 ;
      RECT 0.785 1.075 2.265 1.275 ;
      RECT 0.785 1.275 1.035 1.575 ;
      RECT 1.205 1.575 1.585 2.295 ;
      RECT 1.205 2.295 3.265 2.465 ;
      RECT 1.215 0.085 1.505 0.905 ;
      RECT 1.675 0.255 2.005 0.725 ;
      RECT 1.675 0.725 4.525 0.905 ;
      RECT 1.755 1.445 2.765 1.745 ;
      RECT 1.755 1.745 1.925 2.125 ;
      RECT 2.095 1.935 2.425 2.295 ;
      RECT 2.175 0.085 2.345 0.555 ;
      RECT 2.435 0.905 3.095 0.965 ;
      RECT 2.435 0.965 2.765 1.445 ;
      RECT 2.515 0.255 2.845 0.725 ;
      RECT 2.595 1.745 2.765 2.125 ;
      RECT 2.935 1.455 4.975 1.665 ;
      RECT 2.935 1.665 3.265 2.295 ;
      RECT 3.015 0.085 3.185 0.555 ;
      RECT 3.355 0.255 3.685 0.725 ;
      RECT 3.435 1.835 3.685 2.635 ;
      RECT 3.855 0.085 4.025 0.555 ;
      RECT 3.855 1.665 4.025 2.465 ;
      RECT 4.195 0.255 4.525 0.725 ;
      RECT 4.195 1.835 4.525 2.635 ;
      RECT 4.695 0.085 5.45 0.565 ;
      RECT 4.695 0.565 4.975 0.905 ;
      RECT 4.695 1.665 4.975 2.465 ;
      RECT 5.145 0.735 5.46 1.325 ;
      RECT 5.655 0.265 5.88 1.075 ;
      RECT 5.655 1.075 12.75 1.325 ;
      RECT 5.655 1.325 5.845 2.465 ;
      RECT 6.05 0.085 6.31 0.61 ;
      RECT 6.49 0.265 6.74 1.075 ;
      RECT 6.515 1.325 6.705 2.46 ;
      RECT 6.91 0.085 7.17 0.645 ;
      RECT 7.77 0.085 8.03 0.565 ;
      RECT 8.63 0.085 8.89 0.565 ;
      RECT 9.49 0.085 9.735 0.565 ;
      RECT 10.35 0.085 10.595 0.565 ;
      RECT 11.205 0.085 11.455 0.565 ;
      RECT 12.065 0.085 12.315 0.565 ;
      RECT 12.925 0.085 13.185 0.565 ;
      RECT 13.785 0.085 14.085 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.525 0.765 2.695 0.935 ;
      RECT 2.885 0.765 3.055 0.935 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.21 0.765 5.38 0.935 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
    LAYER met1 ;
      RECT 2.465 0.735 3.115 0.78 ;
      RECT 2.465 0.78 5.44 0.92 ;
      RECT 2.465 0.92 3.115 0.965 ;
      RECT 5.15 0.735 5.44 0.78 ;
      RECT 5.15 0.92 5.44 0.965 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
MACRO sky130_fd_sc_hd__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915 0.255 14.175 0.825 ;
        RECT 13.915 1.605 14.175 2.465 ;
        RECT 13.965 0.825 14.175 1.605 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.5 0.255 12.785 0.715 ;
        RECT 12.5 1.63 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.99 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.025 1.72 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 0.345 2.18 0.845 ;
        RECT 1.96 0.845 2.415 1.015 ;
        RECT 1.96 1.015 2.18 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 5.885 0.965 6.215 1.065 ;
      LAYER mcon ;
        RECT 6.125 0.765 6.295 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
      LAYER mcon ;
        RECT 9.805 0.765 9.975 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 14.45 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.26 0.085 ;
      RECT 0 2.635 14.26 2.805 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.835 0.805 ;
      RECT 0.17 1.795 0.835 1.965 ;
      RECT 0.17 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.455 0.085 1.705 0.635 ;
      RECT 1.455 1.885 1.785 2.635 ;
      RECT 2.235 1.875 2.565 2.385 ;
      RECT 2.35 0.265 2.755 0.595 ;
      RECT 2.35 1.185 3.075 1.365 ;
      RECT 2.35 1.365 2.565 1.875 ;
      RECT 2.585 0.595 2.755 1.075 ;
      RECT 2.585 1.075 3.075 1.185 ;
      RECT 2.745 1.575 3.645 1.745 ;
      RECT 2.745 1.745 3.065 1.905 ;
      RECT 2.895 1.905 3.065 2.465 ;
      RECT 2.925 0.305 3.125 0.625 ;
      RECT 2.925 0.625 3.645 0.765 ;
      RECT 2.925 0.765 3.77 0.795 ;
      RECT 3.31 2.215 3.64 2.635 ;
      RECT 3.37 0.085 3.7 0.445 ;
      RECT 3.475 0.795 3.77 1.095 ;
      RECT 3.475 1.095 3.645 1.575 ;
      RECT 4.23 0.305 4.455 2.465 ;
      RECT 4.625 0.705 4.845 1.575 ;
      RECT 4.625 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 4.7 0.265 5.715 0.465 ;
      RECT 5.025 0.645 5.375 1.015 ;
      RECT 5.295 1.195 5.715 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.545 0.465 5.715 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 5.705 2.205 6.085 2.635 ;
      RECT 5.885 0.085 6.055 0.525 ;
      RECT 6.225 0.255 7.395 0.425 ;
      RECT 6.225 0.425 6.555 0.465 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.7 0.595 7.03 0.765 ;
      RECT 6.815 0.765 7.03 0.895 ;
      RECT 6.815 0.895 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.175 1.915 7.505 2.635 ;
      RECT 7.2 0.425 7.395 0.715 ;
      RECT 7.64 0.085 7.975 0.465 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.33 2.085 ;
      RECT 9.56 0.085 9.82 0.525 ;
      RECT 9.62 2.255 10 2.635 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.43 0.465 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.575 0.645 10.905 0.815 ;
      RECT 10.73 0.815 10.905 1.915 ;
      RECT 10.94 2.255 12.33 2.635 ;
      RECT 11.075 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.765 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.855 1.745 ;
      RECT 11.565 0.265 11.765 0.755 ;
      RECT 12 0.085 12.33 0.805 ;
      RECT 12.16 0.995 12.425 1.325 ;
      RECT 12.16 1.325 12.33 1.915 ;
      RECT 12.96 0.255 13.275 0.995 ;
      RECT 12.96 0.995 13.795 1.325 ;
      RECT 12.96 1.325 13.275 2.415 ;
      RECT 13.45 1.765 13.745 2.635 ;
      RECT 13.455 0.085 13.745 0.545 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 1.785 0.775 1.955 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 1.445 11.355 1.615 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
    LAYER met1 ;
      RECT 0.545 1.755 0.835 1.8 ;
      RECT 0.545 1.8 8.655 1.94 ;
      RECT 0.545 1.94 0.835 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 5.435 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.515 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.22 0.965 5.435 1.12 ;
      RECT 5.22 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbp_1
MACRO sky130_fd_sc_hd__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.77 1.075 1.22 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.38 1.29 0.735 ;
        RECT 1.07 0.735 1.565 0.905 ;
        RECT 1.39 0.905 1.565 1.1 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 1.075 3.595 1.645 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.52 1.075 3.08 1.325 ;
        RECT 2.905 1.325 3.08 2.425 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.825 ;
        RECT 0.085 0.825 0.26 1.795 ;
        RECT 0.085 1.795 0.345 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.43 0.995 0.6 1.445 ;
      RECT 0.43 1.445 0.825 1.615 ;
      RECT 0.515 2.235 0.845 2.635 ;
      RECT 0.62 0.085 0.79 0.75 ;
      RECT 0.655 1.615 0.825 1.885 ;
      RECT 0.655 1.885 2.735 2.055 ;
      RECT 0.995 1.495 2.01 1.715 ;
      RECT 1.46 0.395 1.905 0.565 ;
      RECT 1.715 2.235 2.115 2.635 ;
      RECT 1.735 0.565 1.905 1.355 ;
      RECT 1.735 1.355 2.01 1.495 ;
      RECT 2.075 0.32 2.325 0.69 ;
      RECT 2.155 0.69 2.325 1.075 ;
      RECT 2.155 1.075 2.35 1.245 ;
      RECT 2.18 1.245 2.35 1.495 ;
      RECT 2.18 1.495 2.735 1.885 ;
      RECT 2.405 2.055 2.735 2.29 ;
      RECT 2.495 0.32 2.745 0.725 ;
      RECT 2.495 0.725 3.595 0.905 ;
      RECT 2.915 0.085 3.085 0.555 ;
      RECT 3.25 1.815 3.595 2.635 ;
      RECT 3.255 0.32 3.595 0.725 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o2bb2a_1
MACRO sky130_fd_sc_hd__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.215 1.075 1.685 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 0.38 1.735 0.735 ;
        RECT 1.515 0.735 2.02 0.77 ;
        RECT 1.515 0.77 2.025 0.905 ;
        RECT 1.855 0.905 2.025 1.1 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.7 1.075 4.045 1.645 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.075 3.525 1.325 ;
        RECT 3.355 1.325 3.525 2.425 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.87 0.825 ;
        RECT 0.535 0.825 0.705 1.795 ;
        RECT 0.535 1.795 0.79 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135 -0.085 0.305 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.11 0.085 0.365 0.91 ;
      RECT 0.11 1.41 0.365 2.635 ;
      RECT 0.875 0.995 1.045 1.445 ;
      RECT 0.875 1.445 1.27 1.615 ;
      RECT 0.96 2.235 1.29 2.635 ;
      RECT 1.065 0.085 1.235 0.75 ;
      RECT 1.1 1.615 1.27 1.885 ;
      RECT 1.1 1.885 3.185 2.055 ;
      RECT 1.44 1.495 2.46 1.715 ;
      RECT 1.905 0.395 2.365 0.565 ;
      RECT 2.16 2.235 2.565 2.635 ;
      RECT 2.195 0.565 2.365 1.355 ;
      RECT 2.195 1.355 2.46 1.495 ;
      RECT 2.535 0.32 2.78 0.69 ;
      RECT 2.61 0.69 2.78 1.075 ;
      RECT 2.61 1.075 2.8 1.245 ;
      RECT 2.63 1.245 2.8 1.495 ;
      RECT 2.63 1.495 3.185 1.885 ;
      RECT 2.835 2.055 3.185 2.425 ;
      RECT 2.955 0.32 3.185 0.725 ;
      RECT 2.955 0.725 4.045 0.905 ;
      RECT 3.375 0.085 3.545 0.555 ;
      RECT 3.715 0.32 4.045 0.725 ;
      RECT 3.73 1.815 4.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o2bb2a_2
MACRO sky130_fd_sc_hd__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.075 3.645 1.445 ;
        RECT 3.315 1.445 4.965 1.615 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 0.085 1.445 1.895 1.615 ;
        RECT 1.565 1.075 1.895 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 5.235 0.725 6.91 0.905 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.075 0.275 6.405 0.725 ;
        RECT 6.115 1.415 6.91 1.655 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 6.605 0.905 6.91 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.095 0.255 0.425 0.725 ;
      RECT 0.095 0.725 1.265 0.735 ;
      RECT 0.095 0.735 2.025 0.905 ;
      RECT 0.14 1.795 0.345 2.635 ;
      RECT 0.555 1.785 0.805 2.295 ;
      RECT 0.555 2.295 1.645 2.465 ;
      RECT 0.595 0.085 0.765 0.555 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 0.975 1.785 2.615 1.955 ;
      RECT 0.975 1.955 1.225 2.125 ;
      RECT 1.395 2.125 1.645 2.295 ;
      RECT 1.435 0.085 1.605 0.555 ;
      RECT 1.775 0.255 2.945 0.475 ;
      RECT 1.775 0.475 2.025 0.735 ;
      RECT 1.815 2.125 2.065 2.635 ;
      RECT 2.065 1.075 2.445 1.415 ;
      RECT 2.065 1.415 2.615 1.785 ;
      RECT 2.195 0.645 2.525 0.815 ;
      RECT 2.195 0.815 2.445 1.075 ;
      RECT 2.235 1.955 2.615 1.965 ;
      RECT 2.235 1.965 2.525 2.465 ;
      RECT 2.615 1.075 3.145 1.245 ;
      RECT 2.695 2.135 3.425 2.635 ;
      RECT 2.955 0.725 4.305 0.905 ;
      RECT 2.955 0.905 3.145 1.075 ;
      RECT 2.955 1.245 3.145 1.785 ;
      RECT 2.955 1.785 4.685 1.965 ;
      RECT 3.215 0.085 3.385 0.555 ;
      RECT 3.555 0.305 4.725 0.475 ;
      RECT 3.595 1.965 3.845 2.125 ;
      RECT 3.975 0.645 4.305 0.725 ;
      RECT 4.015 2.135 4.265 2.635 ;
      RECT 4.435 1.965 4.685 2.465 ;
      RECT 4.475 0.475 4.725 0.895 ;
      RECT 4.855 1.795 5.105 2.635 ;
      RECT 4.895 0.085 5.065 0.895 ;
      RECT 5.165 1.075 6.435 1.245 ;
      RECT 5.165 1.245 5.455 1.615 ;
      RECT 5.695 2.165 5.945 2.635 ;
      RECT 5.735 0.085 5.905 0.555 ;
      RECT 6.535 1.825 6.785 2.635 ;
      RECT 6.575 0.085 6.745 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.445 2.615 1.615 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.225 1.445 5.395 1.615 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
    LAYER met1 ;
      RECT 2.385 1.415 2.675 1.46 ;
      RECT 2.385 1.46 5.455 1.6 ;
      RECT 2.385 1.6 2.675 1.645 ;
      RECT 5.165 1.415 5.455 1.46 ;
      RECT 5.165 1.6 5.455 1.645 ;
  END
END sky130_fd_sc_hd__o2bb2a_4
MACRO sky130_fd_sc_hd__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 0.415 5.435 0.745 ;
        RECT 5.15 1.67 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.67 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.77 2.255 3.605 2.425 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.175 1.165 ;
      RECT 3.435 1.165 4.175 1.325 ;
      RECT 3.435 1.325 3.605 2.255 ;
      RECT 3.685 0.085 4.015 0.53 ;
      RECT 3.775 2.135 3.945 2.635 ;
      RECT 3.84 1.535 4.515 1.865 ;
      RECT 4.295 0.415 4.515 0.745 ;
      RECT 4.295 1.865 4.515 2.435 ;
      RECT 4.345 0.745 4.515 0.995 ;
      RECT 4.345 0.995 5.095 1.325 ;
      RECT 4.345 1.325 4.515 1.535 ;
      RECT 4.695 0.085 4.9 0.715 ;
      RECT 4.695 1.57 4.9 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.785 3.1 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.16 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
  END
END sky130_fd_sc_hd__dlxtp_1
MACRO sky130_fd_sc_hd__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.33 1.655 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 0.995 1.245 1.325 ;
        RECT 0.89 0.42 1.245 0.995 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.425 1.7 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905 0.73 2.155 0.935 ;
        RECT 1.905 0.935 2.075 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535 0.255 2.705 0.64 ;
        RECT 2.535 0.64 4.05 0.81 ;
        RECT 2.535 1.795 2.785 2.465 ;
        RECT 2.615 1.485 4.05 1.655 ;
        RECT 2.615 1.655 2.785 1.795 ;
        RECT 3.375 0.255 3.545 0.64 ;
        RECT 3.375 1.655 4.05 1.745 ;
        RECT 3.375 1.745 3.545 2.465 ;
        RECT 3.8 0.81 4.05 1.485 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.105 1.835 0.385 2.635 ;
      RECT 0.175 0.255 0.67 0.585 ;
      RECT 0.5 0.585 0.67 1.495 ;
      RECT 0.5 1.495 2.415 1.665 ;
      RECT 0.555 1.665 0.765 2.465 ;
      RECT 0.955 1.935 1.285 2.635 ;
      RECT 1.455 1.665 1.645 2.465 ;
      RECT 2.025 0.085 2.335 0.55 ;
      RECT 2.025 1.855 2.355 2.635 ;
      RECT 2.245 1.105 3.585 1.305 ;
      RECT 2.245 1.305 2.415 1.495 ;
      RECT 2.575 1.075 3.585 1.105 ;
      RECT 2.875 0.085 3.205 0.47 ;
      RECT 2.955 1.835 3.205 2.635 ;
      RECT 3.715 0.085 4.045 0.47 ;
      RECT 3.715 1.915 4.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__and4_4
MACRO sky130_fd_sc_hd__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.755 0.33 2.075 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.89 0.42 1.245 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.415 1.72 1.305 ;
        RECT 1.42 1.305 1.59 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.9 0.415 2.16 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 0.295 3.065 0.34 ;
        RECT 2.735 0.34 3.07 0.805 ;
        RECT 2.735 1.495 3.07 2.465 ;
        RECT 2.895 0.805 3.07 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.095 2.255 0.425 2.635 ;
      RECT 0.175 0.255 0.67 0.585 ;
      RECT 0.5 0.585 0.67 1.495 ;
      RECT 0.5 1.495 2.555 1.665 ;
      RECT 0.6 1.665 0.85 2.465 ;
      RECT 1.07 1.915 1.4 2.635 ;
      RECT 1.585 1.665 1.835 2.465 ;
      RECT 2.235 1.835 2.565 2.635 ;
      RECT 2.33 0.085 2.565 0.89 ;
      RECT 2.33 1.075 2.725 1.315 ;
      RECT 2.33 1.315 2.555 1.495 ;
      RECT 3.245 1.835 3.575 2.635 ;
      RECT 3.255 0.085 3.585 0.81 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__and4_2
MACRO sky130_fd_sc_hd__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.325 2.075 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885 0.36 1.235 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.355 1.715 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.355 2.175 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795 0.295 3.135 0.805 ;
        RECT 2.795 2.205 3.135 2.465 ;
        RECT 2.875 0.805 3.135 2.205 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 2.255 0.425 2.635 ;
      RECT 0.17 0.255 0.665 0.585 ;
      RECT 0.495 0.585 0.665 1.495 ;
      RECT 0.495 1.495 2.685 1.665 ;
      RECT 0.595 1.665 0.845 2.465 ;
      RECT 1.065 1.915 1.395 2.635 ;
      RECT 1.58 1.665 1.83 2.465 ;
      RECT 2.295 1.835 2.625 2.635 ;
      RECT 2.355 0.085 2.625 0.885 ;
      RECT 2.37 1.075 2.7 1.325 ;
      RECT 2.37 1.325 2.685 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__and4_1
MACRO sky130_fd_sc_hd__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.955 2.985 1.325 ;
        RECT 2.755 0.415 3.105 0.61 ;
        RECT 2.755 0.61 2.985 0.955 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.165 0.995 3.545 1.325 ;
        RECT 3.305 0.425 3.545 0.995 ;
        RECT 3.305 1.325 3.545 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.995 4.055 1.63 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085 1.075 2.515 1.245 ;
        RECT 2.345 1.245 2.515 1.445 ;
        RECT 2.345 1.445 2.55 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.745 1.53 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.695500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.655 0.845 0.825 ;
        RECT 0.135 0.825 0.345 1.785 ;
        RECT 0.135 1.785 1.185 1.955 ;
        RECT 0.135 1.955 0.345 2.465 ;
        RECT 1.015 1.955 1.185 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.085 0.425 0.465 ;
      RECT 0.515 2.125 0.845 2.635 ;
      RECT 0.535 0.995 0.705 1.445 ;
      RECT 0.535 1.445 2.125 1.615 ;
      RECT 0.935 0.085 1.64 0.445 ;
      RECT 1.535 1.785 1.705 2.295 ;
      RECT 1.535 2.295 2.545 2.465 ;
      RECT 1.7 0.615 2.585 0.785 ;
      RECT 1.7 0.785 1.89 1.445 ;
      RECT 1.875 1.615 2.125 1.945 ;
      RECT 1.875 1.945 2.205 2.115 ;
      RECT 2.255 0.275 2.585 0.615 ;
      RECT 2.375 1.795 3.545 1.965 ;
      RECT 2.375 1.965 2.545 2.295 ;
      RECT 2.715 2.14 3.045 2.635 ;
      RECT 3.375 1.965 3.545 2.465 ;
      RECT 3.715 0.085 4.05 0.805 ;
      RECT 3.715 1.915 4.05 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a32o_2
MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.28 1.075 5.075 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.075 4.03 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 3.105 1.295 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.63 1.075 6.78 1.625 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.03 1.075 7.71 1.295 ;
        RECT 7.03 1.295 7.225 1.635 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.635 1.605 0.805 ;
        RECT 0.12 0.805 0.34 1.495 ;
        RECT 0.12 1.495 1.605 1.665 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 1.665 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.435 1.665 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 0.095 1.915 0.425 2.635 ;
      RECT 0.57 0.995 1.97 1.325 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 0.935 1.915 1.265 2.635 ;
      RECT 1.775 0.085 2.105 0.465 ;
      RECT 1.775 1.915 2.105 2.635 ;
      RECT 1.8 1.325 1.97 1.495 ;
      RECT 1.8 1.495 5.45 1.665 ;
      RECT 2.275 0.255 2.445 0.655 ;
      RECT 2.275 0.655 3.885 0.825 ;
      RECT 2.275 1.915 5.065 2.085 ;
      RECT 2.275 2.085 2.445 2.465 ;
      RECT 2.615 0.085 2.945 0.465 ;
      RECT 2.615 2.255 2.945 2.635 ;
      RECT 3.135 0.295 5.145 0.465 ;
      RECT 3.215 2.085 3.385 2.465 ;
      RECT 3.555 2.255 3.885 2.635 ;
      RECT 4.055 2.085 4.225 2.465 ;
      RECT 4.395 0.635 6.425 0.805 ;
      RECT 4.395 2.255 4.725 2.635 ;
      RECT 4.895 2.085 5.065 2.255 ;
      RECT 4.895 2.255 7.725 2.425 ;
      RECT 5.28 0.805 5.45 1.495 ;
      RECT 5.28 1.665 5.45 1.905 ;
      RECT 5.28 1.905 6.2 1.915 ;
      RECT 5.28 1.915 7.305 2.075 ;
      RECT 5.67 0.295 6.805 0.465 ;
      RECT 6.135 2.075 7.305 2.085 ;
      RECT 6.635 0.255 6.805 0.295 ;
      RECT 6.635 0.465 6.805 0.645 ;
      RECT 6.635 0.645 7.645 0.815 ;
      RECT 6.975 0.085 7.305 0.465 ;
      RECT 7.475 0.255 7.645 0.645 ;
      RECT 7.475 1.755 7.725 2.255 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__a32o_4
MACRO sky130_fd_sc_hd__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.665 2.28 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.665 1.8 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.995 1.32 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.66 2.87 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.18 0.995 3.53 1.325 ;
        RECT 3.325 1.325 3.53 1.615 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.3 0.425 0.56 ;
        RECT 0.09 0.56 0.345 1.915 ;
        RECT 0.09 1.915 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.57 0.995 0.875 1.325 ;
      RECT 0.595 0.085 0.925 0.485 ;
      RECT 0.675 1.835 1.005 2.635 ;
      RECT 0.705 0.655 1.265 0.825 ;
      RECT 0.705 0.825 0.875 0.995 ;
      RECT 0.705 1.325 0.875 1.495 ;
      RECT 0.705 1.495 3.075 1.665 ;
      RECT 1.095 0.315 2.71 0.485 ;
      RECT 1.095 0.485 1.265 0.655 ;
      RECT 1.25 1.875 2.675 2.045 ;
      RECT 1.25 2.045 1.535 2.465 ;
      RECT 1.79 2.215 2.12 2.635 ;
      RECT 2.345 2.045 2.675 2.295 ;
      RECT 2.345 2.295 3.505 2.465 ;
      RECT 2.905 1.665 3.075 2.125 ;
      RECT 3.255 0.085 3.585 0.805 ;
      RECT 3.335 1.795 3.505 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a32o_1
MACRO sky130_fd_sc_hd__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.075 3.995 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.075 3.275 2.39 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 2.735 2.39 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865 1.075 2.195 2.39 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.075 1.695 1.285 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.672000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.885 ;
        RECT 0.085 0.885 0.355 1.455 ;
        RECT 0.085 1.455 0.61 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.525 1.075 1.105 1.285 ;
      RECT 0.715 0.085 0.885 0.545 ;
      RECT 0.735 0.715 1.485 0.905 ;
      RECT 0.735 0.905 1.105 1.075 ;
      RECT 0.845 1.285 1.105 1.455 ;
      RECT 0.845 1.455 1.595 1.745 ;
      RECT 0.845 1.915 1.175 2.635 ;
      RECT 1.155 0.27 1.485 0.715 ;
      RECT 1.345 1.745 1.595 2.465 ;
      RECT 1.655 0.415 1.825 0.735 ;
      RECT 1.655 0.735 3.955 0.905 ;
      RECT 2.05 0.085 2.38 0.545 ;
      RECT 2.58 0.255 2.91 0.735 ;
      RECT 3.125 0.085 3.455 0.545 ;
      RECT 3.605 1.515 3.935 2.635 ;
      RECT 3.625 0.255 3.955 0.735 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o41a_1
MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.65 1.075 7.735 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 1.075 6.36 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.33 1.075 4.96 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.41 1.075 4.04 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.165 1.275 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 1.685 0.905 ;
        RECT 0.085 0.905 0.345 1.465 ;
        RECT 0.085 1.465 1.685 1.665 ;
        RECT 0.515 0.255 0.845 0.715 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 0.255 1.685 0.715 ;
        RECT 1.355 1.665 1.685 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.085 0.085 0.345 0.545 ;
      RECT 0.085 1.835 0.345 2.635 ;
      RECT 0.515 1.075 2.665 1.245 ;
      RECT 0.515 1.245 2.545 1.295 ;
      RECT 1.015 0.085 1.185 0.545 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.855 0.085 2.105 0.885 ;
      RECT 1.855 1.465 2.025 2.635 ;
      RECT 2.195 1.295 2.545 1.445 ;
      RECT 2.195 1.445 3.825 1.615 ;
      RECT 2.195 1.615 2.545 2.465 ;
      RECT 2.295 0.255 3.485 0.465 ;
      RECT 2.295 0.635 3.045 0.905 ;
      RECT 2.295 0.905 2.665 1.075 ;
      RECT 2.715 1.835 2.965 2.635 ;
      RECT 3.135 1.835 3.405 2.295 ;
      RECT 3.135 2.295 4.325 2.465 ;
      RECT 3.235 0.465 3.485 0.735 ;
      RECT 3.235 0.735 7.595 0.905 ;
      RECT 3.575 1.615 3.825 2.125 ;
      RECT 3.655 0.085 3.875 0.545 ;
      RECT 3.995 1.445 5.165 1.615 ;
      RECT 3.995 1.615 4.325 2.295 ;
      RECT 4.075 0.255 4.245 0.735 ;
      RECT 4.445 0.085 4.715 0.545 ;
      RECT 4.495 1.785 4.665 2.295 ;
      RECT 4.495 2.295 6.145 2.465 ;
      RECT 4.835 1.615 5.165 2.115 ;
      RECT 4.915 0.255 5.085 0.735 ;
      RECT 5.305 0.085 5.915 0.545 ;
      RECT 5.395 1.445 7.595 1.615 ;
      RECT 5.395 1.615 5.645 2.115 ;
      RECT 5.815 1.785 6.145 2.295 ;
      RECT 6.24 0.255 6.41 0.735 ;
      RECT 6.315 1.615 6.485 2.455 ;
      RECT 6.655 1.785 6.985 2.635 ;
      RECT 6.685 0.085 6.955 0.545 ;
      RECT 7.265 0.255 7.595 0.735 ;
      RECT 7.265 1.615 7.595 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__o41a_4
MACRO sky130_fd_sc_hd__o41a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.515 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.075 3.655 2.335 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.825 1.075 3.155 2.34 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.075 2.655 2.34 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.155 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.88 ;
        RECT 0.515 0.88 0.79 1.495 ;
        RECT 0.515 1.495 0.845 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.085 0.345 0.885 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 0.96 1.075 1.6 1.325 ;
      RECT 1.015 0.085 1.26 0.885 ;
      RECT 1.015 1.495 1.185 1.835 ;
      RECT 1.015 1.835 1.525 2.635 ;
      RECT 1.355 1.325 1.6 1.495 ;
      RECT 1.355 1.495 2.145 1.665 ;
      RECT 1.43 0.255 1.785 0.85 ;
      RECT 1.43 0.85 1.6 1.075 ;
      RECT 1.695 1.665 2.145 2.465 ;
      RECT 1.985 0.255 2.315 0.715 ;
      RECT 1.985 0.715 4.395 0.905 ;
      RECT 2.485 0.085 2.75 0.545 ;
      RECT 2.955 0.255 3.285 0.715 ;
      RECT 3.505 0.085 3.775 0.545 ;
      RECT 4.065 0.255 4.395 0.715 ;
      RECT 4.065 1.495 4.395 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__o41a_2
MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.75 1.075 5.865 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.37 1.075 4.48 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 3.065 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.705 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.845 1.325 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 2.045 0.905 ;
        RECT 0.515 1.495 3.105 1.665 ;
        RECT 0.515 1.665 0.845 2.095 ;
        RECT 1.875 0.905 2.045 1.105 ;
        RECT 1.875 1.105 2.17 1.495 ;
        RECT 2.775 1.665 3.105 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.09 0.255 2.405 0.485 ;
      RECT 0.09 0.485 0.345 0.905 ;
      RECT 0.09 1.495 0.345 2.295 ;
      RECT 0.09 2.295 1.265 2.465 ;
      RECT 1.015 1.835 2.105 2.005 ;
      RECT 1.015 2.005 1.265 2.295 ;
      RECT 1.435 2.175 1.605 2.635 ;
      RECT 1.775 2.005 2.105 2.455 ;
      RECT 2.235 0.485 2.405 0.715 ;
      RECT 2.235 0.715 5.755 0.905 ;
      RECT 2.335 1.835 2.585 2.255 ;
      RECT 2.335 2.255 4.385 2.445 ;
      RECT 2.62 0.085 2.95 0.545 ;
      RECT 3.135 0.255 3.465 0.715 ;
      RECT 3.275 1.495 3.445 2.255 ;
      RECT 3.615 1.495 5.325 1.665 ;
      RECT 3.615 1.665 3.945 2.085 ;
      RECT 3.635 0.085 3.805 0.545 ;
      RECT 4.055 0.255 4.725 0.715 ;
      RECT 4.135 1.835 4.385 2.255 ;
      RECT 4.62 1.835 4.825 2.635 ;
      RECT 4.905 0.085 5.235 0.545 ;
      RECT 4.995 1.665 5.325 2.46 ;
      RECT 5.425 0.255 5.755 0.715 ;
      RECT 5.495 1.495 5.715 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__o32ai_2
MACRO sky130_fd_sc_hd__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.575 0.995 3.135 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.93 0.995 2.225 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 0.995 1.7 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.685 0.345 0.995 ;
        RECT 0.09 0.995 0.36 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.87 0.995 1.24 1.615 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.821250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 0.845 0.825 ;
        RECT 0.53 0.825 0.7 1.785 ;
        RECT 0.53 1.785 1.545 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 0.255 1.345 0.485 ;
      RECT 0.09 1.495 0.36 2.635 ;
      RECT 1.015 0.485 1.345 0.655 ;
      RECT 1.015 0.655 2.525 0.825 ;
      RECT 1.515 0.085 2.185 0.485 ;
      RECT 2.355 0.375 2.525 0.655 ;
      RECT 2.695 0.085 3.135 0.825 ;
      RECT 2.695 1.495 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o32ai_1
MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.29 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.09 1.075 7.26 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.77 1.075 5.38 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 3.54 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.685 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 3.38 0.905 ;
        RECT 0.515 1.495 5.58 1.665 ;
        RECT 0.515 1.665 0.845 2.085 ;
        RECT 1.355 1.665 1.7 2.085 ;
        RECT 1.855 0.905 2.035 1.495 ;
        RECT 4.41 1.665 4.74 2.085 ;
        RECT 5.25 1.665 5.58 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.09 0.255 3.8 0.465 ;
      RECT 0.09 0.465 0.345 0.905 ;
      RECT 0.09 1.495 0.345 2.255 ;
      RECT 0.09 2.255 2.04 2.465 ;
      RECT 1.015 1.835 1.185 2.255 ;
      RECT 1.87 1.835 3.8 2.005 ;
      RECT 1.87 2.005 2.04 2.255 ;
      RECT 2.21 2.175 2.54 2.635 ;
      RECT 2.71 2.005 2.88 2.425 ;
      RECT 3.05 2.175 3.38 2.635 ;
      RECT 3.55 0.465 3.8 0.735 ;
      RECT 3.55 0.735 10.035 0.905 ;
      RECT 3.55 2.005 3.8 2.465 ;
      RECT 3.97 0.085 4.14 0.545 ;
      RECT 3.99 1.835 4.24 2.255 ;
      RECT 3.99 2.255 7.68 2.465 ;
      RECT 4.31 0.255 4.64 0.735 ;
      RECT 4.81 0.085 5.14 0.545 ;
      RECT 4.91 1.835 5.08 2.255 ;
      RECT 5.31 0.255 5.98 0.735 ;
      RECT 5.75 1.835 5.92 2.255 ;
      RECT 6.09 1.495 9.46 1.665 ;
      RECT 6.09 1.665 6.42 2.085 ;
      RECT 6.17 0.085 6.34 0.545 ;
      RECT 6.51 0.255 6.84 0.735 ;
      RECT 6.59 1.835 6.76 2.255 ;
      RECT 6.93 1.665 7.26 2.085 ;
      RECT 7.01 0.085 7.18 0.545 ;
      RECT 7.35 0.255 8.04 0.735 ;
      RECT 7.43 1.835 7.68 2.255 ;
      RECT 7.87 1.835 8.12 2.635 ;
      RECT 8.29 1.665 8.62 2.465 ;
      RECT 8.37 0.085 8.54 0.545 ;
      RECT 8.71 0.255 9.04 0.735 ;
      RECT 8.79 1.835 8.96 2.635 ;
      RECT 9.13 1.665 9.46 2.465 ;
      RECT 9.21 0.085 9.47 0.545 ;
      RECT 9.63 1.495 10.035 2.635 ;
      RECT 9.645 0.255 10.035 0.735 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__o32ai_4
MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.765 1.95 1.015 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.039500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.04 0.255 6.46 0.545 ;
        RECT 6.04 1.835 7.3 2.005 ;
        RECT 6.04 2.005 6.37 2.455 ;
        RECT 6.29 0.545 6.46 0.715 ;
        RECT 6.29 0.715 7.3 0.885 ;
        RECT 6.585 1.785 7.3 1.835 ;
        RECT 6.75 0.885 7.3 1.785 ;
        RECT 6.97 0.255 7.3 0.715 ;
        RECT 6.97 2.005 7.3 2.465 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
      LAYER mcon ;
        RECT 0.15 1.105 0.32 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.23 1.055 5.74 1.325 ;
      LAYER mcon ;
        RECT 5.23 1.105 5.4 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.09 1.075 0.38 1.12 ;
        RECT 0.09 1.12 5.46 1.26 ;
        RECT 0.09 1.26 0.38 1.305 ;
        RECT 5.17 1.075 5.46 1.12 ;
        RECT 5.17 1.26 5.46 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.28 1.355 ;
      RECT 1.015 1.355 2.335 1.585 ;
      RECT 1.015 1.585 1.24 2.465 ;
      RECT 1.45 0.085 1.785 0.465 ;
      RECT 1.45 2.195 1.815 2.635 ;
      RECT 1.525 1.785 1.695 1.855 ;
      RECT 1.525 1.855 2.845 1.905 ;
      RECT 1.525 1.905 2.735 2.025 ;
      RECT 2.045 1.585 2.335 1.685 ;
      RECT 2.29 0.705 2.735 1.035 ;
      RECT 2.415 0.365 3.075 0.535 ;
      RECT 2.475 2.195 3.165 2.425 ;
      RECT 2.505 1.575 2.845 1.855 ;
      RECT 2.565 1.035 2.735 1.575 ;
      RECT 2.905 0.535 3.075 0.995 ;
      RECT 2.905 0.995 3.775 1.165 ;
      RECT 2.915 2.06 3.185 2.09 ;
      RECT 2.915 2.09 3.18 2.105 ;
      RECT 2.915 2.105 3.165 2.195 ;
      RECT 2.98 2.015 3.185 2.06 ;
      RECT 3.015 1.165 3.775 1.325 ;
      RECT 3.015 1.325 3.185 2.015 ;
      RECT 3.315 0.085 3.65 0.53 ;
      RECT 3.335 2.175 3.695 2.635 ;
      RECT 3.355 1.535 4.115 1.865 ;
      RECT 3.895 0.415 4.115 0.745 ;
      RECT 3.895 1.865 4.115 2.435 ;
      RECT 3.945 0.745 4.115 0.995 ;
      RECT 3.945 0.995 4.72 1.325 ;
      RECT 3.945 1.325 4.115 1.535 ;
      RECT 4.295 0.085 4.58 0.715 ;
      RECT 4.295 2.01 4.58 2.635 ;
      RECT 4.75 0.29 5.06 0.715 ;
      RECT 4.75 0.715 6.12 0.825 ;
      RECT 4.75 1.495 6.14 1.665 ;
      RECT 4.75 1.665 5.035 2.465 ;
      RECT 4.89 0.825 6.12 0.885 ;
      RECT 4.89 0.885 5.06 1.495 ;
      RECT 5.575 1.835 5.84 2.635 ;
      RECT 5.59 0.085 5.87 0.545 ;
      RECT 5.91 0.885 6.12 1.055 ;
      RECT 5.91 1.055 6.58 1.29 ;
      RECT 5.91 1.29 6.14 1.495 ;
      RECT 6.54 2.175 6.8 2.635 ;
      RECT 6.63 0.085 6.8 0.545 ;
      RECT 7.47 0.085 7.735 0.885 ;
      RECT 7.47 1.485 7.735 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 1.755 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.465 1.755 1.755 1.8 ;
      RECT 1.465 1.94 1.755 1.985 ;
  END
END sky130_fd_sc_hd__dlclkp_4
MACRO sky130_fd_sc_hd__dlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 1.435 2.215 1.685 ;
        RECT 1.985 0.285 2.215 1.435 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.36 0.595 ;
        RECT 6.095 1.495 6.36 2.455 ;
        RECT 6.165 0.595 6.36 1.495 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
      LAYER mcon ;
        RECT 0.15 1.105 0.32 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.21 1.105 5.485 1.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.09 1.075 0.38 1.12 ;
        RECT 0.09 1.12 5.44 1.26 ;
        RECT 0.09 1.26 0.38 1.305 ;
        RECT 5.15 1.075 5.44 1.12 ;
        RECT 5.15 1.26 5.44 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 0.995 1.355 ;
        RECT -0.19 1.355 7.09 2.91 ;
        RECT 2.625 1.305 7.09 1.355 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.175 0.26 0.345 0.615 ;
      RECT 0.175 0.615 0.78 0.785 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.785 0.78 1.06 ;
      RECT 0.61 1.06 0.84 1.39 ;
      RECT 0.61 1.39 0.78 1.795 ;
      RECT 1.015 0.26 1.28 1.855 ;
      RECT 1.015 1.855 2.645 2.025 ;
      RECT 1.015 2.025 1.24 2.465 ;
      RECT 1.455 2.195 1.82 2.635 ;
      RECT 1.485 0.085 1.815 0.905 ;
      RECT 2.395 0.815 3.225 0.985 ;
      RECT 2.395 0.985 2.645 1.855 ;
      RECT 2.48 2.255 3.23 2.425 ;
      RECT 2.795 0.39 3.725 0.56 ;
      RECT 3.06 1.155 4.18 1.325 ;
      RECT 3.06 1.325 3.23 2.255 ;
      RECT 3.4 2.135 3.7 2.635 ;
      RECT 3.435 1.535 4.735 1.84 ;
      RECT 3.435 1.84 4.135 1.865 ;
      RECT 3.555 0.56 3.725 0.995 ;
      RECT 3.555 0.995 4.18 1.155 ;
      RECT 3.895 0.085 4.145 0.61 ;
      RECT 3.915 1.865 4.135 2.435 ;
      RECT 4.315 0.255 4.585 0.615 ;
      RECT 4.315 2.01 4.6 2.635 ;
      RECT 4.35 0.615 4.585 0.995 ;
      RECT 4.35 0.995 4.735 1.535 ;
      RECT 4.835 0.29 5.15 0.62 ;
      RECT 4.93 0.62 5.15 0.765 ;
      RECT 4.93 0.765 5.995 0.935 ;
      RECT 5.01 1.725 5.925 1.895 ;
      RECT 5.01 1.895 5.34 2.465 ;
      RECT 5.575 2.13 5.925 2.635 ;
      RECT 5.675 0.085 5.845 0.545 ;
      RECT 5.755 0.935 5.995 1.325 ;
      RECT 5.755 1.325 5.925 1.725 ;
      RECT 6.53 0.085 6.81 0.885 ;
      RECT 6.53 1.485 6.81 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
  END
END sky130_fd_sc_hd__dlclkp_2
MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.435 2.185 1.685 ;
        RECT 1.985 0.385 2.185 1.435 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 0.255 6.355 0.595 ;
        RECT 6.09 1.495 6.355 2.455 ;
        RECT 6.17 0.595 6.355 1.495 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
      LAYER mcon ;
        RECT 0.145 1.105 0.315 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.19 1.105 5.51 1.435 ;
      LAYER mcon ;
        RECT 5.21 1.105 5.38 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.075 0.38 1.12 ;
        RECT 0.085 1.12 5.44 1.26 ;
        RECT 0.085 1.26 0.38 1.305 ;
        RECT 5.15 1.075 5.44 1.12 ;
        RECT 5.15 1.26 5.44 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 0.995 1.355 ;
        RECT -0.19 1.355 6.63 2.91 ;
        RECT 2.62 1.305 6.63 1.355 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.175 0.26 0.345 0.615 ;
      RECT 0.175 0.615 0.78 0.785 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.785 0.78 1.06 ;
      RECT 0.61 1.06 0.84 1.39 ;
      RECT 0.61 1.39 0.78 1.795 ;
      RECT 1.015 0.26 1.28 1.855 ;
      RECT 1.015 1.855 2.59 2.025 ;
      RECT 1.015 2.025 1.24 2.465 ;
      RECT 1.45 2.195 1.815 2.635 ;
      RECT 1.48 0.085 1.81 0.905 ;
      RECT 2.39 0.815 3.22 0.985 ;
      RECT 2.39 0.985 2.59 1.855 ;
      RECT 2.475 2.255 3.225 2.425 ;
      RECT 2.79 0.39 3.725 0.56 ;
      RECT 3.055 1.155 4.175 1.325 ;
      RECT 3.055 1.325 3.225 2.255 ;
      RECT 3.395 2.135 3.695 2.635 ;
      RECT 3.43 1.535 4.71 1.84 ;
      RECT 3.43 1.84 4.13 1.865 ;
      RECT 3.555 0.56 3.725 0.995 ;
      RECT 3.555 0.995 4.175 1.155 ;
      RECT 3.895 0.085 4.145 0.61 ;
      RECT 3.91 1.865 4.13 2.435 ;
      RECT 4.31 2.01 4.595 2.635 ;
      RECT 4.32 0.255 4.58 0.615 ;
      RECT 4.345 0.615 4.58 0.995 ;
      RECT 4.345 0.995 4.74 1.325 ;
      RECT 4.345 1.325 4.71 1.535 ;
      RECT 4.84 0.29 5.155 0.62 ;
      RECT 4.935 0.62 5.155 0.765 ;
      RECT 4.935 0.765 6 0.935 ;
      RECT 5.005 1.725 5.92 1.895 ;
      RECT 5.005 1.895 5.335 2.465 ;
      RECT 5.57 2.13 5.92 2.635 ;
      RECT 5.67 0.085 5.84 0.545 ;
      RECT 5.75 0.935 6 1.325 ;
      RECT 5.75 1.325 5.92 1.725 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__dlclkp_1
MACRO sky130_fd_sc_hd__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.16 0.265 9.495 1.695 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.03 1.535 10.42 2.08 ;
        RECT 10.04 0.31 10.42 0.825 ;
        RECT 10.12 2.08 10.42 2.465 ;
        RECT 10.25 0.825 10.42 1.535 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 7.985 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.055 2.635 ;
      RECT 7.815 0.465 7.985 0.995 ;
      RECT 7.815 0.995 8.16 1.075 ;
      RECT 7.815 1.075 8.65 1.295 ;
      RECT 7.99 1.295 8.65 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.335 0.345 8.585 0.715 ;
      RECT 8.335 0.715 8.99 0.885 ;
      RECT 8.335 1.795 8.99 1.865 ;
      RECT 8.335 1.865 9.835 2.035 ;
      RECT 8.335 2.035 8.56 2.465 ;
      RECT 8.73 2.205 9.07 2.635 ;
      RECT 8.755 0.085 8.99 0.545 ;
      RECT 8.82 0.885 8.99 1.795 ;
      RECT 9.62 2.255 9.95 2.635 ;
      RECT 9.665 0.995 10.08 1.325 ;
      RECT 9.665 1.325 9.835 1.865 ;
      RECT 9.7 0.085 9.87 0.825 ;
      RECT 10.59 0.085 10.76 0.93 ;
      RECT 10.59 1.445 10.76 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrbp_2
MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.6 1.455 9.005 2.465 ;
        RECT 8.675 0.275 9.005 1.455 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.18 0.265 10.435 0.795 ;
        RECT 10.18 1.445 10.435 2.325 ;
        RECT 10.225 0.795 10.435 1.445 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.77 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.58 0.085 ;
      RECT 0 2.635 10.58 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.43 2.635 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.435 1.295 ;
      RECT 7.99 1.295 8.435 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.335 0.085 8.505 0.77 ;
      RECT 9.195 0.345 9.445 0.995 ;
      RECT 9.195 0.995 10.055 1.325 ;
      RECT 9.195 1.325 9.525 2.425 ;
      RECT 9.76 0.085 9.93 0.68 ;
      RECT 9.76 1.495 9.93 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrbp_1
MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.4 1.075 1.41 1.33 ;
        RECT 0.965 1.33 1.41 1.515 ;
        RECT 0.965 1.515 3.63 1.685 ;
        RECT 3.35 0.995 3.63 1.515 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705 1.075 3.18 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.8 0.995 4.975 1.41 ;
        RECT 4.26 1.41 4.975 1.515 ;
        RECT 4.26 1.515 7 1.685 ;
        RECT 6.83 0.995 7 1.515 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.37 1.075 6.44 1.345 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.001000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805 1.855 7.68 2.025 ;
        RECT 1.805 2.025 3.47 2.105 ;
        RECT 4.045 2.025 7.68 2.105 ;
        RECT 5.28 0.27 6.735 0.45 ;
        RECT 6.565 0.45 6.735 0.655 ;
        RECT 6.565 0.655 7.35 0.825 ;
        RECT 7.17 0.825 7.35 1.34 ;
        RECT 7.17 1.34 7.68 1.855 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.09 1.665 0.385 2.635 ;
      RECT 0.155 0.535 0.355 0.625 ;
      RECT 0.155 0.625 1.24 0.695 ;
      RECT 0.155 0.695 3.835 0.795 ;
      RECT 0.155 0.795 3.13 0.865 ;
      RECT 0.155 0.865 1.795 0.905 ;
      RECT 0.525 0.085 0.855 0.445 ;
      RECT 0.555 1.86 0.775 1.935 ;
      RECT 0.555 1.935 1.635 2.105 ;
      RECT 0.555 2.105 0.775 2.19 ;
      RECT 0.955 2.275 1.285 2.635 ;
      RECT 1.025 0.425 1.24 0.625 ;
      RECT 1.455 2.105 1.635 2.275 ;
      RECT 1.455 2.275 3.435 2.465 ;
      RECT 1.465 0.085 1.635 0.525 ;
      RECT 1.775 0.625 3.835 0.695 ;
      RECT 2.245 0.085 2.575 0.445 ;
      RECT 3.105 0.085 3.435 0.445 ;
      RECT 3.605 0.255 4.92 0.455 ;
      RECT 3.605 0.455 3.835 0.625 ;
      RECT 3.615 2.195 3.885 2.635 ;
      RECT 4.005 0.635 6.17 0.815 ;
      RECT 4.435 2.275 4.765 2.635 ;
      RECT 5.28 2.275 5.61 2.635 ;
      RECT 6.12 2.275 6.455 2.635 ;
      RECT 6.98 0.31 7.68 0.48 ;
      RECT 7.355 2.275 7.685 2.635 ;
      RECT 7.51 0.48 7.68 0.595 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 0.425 1.24 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 0.425 7.68 0.595 ;
    LAYER met1 ;
      RECT 1.01 0.395 1.3 0.44 ;
      RECT 1.01 0.44 7.74 0.58 ;
      RECT 1.01 0.58 1.3 0.625 ;
      RECT 7.45 0.395 7.74 0.44 ;
      RECT 7.45 0.58 7.74 0.625 ;
  END
END sky130_fd_sc_hd__o211ai_4
MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505 1.075 4.455 1.245 ;
        RECT 3.56 1.245 4.455 1.295 ;
        RECT 4.115 0.765 4.455 1.075 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.075 3.335 1.355 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.905 1.365 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.375 1.97 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.022000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.67 0.875 1.54 ;
        RECT 0.545 1.54 3.155 1.71 ;
        RECT 0.545 1.71 0.805 2.465 ;
        RECT 1.475 1.71 1.665 2.465 ;
        RECT 2.825 1.71 3.155 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.095 0.255 2.165 0.445 ;
      RECT 0.115 2.175 0.375 2.635 ;
      RECT 0.975 1.915 1.305 2.635 ;
      RECT 1.045 0.445 2.165 0.465 ;
      RECT 1.045 0.465 1.235 0.89 ;
      RECT 1.405 0.635 3.945 0.845 ;
      RECT 1.835 1.915 2.165 2.635 ;
      RECT 2.395 0.085 2.725 0.445 ;
      RECT 2.395 2.1 2.655 2.295 ;
      RECT 2.395 2.295 3.515 2.465 ;
      RECT 3.255 0.085 3.585 0.445 ;
      RECT 3.325 1.525 4.445 1.695 ;
      RECT 3.325 1.695 3.515 2.295 ;
      RECT 3.685 1.865 4.015 2.635 ;
      RECT 3.755 0.515 3.945 0.635 ;
      RECT 4.115 0.085 4.445 0.445 ;
      RECT 4.185 1.695 4.445 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__o211ai_2
MACRO sky130_fd_sc_hd__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.395 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 0.98 1.325 ;
        RECT 0.605 1.325 0.775 2.25 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 0.995 1.795 1.325 ;
        RECT 1.47 1.325 1.795 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 1.075 2.3 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.418250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.595 1.275 1.815 ;
        RECT 0.945 1.815 2.675 2.045 ;
        RECT 0.945 2.045 1.275 2.445 ;
        RECT 1.965 0.255 2.675 0.845 ;
        RECT 1.975 2.045 2.675 2.465 ;
        RECT 2.47 0.845 2.675 1.815 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 0.255 0.425 0.615 ;
      RECT 0.095 0.615 1.455 0.825 ;
      RECT 0.095 1.575 0.425 2.635 ;
      RECT 0.595 0.085 0.925 0.445 ;
      RECT 1.125 0.255 1.455 0.615 ;
      RECT 1.445 2.275 1.775 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__o211ai_1
MACRO sky130_fd_sc_hd__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 1.075 2.675 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 2.025 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.535 1.345 ;
        RECT 0.085 1.345 0.355 2.445 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.474000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.255 1.285 0.645 ;
        RECT 1.115 0.645 1.355 0.825 ;
        RECT 1.185 0.825 1.355 1.455 ;
        RECT 1.185 1.455 1.795 1.625 ;
        RECT 1.47 1.625 1.795 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.085 0.36 0.825 ;
      RECT 0.525 1.535 1.015 1.705 ;
      RECT 0.525 1.705 0.8 2.21 ;
      RECT 0.58 0.495 0.77 0.655 ;
      RECT 0.58 0.655 0.89 0.825 ;
      RECT 0.72 0.825 0.89 0.995 ;
      RECT 0.72 0.995 1.015 1.535 ;
      RECT 0.97 1.875 1.3 2.635 ;
      RECT 1.49 0.255 1.82 0.485 ;
      RECT 1.57 0.485 1.74 0.735 ;
      RECT 1.57 0.735 2.665 0.905 ;
      RECT 1.995 0.085 2.165 0.555 ;
      RECT 2.27 1.535 2.645 2.635 ;
      RECT 2.335 0.27 2.665 0.735 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__o21bai_1
MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645 1.075 6.81 1.285 ;
        RECT 6.585 1.285 6.81 2.455 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.555 1.285 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.455 4.315 1.625 ;
        RECT 1.065 1.625 1.275 2.465 ;
        RECT 1.42 0.645 2.675 0.815 ;
        RECT 1.865 1.625 2.115 2.465 ;
        RECT 2.445 0.815 2.675 1.075 ;
        RECT 2.445 1.075 2.895 1.445 ;
        RECT 2.445 1.445 4.315 1.455 ;
        RECT 3.225 1.625 3.475 2.125 ;
        RECT 4.065 1.625 4.315 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.145 1.455 0.895 1.625 ;
      RECT 0.145 1.625 0.475 2.435 ;
      RECT 0.225 0.085 0.395 0.895 ;
      RECT 0.565 0.29 0.895 0.895 ;
      RECT 0.645 1.795 0.855 2.635 ;
      RECT 0.725 0.895 0.895 1.075 ;
      RECT 0.725 1.075 2.275 1.285 ;
      RECT 0.725 1.285 0.895 1.455 ;
      RECT 1.08 0.305 3.095 0.475 ;
      RECT 1.445 1.795 1.695 2.635 ;
      RECT 2.285 1.795 2.535 2.635 ;
      RECT 2.775 1.795 3.055 2.295 ;
      RECT 2.775 2.295 4.735 2.465 ;
      RECT 2.845 0.475 3.095 0.725 ;
      RECT 2.845 0.725 6.455 0.905 ;
      RECT 3.265 0.085 3.435 0.555 ;
      RECT 3.605 0.255 3.935 0.725 ;
      RECT 3.645 1.795 3.895 2.295 ;
      RECT 4.105 0.085 4.275 0.555 ;
      RECT 4.445 0.255 4.775 0.725 ;
      RECT 4.485 1.455 6.415 1.625 ;
      RECT 4.485 1.625 4.735 2.295 ;
      RECT 4.905 1.795 5.155 2.635 ;
      RECT 4.945 0.085 5.115 0.555 ;
      RECT 5.285 0.255 5.615 0.725 ;
      RECT 5.325 1.625 5.575 2.465 ;
      RECT 5.745 1.795 5.995 2.635 ;
      RECT 5.785 0.085 5.955 0.555 ;
      RECT 6.125 0.255 6.455 0.725 ;
      RECT 6.165 1.625 6.415 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
  END
END sky130_fd_sc_hd__o21bai_4
MACRO sky130_fd_sc_hd__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.075 4.055 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.075 3.09 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.525 1.325 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.445 2.65 1.615 ;
        RECT 1.085 1.615 1.255 2.465 ;
        RECT 1.525 0.645 1.855 0.905 ;
        RECT 1.525 0.905 1.78 1.445 ;
        RECT 2.405 1.615 2.65 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.18 0.085 0.35 0.825 ;
      RECT 0.18 1.495 0.865 1.665 ;
      RECT 0.18 1.665 0.35 1.915 ;
      RECT 0.585 1.875 0.915 2.635 ;
      RECT 0.6 0.445 0.865 0.825 ;
      RECT 0.695 0.825 0.865 1.075 ;
      RECT 0.695 1.075 1.335 1.245 ;
      RECT 0.695 1.245 0.865 1.495 ;
      RECT 1.075 0.255 2.275 0.475 ;
      RECT 1.075 0.475 1.355 0.905 ;
      RECT 1.47 1.795 1.72 2.635 ;
      RECT 1.955 1.795 2.235 2.295 ;
      RECT 1.955 2.295 3.035 2.465 ;
      RECT 2.025 0.475 2.275 0.725 ;
      RECT 2.025 0.725 3.98 0.905 ;
      RECT 2.445 0.085 2.615 0.555 ;
      RECT 2.785 0.255 3.115 0.725 ;
      RECT 2.865 1.455 3.98 1.665 ;
      RECT 2.865 1.665 3.035 2.295 ;
      RECT 3.205 1.835 3.535 2.635 ;
      RECT 3.285 0.085 3.455 0.555 ;
      RECT 3.625 0.265 3.98 0.725 ;
      RECT 3.705 1.665 3.98 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o21bai_2
MACRO sky130_fd_sc_hd__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 2.35 1.325 ;
        RECT 1.525 1.325 1.77 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585 2.125 2.2 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.86 0.415 3.135 0.76 ;
        RECT 2.86 1.495 3.135 2.465 ;
        RECT 2.965 0.76 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.345 0.905 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 0.515 0.485 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.31 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 1.025 0.255 1.285 0.655 ;
      RECT 1.025 0.655 2.69 0.825 ;
      RECT 1.025 1.495 1.355 1.785 ;
      RECT 1.025 1.785 2.2 1.955 ;
      RECT 1.455 0.085 1.785 0.485 ;
      RECT 1.955 0.305 2.125 0.655 ;
      RECT 2.03 1.495 2.69 1.665 ;
      RECT 2.03 1.665 2.2 1.785 ;
      RECT 2.295 0.085 2.67 0.485 ;
      RECT 2.37 1.835 2.65 2.635 ;
      RECT 2.52 0.825 2.69 0.995 ;
      RECT 2.52 0.995 2.795 1.325 ;
      RECT 2.52 1.325 2.69 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__or3b_1
MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.075 2.23 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 2.125 3.135 2.365 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.64 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.265 1.285 0.595 ;
        RECT 0.935 0.595 1.105 1.495 ;
        RECT 0.935 1.495 1.33 1.7 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.29 0.345 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.81 0.765 1.87 ;
      RECT 0.085 1.87 2.66 1.955 ;
      RECT 0.085 1.955 1.72 2.04 ;
      RECT 0.085 2.04 0.345 2.22 ;
      RECT 0.55 2.21 0.91 2.635 ;
      RECT 0.595 0.085 0.765 0.565 ;
      RECT 0.595 0.905 0.765 1.81 ;
      RECT 1.275 0.765 3.135 0.825 ;
      RECT 1.275 0.825 2.16 0.905 ;
      RECT 1.275 0.905 1.595 0.935 ;
      RECT 1.275 0.935 1.445 1.325 ;
      RECT 1.425 0.735 3.135 0.765 ;
      RECT 1.425 2.21 1.755 2.635 ;
      RECT 1.52 0.085 1.69 0.565 ;
      RECT 1.55 1.785 2.66 1.87 ;
      RECT 1.99 0.305 2.16 0.655 ;
      RECT 1.99 0.655 3.135 0.735 ;
      RECT 2.33 0.085 2.66 0.485 ;
      RECT 2.49 0.995 2.79 1.325 ;
      RECT 2.49 1.325 2.66 1.785 ;
      RECT 2.83 0.305 3.085 0.605 ;
      RECT 2.83 0.605 3.135 0.655 ;
      RECT 2.83 1.495 3.135 1.925 ;
      RECT 2.965 0.825 3.135 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__or3b_2
MACRO sky130_fd_sc_hd__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 1.415 2.72 1.7 ;
        RECT 2.535 0.995 2.72 1.415 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.89 0.995 3.2 1.7 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.64 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.735 2.025 0.905 ;
        RECT 0.935 0.905 1.105 1.415 ;
        RECT 0.935 1.415 2.22 1.7 ;
        RECT 1 0.285 1.33 0.735 ;
        RECT 1.855 0.255 2.09 0.585 ;
        RECT 1.855 0.585 2.025 0.735 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.29 0.345 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.81 0.765 1.87 ;
      RECT 0.085 1.87 3.62 2.04 ;
      RECT 0.085 2.04 0.345 2.22 ;
      RECT 0.55 2.21 0.91 2.635 ;
      RECT 0.595 0.905 0.765 1.81 ;
      RECT 0.62 0.085 0.79 0.565 ;
      RECT 1.275 1.075 2.365 1.245 ;
      RECT 1.42 2.21 1.75 2.635 ;
      RECT 1.5 0.085 1.67 0.565 ;
      RECT 2.195 0.72 4.055 0.825 ;
      RECT 2.195 0.825 2.4 0.89 ;
      RECT 2.195 0.89 2.365 1.075 ;
      RECT 2.25 0.655 4.055 0.72 ;
      RECT 2.255 2.21 2.595 2.635 ;
      RECT 2.26 0.085 2.59 0.485 ;
      RECT 2.76 0.305 2.93 0.655 ;
      RECT 3.1 0.085 3.49 0.485 ;
      RECT 3.39 0.995 3.68 1.325 ;
      RECT 3.39 1.325 3.62 1.87 ;
      RECT 3.52 2.21 4.055 2.425 ;
      RECT 3.66 0.305 3.915 0.605 ;
      RECT 3.66 0.605 4.055 0.655 ;
      RECT 3.85 0.825 4.055 2.21 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__or3b_4
MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.495 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.075 3.08 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.845 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 3.925 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.355 1.665 2.685 2.465 ;
        RECT 3.37 1.055 3.925 1.445 ;
        RECT 3.595 0.635 3.925 1.055 ;
        RECT 3.595 1.665 3.925 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 1.185 0.905 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.935 0.255 2.125 0.465 ;
      RECT 0.935 0.465 1.185 0.735 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.355 0.635 3.085 0.905 ;
      RECT 1.855 1.835 2.185 2.635 ;
      RECT 2.315 0.255 4.425 0.465 ;
      RECT 2.995 1.835 3.325 2.635 ;
      RECT 3.255 0.465 3.425 0.885 ;
      RECT 4.095 0.465 4.425 0.905 ;
      RECT 4.095 1.445 4.425 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__nand4_2
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.995 2.215 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 0.3 1.35 0.825 ;
        RECT 1.145 0.825 1.35 0.995 ;
        RECT 1.145 0.995 1.455 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.3 0.81 0.995 ;
        RECT 0.595 0.995 0.975 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 0.995 0.395 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.795000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 1.795 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.385 1.665 1.715 2.465 ;
        RECT 1.52 0.255 2.215 0.825 ;
        RECT 1.625 0.825 1.795 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 0.09 0.085 0.425 0.825 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.915 1.835 2.195 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nand4_1
MACRO sky130_fd_sc_hd__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.71 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.85 1.075 5.565 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.54 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.7 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 7.305 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 6.11 0.655 7.305 0.905 ;
        RECT 6.11 0.905 6.29 1.445 ;
        RECT 6.135 1.665 6.465 2.465 ;
        RECT 6.975 1.665 7.305 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.09 0.255 0.345 0.655 ;
      RECT 0.09 0.655 2.025 0.905 ;
      RECT 0.09 1.445 0.345 2.635 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 1.015 0.255 1.185 0.655 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.355 0.085 1.685 0.485 ;
      RECT 1.855 0.255 3.785 0.485 ;
      RECT 1.855 0.485 2.025 0.655 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.195 0.655 5.565 0.905 ;
      RECT 2.695 1.835 2.865 2.635 ;
      RECT 3.535 1.835 4.225 2.635 ;
      RECT 3.975 0.255 7.73 0.485 ;
      RECT 4.895 1.835 5.065 2.635 ;
      RECT 5.77 0.485 5.94 0.905 ;
      RECT 5.77 1.835 5.94 2.635 ;
      RECT 6.635 1.835 6.805 2.635 ;
      RECT 7.475 0.485 7.73 0.905 ;
      RECT 7.475 1.445 7.735 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__nand4_4
MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 1.005 2.16 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615 0.255 11.875 0.825 ;
        RECT 11.615 1.445 11.875 2.465 ;
        RECT 11.66 0.825 11.875 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.2 0.255 10.485 0.715 ;
        RECT 10.2 1.63 10.485 2.465 ;
        RECT 10.28 0.715 10.485 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315 1.095 9.69 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.59 0.735 4 0.965 ;
        RECT 3.59 0.965 3.92 1.065 ;
      LAYER mcon ;
        RECT 3.83 0.765 4 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.46 0.735 7.835 1.065 ;
      LAYER mcon ;
        RECT 7.51 0.765 7.68 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.77 0.735 4.06 0.78 ;
        RECT 3.77 0.78 7.74 0.92 ;
        RECT 3.77 0.92 4.06 0.965 ;
        RECT 7.45 0.735 7.74 0.78 ;
        RECT 7.45 0.92 7.74 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.15 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.84 0.805 ;
      RECT 0.085 1.795 0.84 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.41 0.635 2.125 0.825 ;
      RECT 1.41 0.825 1.58 1.795 ;
      RECT 1.41 1.795 2.125 1.965 ;
      RECT 1.435 0.085 1.785 0.465 ;
      RECT 1.435 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.33 0.705 2.55 1.575 ;
      RECT 2.33 1.575 2.83 1.955 ;
      RECT 2.34 2.25 3.17 2.42 ;
      RECT 2.405 0.265 3.4 0.465 ;
      RECT 2.73 0.645 3.06 1.015 ;
      RECT 3 1.195 3.4 1.235 ;
      RECT 3 1.235 4.35 1.405 ;
      RECT 3 1.405 3.17 2.25 ;
      RECT 3.23 0.465 3.4 1.195 ;
      RECT 3.34 1.575 3.59 1.785 ;
      RECT 3.34 1.785 4.69 2.035 ;
      RECT 3.41 2.205 3.79 2.635 ;
      RECT 3.57 0.085 3.74 0.525 ;
      RECT 3.91 0.255 5.08 0.425 ;
      RECT 3.91 0.425 4.24 0.545 ;
      RECT 4.09 2.035 4.26 2.375 ;
      RECT 4.1 1.405 4.35 1.485 ;
      RECT 4.13 1.155 4.35 1.235 ;
      RECT 4.41 0.595 4.74 0.765 ;
      RECT 4.52 0.765 4.74 0.895 ;
      RECT 4.52 0.895 5.83 1.065 ;
      RECT 4.52 1.065 4.69 1.785 ;
      RECT 4.86 1.235 5.19 1.415 ;
      RECT 4.86 1.415 5.865 1.655 ;
      RECT 4.88 1.915 5.21 2.635 ;
      RECT 4.91 0.425 5.08 0.715 ;
      RECT 5.35 0.085 5.68 0.465 ;
      RECT 5.5 1.065 5.83 1.235 ;
      RECT 6.065 1.575 6.3 1.985 ;
      RECT 6.125 0.705 6.41 1.125 ;
      RECT 6.125 1.125 6.745 1.305 ;
      RECT 6.255 2.25 7.085 2.42 ;
      RECT 6.32 0.265 7.085 0.465 ;
      RECT 6.54 1.305 6.745 1.905 ;
      RECT 6.915 0.465 7.085 1.235 ;
      RECT 6.915 1.235 8.265 1.405 ;
      RECT 6.915 1.405 7.085 2.25 ;
      RECT 7.255 1.575 7.505 1.915 ;
      RECT 7.255 1.915 10.03 2.085 ;
      RECT 7.265 0.085 7.525 0.525 ;
      RECT 7.325 2.255 7.705 2.635 ;
      RECT 7.785 0.255 8.955 0.425 ;
      RECT 7.785 0.425 8.115 0.545 ;
      RECT 7.945 2.085 8.115 2.375 ;
      RECT 8.045 1.075 8.265 1.235 ;
      RECT 8.285 0.595 8.615 0.78 ;
      RECT 8.435 0.78 8.615 1.915 ;
      RECT 8.645 2.255 10.03 2.635 ;
      RECT 8.785 0.425 8.955 0.585 ;
      RECT 8.785 0.755 9.475 0.925 ;
      RECT 8.785 0.925 9.06 1.575 ;
      RECT 8.785 1.575 9.545 1.745 ;
      RECT 9.24 0.265 9.475 0.755 ;
      RECT 9.7 0.085 10.03 0.805 ;
      RECT 9.86 0.995 10.11 1.325 ;
      RECT 9.86 1.325 10.03 1.915 ;
      RECT 10.655 0.255 10.97 0.995 ;
      RECT 10.655 0.995 11.49 1.325 ;
      RECT 10.655 1.325 10.97 2.415 ;
      RECT 11.15 0.085 11.445 0.545 ;
      RECT 11.15 1.765 11.445 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.45 1.785 2.62 1.955 ;
      RECT 2.89 0.765 3.06 0.935 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.67 1.445 5.84 1.615 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.13 1.105 6.3 1.275 ;
      RECT 6.13 1.785 6.3 1.955 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.89 1.445 9.06 1.615 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 6.36 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 3.12 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.39 1.755 2.68 1.8 ;
      RECT 2.39 1.94 2.68 1.985 ;
      RECT 2.83 0.735 3.12 0.78 ;
      RECT 2.83 0.92 3.12 0.965 ;
      RECT 2.925 0.965 3.12 1.12 ;
      RECT 2.925 1.12 6.36 1.26 ;
      RECT 5.61 1.415 5.9 1.46 ;
      RECT 5.61 1.46 9.12 1.6 ;
      RECT 5.61 1.6 5.9 1.645 ;
      RECT 6.07 1.075 6.36 1.12 ;
      RECT 6.07 1.26 6.36 1.305 ;
      RECT 6.07 1.755 6.36 1.8 ;
      RECT 6.07 1.94 6.36 1.985 ;
      RECT 8.83 1.415 9.12 1.46 ;
      RECT 8.83 1.6 9.12 1.645 ;
  END
END sky130_fd_sc_hd__dfbbp_1
MACRO sky130_fd_sc_hd__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.285 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.28 0.825 0.995 ;
        RECT 0.605 0.995 1 1.325 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.03 1.075 2.615 1.325 ;
        RECT 2.445 1.325 2.615 2.425 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.56 0.43 1.81 0.79 ;
        RECT 1.64 0.79 1.81 1.495 ;
        RECT 1.64 1.495 2.27 1.665 ;
        RECT 1.94 1.665 2.27 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 0.085 0.425 0.815 ;
      RECT 0.15 1.455 0.4 2.635 ;
      RECT 0.57 1.495 1.34 1.665 ;
      RECT 0.57 1.665 0.82 2.465 ;
      RECT 0.99 1.835 1.77 2.635 ;
      RECT 1 0.28 1.34 0.825 ;
      RECT 1.17 0.825 1.34 0.995 ;
      RECT 1.17 0.995 1.47 1.325 ;
      RECT 1.17 1.325 1.34 1.495 ;
      RECT 1.98 0.425 2.27 0.725 ;
      RECT 1.98 0.725 3.11 0.905 ;
      RECT 2.44 0.085 2.61 0.555 ;
      RECT 2.78 0.275 3.11 0.725 ;
      RECT 2.82 1.455 3.07 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o2bb2ai_1
MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 3.505 1.285 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 1.825 1.285 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.045 1.075 10.005 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.875 1.285 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415 0.645 6.155 0.905 ;
        RECT 4.425 1.455 7.715 1.625 ;
        RECT 4.425 1.625 4.675 2.465 ;
        RECT 5.265 1.625 5.515 2.465 ;
        RECT 5.875 0.905 6.155 1.455 ;
        RECT 6.625 1.625 6.875 2.125 ;
        RECT 7.465 1.625 7.715 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135 -0.085 0.305 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.085 0.645 1.705 0.905 ;
      RECT 0.085 0.905 0.255 1.455 ;
      RECT 0.085 1.455 3.915 1.625 ;
      RECT 0.1 0.255 2.125 0.475 ;
      RECT 0.155 1.795 0.405 2.635 ;
      RECT 0.575 1.625 0.825 2.465 ;
      RECT 0.995 1.795 1.245 2.635 ;
      RECT 1.415 1.625 1.665 2.465 ;
      RECT 1.835 1.795 2.085 2.635 ;
      RECT 1.875 0.475 2.125 0.725 ;
      RECT 1.875 0.725 3.805 0.905 ;
      RECT 2.255 1.625 2.505 2.465 ;
      RECT 2.295 0.085 2.465 0.555 ;
      RECT 2.635 0.255 2.965 0.725 ;
      RECT 2.675 1.795 2.925 2.635 ;
      RECT 3.095 1.625 3.345 2.465 ;
      RECT 3.135 0.085 3.305 0.555 ;
      RECT 3.475 0.255 3.805 0.725 ;
      RECT 3.515 1.795 4.255 2.635 ;
      RECT 3.745 1.075 5.705 1.285 ;
      RECT 3.745 1.285 3.915 1.455 ;
      RECT 4.06 0.255 6.495 0.475 ;
      RECT 4.06 0.475 4.245 0.835 ;
      RECT 4.845 1.795 5.095 2.635 ;
      RECT 5.685 1.795 5.935 2.635 ;
      RECT 6.175 1.795 6.455 2.295 ;
      RECT 6.175 2.295 8.135 2.465 ;
      RECT 6.325 0.475 6.495 0.735 ;
      RECT 6.325 0.735 9.855 0.905 ;
      RECT 6.665 0.085 6.835 0.555 ;
      RECT 7.005 0.255 7.335 0.725 ;
      RECT 7.005 0.725 9.855 0.735 ;
      RECT 7.045 1.795 7.295 2.295 ;
      RECT 7.505 0.085 7.675 0.555 ;
      RECT 7.845 0.255 8.175 0.725 ;
      RECT 7.885 1.455 9.875 1.625 ;
      RECT 7.885 1.625 8.135 2.295 ;
      RECT 8.305 1.795 8.555 2.635 ;
      RECT 8.345 0.085 8.515 0.555 ;
      RECT 8.685 0.255 9.015 0.725 ;
      RECT 8.725 1.625 8.975 2.465 ;
      RECT 9.145 1.795 9.395 2.635 ;
      RECT 9.185 0.085 9.355 0.555 ;
      RECT 9.525 0.255 9.855 0.725 ;
      RECT 9.565 1.625 9.875 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4
MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.625 1.445 ;
        RECT 0.09 1.445 1.945 1.615 ;
        RECT 1.615 1.075 1.945 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795 1.075 1.4 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.41 1.075 3.74 1.445 ;
        RECT 3.41 1.445 5.435 1.615 ;
        RECT 4.73 1.075 5.435 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.96 1.075 4.5 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745 0.645 3.075 1.075 ;
        RECT 2.745 1.075 3.215 1.785 ;
        RECT 2.745 1.785 4.33 1.955 ;
        RECT 2.745 1.955 3.035 2.465 ;
        RECT 4.08 1.955 4.33 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.15 1.795 0.4 2.635 ;
      RECT 0.195 0.085 0.365 0.895 ;
      RECT 0.535 0.305 1.705 0.475 ;
      RECT 0.535 0.475 0.785 0.895 ;
      RECT 0.575 1.785 2.285 1.965 ;
      RECT 0.575 1.965 0.825 2.465 ;
      RECT 0.955 0.645 1.285 0.725 ;
      RECT 0.955 0.725 2.285 0.905 ;
      RECT 0.995 2.135 1.245 2.635 ;
      RECT 1.415 1.965 1.665 2.125 ;
      RECT 1.835 2.135 2.575 2.635 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.115 0.905 2.285 0.995 ;
      RECT 2.115 0.995 2.575 1.325 ;
      RECT 2.115 1.325 2.285 1.785 ;
      RECT 2.325 0.255 3.53 0.475 ;
      RECT 2.325 0.475 2.575 0.555 ;
      RECT 3.205 2.125 3.49 2.635 ;
      RECT 3.245 0.475 3.53 0.735 ;
      RECT 3.245 0.735 5.21 0.905 ;
      RECT 3.66 2.125 3.91 2.295 ;
      RECT 3.66 2.295 4.75 2.465 ;
      RECT 3.7 0.085 3.87 0.555 ;
      RECT 4.04 0.255 4.37 0.725 ;
      RECT 4.04 0.725 5.21 0.735 ;
      RECT 4.5 1.785 4.75 2.295 ;
      RECT 4.54 0.085 4.71 0.555 ;
      RECT 4.88 0.255 5.21 0.725 ;
      RECT 4.965 1.795 5.17 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2
MACRO sky130_fd_sc_hd__a41oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 0.995 3.085 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 0.755 2.21 1.665 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 0.755 1.71 1.665 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 0.965 1.25 1.665 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.965 0.78 1.665 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.669500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.285 0.345 0.615 ;
        RECT 0.09 0.615 1.29 0.785 ;
        RECT 0.09 0.785 0.36 1.845 ;
        RECT 0.09 1.845 0.425 2.425 ;
        RECT 1.12 0.295 3.015 0.465 ;
        RECT 1.12 0.465 1.29 0.615 ;
        RECT 2.685 0.465 3.015 0.805 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.595 1.845 3.015 2.015 ;
      RECT 0.595 2.015 0.845 2.465 ;
      RECT 0.62 0.085 0.95 0.445 ;
      RECT 1.12 2.195 1.45 2.635 ;
      RECT 1.76 2.015 1.93 2.465 ;
      RECT 2.215 2.195 2.545 2.635 ;
      RECT 2.765 2.015 3.015 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a41oi_1
MACRO sky130_fd_sc_hd__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785 1.075 2.455 1.295 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665 1.075 3.365 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.075 4.575 1.295 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.755 1.075 5.895 1.295 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.555 1.28 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.645 2.295 0.815 ;
        RECT 0.145 0.815 0.315 1.455 ;
        RECT 0.145 1.455 1.455 1.625 ;
        RECT 0.685 0.255 0.855 0.645 ;
        RECT 1.125 1.625 1.455 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.185 0.085 0.515 0.465 ;
      RECT 0.785 1.795 0.955 2.295 ;
      RECT 0.785 2.295 1.795 2.465 ;
      RECT 1.025 0.085 1.375 0.465 ;
      RECT 1.545 0.295 2.635 0.465 ;
      RECT 1.625 1.535 5.76 1.705 ;
      RECT 1.625 1.705 1.795 2.295 ;
      RECT 1.965 1.915 2.295 2.635 ;
      RECT 2.465 0.465 2.635 0.645 ;
      RECT 2.465 0.645 3.555 0.815 ;
      RECT 2.465 1.705 2.635 2.465 ;
      RECT 2.805 0.295 4.495 0.465 ;
      RECT 2.805 1.915 3.135 2.635 ;
      RECT 3.325 1.705 3.495 2.465 ;
      RECT 3.745 0.645 5.675 0.815 ;
      RECT 3.755 1.915 4.425 2.635 ;
      RECT 4.665 1.705 4.835 2.465 ;
      RECT 5.005 0.085 5.335 0.465 ;
      RECT 5.005 1.915 5.335 2.635 ;
      RECT 5.505 0.255 5.675 0.645 ;
      RECT 5.505 1.705 5.675 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__a41oi_2
MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.995 4.205 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405 1.075 6.315 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.56 1.075 7.955 1.3 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.075 9.975 1.28 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.745 1.305 ;
        RECT 0.105 1.305 0.325 1.965 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.575 2.155 1.685 ;
        RECT 0.515 1.685 1.685 1.745 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 0.635 4.015 0.805 ;
        RECT 1.35 1.495 2.155 1.575 ;
        RECT 1.35 1.745 1.685 2.085 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.935 0.805 2.155 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.09 0.085 0.425 0.465 ;
      RECT 0.09 2.255 2.335 2.425 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 1.775 0.085 2.105 0.465 ;
      RECT 2.165 1.905 3.515 2.075 ;
      RECT 2.165 2.075 2.335 2.255 ;
      RECT 2.165 2.425 2.335 2.465 ;
      RECT 2.425 0.295 6.115 0.465 ;
      RECT 2.505 2.255 3.175 2.635 ;
      RECT 3.345 1.575 9.945 1.745 ;
      RECT 3.345 1.745 3.515 1.905 ;
      RECT 3.345 2.075 3.515 2.465 ;
      RECT 3.685 1.915 4.015 2.635 ;
      RECT 4.185 1.745 4.355 2.425 ;
      RECT 4.525 0.635 7.895 0.805 ;
      RECT 4.62 1.915 4.95 2.635 ;
      RECT 5.12 1.745 5.29 2.465 ;
      RECT 5.495 1.915 6.165 2.635 ;
      RECT 6.305 0.295 8.235 0.465 ;
      RECT 6.385 1.745 6.555 2.465 ;
      RECT 6.725 1.915 7.055 2.635 ;
      RECT 7.225 1.745 7.395 2.465 ;
      RECT 7.565 1.915 7.895 2.635 ;
      RECT 8.065 0.255 8.235 0.295 ;
      RECT 8.065 0.465 8.235 0.635 ;
      RECT 8.065 0.635 9.915 0.805 ;
      RECT 8.065 1.745 8.235 2.465 ;
      RECT 8.405 0.085 8.735 0.465 ;
      RECT 8.405 1.915 8.735 2.635 ;
      RECT 8.905 0.255 9.075 0.635 ;
      RECT 8.905 1.745 9.075 2.465 ;
      RECT 9.245 0.085 9.575 0.465 ;
      RECT 9.245 1.915 9.575 2.635 ;
      RECT 9.745 0.255 9.915 0.635 ;
      RECT 9.775 1.745 9.945 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__a41oi_4
MACRO sky130_fd_sc_hd__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345 1.075 2.675 1.275 ;
        RECT 2.445 1.275 2.675 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705 1.075 2.035 1.095 ;
        RECT 1.705 1.095 2.155 1.275 ;
        RECT 1.94 1.275 2.155 2.39 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.535 1.305 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 1.03 ;
        RECT 0.085 1.03 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.535 1.86 1.245 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.595 0.715 1.305 0.905 ;
      RECT 0.595 0.905 0.88 1.475 ;
      RECT 0.595 1.475 1.745 1.69 ;
      RECT 1.005 0.255 1.365 0.52 ;
      RECT 1.005 0.52 1.36 0.525 ;
      RECT 1.005 0.525 1.355 0.535 ;
      RECT 1.005 0.535 1.35 0.54 ;
      RECT 1.005 0.54 1.345 0.55 ;
      RECT 1.005 0.55 1.34 0.555 ;
      RECT 1.005 0.555 1.33 0.565 ;
      RECT 1.005 0.565 1.32 0.575 ;
      RECT 1.005 0.575 1.305 0.715 ;
      RECT 1.415 1.69 1.745 2.465 ;
      RECT 1.495 0.635 1.825 0.715 ;
      RECT 1.495 0.715 2.675 0.905 ;
      RECT 1.995 0.085 2.165 0.545 ;
      RECT 2.335 0.255 2.675 0.715 ;
      RECT 2.335 1.915 2.665 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__o21a_1
MACRO sky130_fd_sc_hd__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.48 0.99 3.785 1.495 ;
        RECT 3.48 1.495 5.4 1.705 ;
        RECT 5.03 0.995 5.4 1.495 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.14 0.995 4.69 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.075 3.155 1.615 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.635 1.715 0.805 ;
        RECT 0.09 0.805 0.32 1.53 ;
        RECT 0.09 1.53 1.955 1.7 ;
        RECT 0.595 0.615 1.715 0.635 ;
        RECT 0.915 1.7 1.105 2.465 ;
        RECT 1.775 1.7 1.955 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 0.415 1.87 0.745 2.635 ;
      RECT 0.49 0.995 2.315 1.335 ;
      RECT 0.955 0.085 1.285 0.445 ;
      RECT 1.275 1.87 1.605 2.635 ;
      RECT 1.815 0.085 2.145 0.465 ;
      RECT 2.115 0.655 3.095 0.87 ;
      RECT 2.115 0.87 2.315 0.995 ;
      RECT 2.125 1.335 2.315 1.83 ;
      RECT 2.125 1.83 2.845 1.875 ;
      RECT 2.125 1.875 4.545 2.085 ;
      RECT 2.135 2.255 2.485 2.635 ;
      RECT 2.335 0.255 3.605 0.485 ;
      RECT 2.655 2.085 4.545 2.105 ;
      RECT 2.655 2.105 2.845 2.465 ;
      RECT 3.015 2.275 3.685 2.635 ;
      RECT 3.275 0.485 3.605 0.615 ;
      RECT 3.275 0.615 5.405 0.785 ;
      RECT 3.775 0.085 4.115 0.445 ;
      RECT 4.215 2.105 4.545 2.445 ;
      RECT 4.645 0.085 4.975 0.445 ;
      RECT 5.075 1.935 5.435 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__o21a_4
MACRO sky130_fd_sc_hd__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.125 1.45 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.025 2.61 1.4 ;
        RECT 2.405 1.4 2.61 1.985 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 1.01 1.855 1.615 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.53 0.255 0.775 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 1.635 0.345 2.635 ;
      RECT 0.105 0.085 0.345 0.885 ;
      RECT 0.945 0.085 1.275 0.465 ;
      RECT 0.945 0.635 1.795 0.84 ;
      RECT 0.945 0.84 1.275 1.33 ;
      RECT 0.945 2.185 1.795 2.635 ;
      RECT 1.105 1.33 1.275 1.785 ;
      RECT 1.105 1.785 2.225 2.005 ;
      RECT 1.465 0.255 1.795 0.635 ;
      RECT 1.965 0.465 2.175 0.635 ;
      RECT 1.965 0.635 3.12 0.825 ;
      RECT 1.965 2.005 2.225 2.465 ;
      RECT 2.345 0.085 2.675 0.465 ;
      RECT 2.795 1.65 3.12 2.635 ;
      RECT 2.845 0.495 3.12 0.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o21a_2
MACRO sky130_fd_sc_hd__clkdlybuf4s15_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.56 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.285 3.595 0.545 ;
        RECT 3.21 1.76 3.595 2.465 ;
        RECT 3.365 0.545 3.595 1.76 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.215 0.885 ;
      RECT 0.085 1.495 1.215 1.665 ;
      RECT 0.085 1.665 0.425 2.465 ;
      RECT 0.595 0.085 0.91 0.545 ;
      RECT 0.595 1.835 0.925 2.635 ;
      RECT 0.73 0.885 1.215 1.495 ;
      RECT 1.385 0.255 1.76 0.825 ;
      RECT 1.385 1.835 1.76 2.465 ;
      RECT 1.59 0.825 1.76 1.055 ;
      RECT 1.59 1.055 2.685 1.25 ;
      RECT 1.59 1.25 1.76 1.835 ;
      RECT 1.93 0.255 2.26 0.715 ;
      RECT 1.93 0.715 3.195 0.885 ;
      RECT 1.93 1.42 3.195 1.59 ;
      RECT 1.93 1.59 2.41 2.465 ;
      RECT 2.64 1.76 3.04 2.635 ;
      RECT 2.71 0.085 3.04 0.545 ;
      RECT 2.855 0.885 3.195 1.42 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_1
MACRO sky130_fd_sc_hd__clkdlybuf4s15_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.06 0.555 1.625 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 0.255 3.55 0.64 ;
        RECT 3.07 1.485 3.55 2.465 ;
        RECT 3.355 0.64 3.55 1.485 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.255 0.415 0.72 ;
      RECT 0.085 0.72 1.06 0.89 ;
      RECT 0.085 1.795 1.06 1.965 ;
      RECT 0.085 1.965 0.43 2.465 ;
      RECT 0.585 0.085 0.915 0.55 ;
      RECT 0.6 2.135 0.93 2.635 ;
      RECT 0.89 0.89 1.06 1.075 ;
      RECT 0.89 1.075 1.32 1.245 ;
      RECT 0.89 1.245 1.06 1.795 ;
      RECT 1.23 1.785 1.66 2.465 ;
      RECT 1.28 0.255 1.66 0.905 ;
      RECT 1.49 0.905 1.66 1.075 ;
      RECT 1.49 1.075 2.415 1.485 ;
      RECT 1.49 1.485 1.66 1.785 ;
      RECT 1.83 0.255 2.1 0.735 ;
      RECT 1.83 0.735 2.9 0.905 ;
      RECT 1.83 1.79 2.9 1.965 ;
      RECT 1.83 1.965 2.1 2.465 ;
      RECT 2.55 0.085 2.88 0.565 ;
      RECT 2.55 2.135 2.88 2.635 ;
      RECT 2.73 0.905 2.9 1.075 ;
      RECT 2.73 1.075 3.185 1.245 ;
      RECT 2.73 1.245 2.9 1.79 ;
      RECT 3.72 0.085 4.055 0.645 ;
      RECT 3.72 1.485 4.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_2
MACRO sky130_fd_sc_hd__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.075 3.005 1.245 ;
        RECT 1.66 1.035 3.005 1.075 ;
        RECT 1.66 1.245 3.005 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.035 1.385 1.445 ;
        RECT 0.1 1.445 3.575 1.625 ;
        RECT 3.245 1.035 3.575 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.745 1.035 4.755 1.275 ;
        RECT 3.745 1.275 4.46 1.615 ;
      LAYER mcon ;
        RECT 3.83 1.445 4 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.59 0.995 6.935 1.325 ;
        RECT 6.59 1.325 6.76 1.615 ;
      LAYER mcon ;
        RECT 6.59 1.445 6.76 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.77 1.415 4.06 1.46 ;
        RECT 3.77 1.46 6.82 1.6 ;
        RECT 3.77 1.6 4.06 1.645 ;
        RECT 6.53 1.415 6.82 1.46 ;
        RECT 6.53 1.6 6.82 1.645 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5 1.035 6.35 1.275 ;
        RECT 6.13 1.275 6.35 1.695 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 0.675 3.33 0.695 ;
        RECT 1.775 0.695 7.275 0.825 ;
        RECT 1.775 0.825 6.355 0.865 ;
        RECT 3.875 0.255 4.195 0.615 ;
        RECT 3.875 0.615 5.045 0.625 ;
        RECT 3.875 0.625 7.275 0.695 ;
        RECT 4.875 0.255 5.045 0.615 ;
        RECT 5.17 1.865 7.275 2.085 ;
        RECT 5.715 0.255 5.885 0.615 ;
        RECT 5.715 0.615 7.275 0.625 ;
        RECT 6.93 1.495 7.275 1.865 ;
        RECT 7.105 0.825 7.275 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.095 0.085 0.395 0.585 ;
      RECT 0.095 1.795 3.705 2.085 ;
      RECT 0.095 2.085 0.345 2.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 0.565 0.53 0.775 0.695 ;
      RECT 0.565 0.695 1.605 0.865 ;
      RECT 0.95 0.085 1.185 0.525 ;
      RECT 1.015 2.085 3.705 2.105 ;
      RECT 1.015 2.105 1.185 2.465 ;
      RECT 1.355 0.255 3.365 0.505 ;
      RECT 1.355 0.505 1.605 0.695 ;
      RECT 1.355 2.275 1.685 2.635 ;
      RECT 1.855 2.105 2.025 2.465 ;
      RECT 2.195 2.275 2.525 2.635 ;
      RECT 2.695 2.105 2.865 2.465 ;
      RECT 3.035 2.275 3.365 2.635 ;
      RECT 3.535 0.085 3.705 0.525 ;
      RECT 3.535 2.105 3.705 2.255 ;
      RECT 3.535 2.255 7.27 2.465 ;
      RECT 3.875 1.785 4.91 2.085 ;
      RECT 4.365 0.085 4.695 0.445 ;
      RECT 4.63 1.445 5.96 1.695 ;
      RECT 4.63 1.695 4.91 1.785 ;
      RECT 5.215 0.085 5.545 0.445 ;
      RECT 6.055 0.085 6.385 0.445 ;
      RECT 6.915 0.085 7.27 0.445 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__a211oi_4
MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.37 1.035 3.08 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.74 1.035 4.5 1.285 ;
        RECT 4.175 1.285 4.5 1.655 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.035 1.785 1.285 ;
        RECT 1.035 1.285 1.255 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.995 0.405 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.826000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 0.255 0.835 0.655 ;
        RECT 0.575 0.655 3.145 0.855 ;
        RECT 0.575 0.855 0.855 1.785 ;
        RECT 0.575 1.785 0.905 2.105 ;
        RECT 1.505 0.285 1.695 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.145 0.085 0.395 0.815 ;
      RECT 0.145 1.785 0.405 2.285 ;
      RECT 0.145 2.285 2.215 2.455 ;
      RECT 1.005 0.085 1.335 0.475 ;
      RECT 1.075 1.785 1.265 2.255 ;
      RECT 1.075 2.255 2.215 2.285 ;
      RECT 1.435 1.455 3.975 1.655 ;
      RECT 1.435 1.655 1.765 2.075 ;
      RECT 1.865 0.085 2.195 0.475 ;
      RECT 1.935 1.835 2.215 2.255 ;
      RECT 2.385 0.265 3.495 0.475 ;
      RECT 2.435 1.835 2.665 2.635 ;
      RECT 2.845 1.655 3.115 2.465 ;
      RECT 3.295 1.835 3.525 2.635 ;
      RECT 3.325 0.475 3.495 0.635 ;
      RECT 3.325 0.635 4.435 0.855 ;
      RECT 3.675 0.085 4.005 0.455 ;
      RECT 3.705 1.655 3.975 2.465 ;
      RECT 4.155 1.835 4.385 2.635 ;
      RECT 4.185 0.265 4.435 0.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__a211oi_2
MACRO sky130_fd_sc_hd__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.265 0.855 0.995 ;
        RECT 0.605 0.995 1.245 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.765 0.435 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425 0.995 1.755 1.325 ;
        RECT 1.525 1.325 1.755 2.455 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 2.235 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.619250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.18 0.265 1.365 0.625 ;
        RECT 1.18 0.625 2.66 0.815 ;
        RECT 1.935 1.785 2.66 2.455 ;
        RECT 2.055 0.265 2.28 0.625 ;
        RECT 2.445 0.815 2.66 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.085 0.425 0.595 ;
      RECT 0.25 1.525 1.355 1.725 ;
      RECT 0.25 1.725 0.5 2.455 ;
      RECT 0.67 1.905 1 2.635 ;
      RECT 1.17 1.725 1.355 2.455 ;
      RECT 1.545 0.085 1.875 0.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__a211oi_1
MACRO sky130_fd_sc_hd__a2111o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.495 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675 1.075 5.625 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.975 3.255 1.285 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.975 2.28 1.285 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.37 1.625 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.165 0.255 6.355 0.635 ;
        RECT 6.165 0.635 7.735 0.805 ;
        RECT 6.165 1.465 7.735 1.635 ;
        RECT 6.165 1.635 7.215 1.715 ;
        RECT 6.165 1.715 6.355 2.465 ;
        RECT 7.025 0.255 7.215 0.635 ;
        RECT 7.025 1.715 7.215 2.465 ;
        RECT 7.49 0.805 7.735 1.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.11 1.795 0.37 2.295 ;
      RECT 0.11 2.295 2.16 2.465 ;
      RECT 0.18 0.255 0.44 0.635 ;
      RECT 0.18 0.635 3.655 0.805 ;
      RECT 0.54 0.805 0.87 2.125 ;
      RECT 0.61 0.085 0.94 0.465 ;
      RECT 1.04 1.455 1.23 2.295 ;
      RECT 1.11 0.255 1.34 0.615 ;
      RECT 1.11 0.615 3.655 0.635 ;
      RECT 1.4 1.455 3.1 1.625 ;
      RECT 1.4 1.625 1.73 2.125 ;
      RECT 1.51 0.085 1.84 0.445 ;
      RECT 1.9 1.795 2.16 2.295 ;
      RECT 2.015 0.255 2.24 0.615 ;
      RECT 2.34 1.795 2.675 2.295 ;
      RECT 2.34 2.295 3.65 2.465 ;
      RECT 2.42 0.085 3.295 0.445 ;
      RECT 2.845 1.625 3.1 2.125 ;
      RECT 3.32 1.795 5.495 1.995 ;
      RECT 3.32 1.995 3.65 2.295 ;
      RECT 3.465 0.255 4.585 0.445 ;
      RECT 3.465 0.445 3.655 0.615 ;
      RECT 3.465 0.805 3.655 1.445 ;
      RECT 3.465 1.445 5.975 1.625 ;
      RECT 3.825 0.615 5.495 0.785 ;
      RECT 3.865 2.165 4.195 2.635 ;
      RECT 4.365 1.995 4.625 2.415 ;
      RECT 4.805 0.085 5.14 0.445 ;
      RECT 4.805 2.255 5.14 2.635 ;
      RECT 5.31 0.255 5.495 0.615 ;
      RECT 5.31 1.995 5.495 2.465 ;
      RECT 5.665 0.085 5.995 0.515 ;
      RECT 5.665 1.8 5.995 2.635 ;
      RECT 5.795 1.075 7.32 1.245 ;
      RECT 5.795 1.245 5.975 1.445 ;
      RECT 6.525 0.085 6.855 0.445 ;
      RECT 6.525 1.885 6.855 2.635 ;
      RECT 7.385 0.085 7.715 0.465 ;
      RECT 7.385 1.805 7.715 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__a2111o_4
MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.955 3.775 1.74 ;
        RECT 3.505 0.29 3.995 0.825 ;
        RECT 3.505 0.825 3.775 0.955 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945 0.995 4.515 1.74 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.195 1.74 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425 0.995 2.735 2.355 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.995 2.255 1.325 ;
        RECT 1.96 1.325 2.255 2.355 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.255 0.895 2.39 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.085 0.435 0.885 ;
      RECT 0.085 1.635 0.435 2.635 ;
      RECT 1.065 0.085 2.01 0.445 ;
      RECT 1.065 0.445 1.325 0.865 ;
      RECT 1.065 1.075 1.705 1.325 ;
      RECT 1.065 1.495 1.315 2.635 ;
      RECT 1.495 0.615 3.335 0.785 ;
      RECT 1.495 0.785 1.705 1.075 ;
      RECT 1.495 1.325 1.705 1.495 ;
      RECT 1.495 1.495 1.785 2.465 ;
      RECT 2.18 0.255 2.42 0.615 ;
      RECT 2.59 0.085 2.92 0.445 ;
      RECT 3.07 1.915 4.515 2.085 ;
      RECT 3.07 2.085 3.4 2.465 ;
      RECT 3.09 0.255 3.335 0.615 ;
      RECT 3.59 2.255 3.92 2.635 ;
      RECT 4.09 2.085 4.515 2.465 ;
      RECT 4.165 0.085 4.515 0.805 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__a2111o_2
MACRO sky130_fd_sc_hd__a2111o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.29 1.325 ;
        RECT 2.985 0.285 3.54 0.845 ;
        RECT 2.985 0.845 3.29 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.51 1.025 4.01 1.29 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 0.995 2.68 2.465 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 1.05 2.22 2.465 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.29 1.05 1.72 1.29 ;
        RECT 1.515 1.29 1.72 2.465 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.255 0.465 1.62 ;
        RECT 0.135 1.62 0.39 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975 -0.065 2.145 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.565 1.815 0.895 2.635 ;
      RECT 0.635 0.085 1.31 0.47 ;
      RECT 0.695 0.65 1.915 0.655 ;
      RECT 0.695 0.655 2.805 0.825 ;
      RECT 0.695 0.825 0.915 1.465 ;
      RECT 0.695 1.465 1.345 1.645 ;
      RECT 1.135 1.645 1.345 2.46 ;
      RECT 1.585 0.26 1.915 0.65 ;
      RECT 2.085 0.085 2.43 0.485 ;
      RECT 2.6 0.26 2.805 0.655 ;
      RECT 2.86 1.495 3.99 1.665 ;
      RECT 2.86 1.665 3.145 2.46 ;
      RECT 3.325 1.835 3.54 2.635 ;
      RECT 3.715 0.085 3.955 0.76 ;
      RECT 3.72 1.665 3.99 2.46 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a2111o_1
MACRO sky130_fd_sc_hd__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 3.685 1.285 ;
        RECT 3.515 1.285 3.685 1.445 ;
        RECT 3.515 1.445 5.165 1.615 ;
        RECT 4.995 1.075 5.415 1.285 ;
        RECT 4.995 1.285 5.165 1.445 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.075 4.765 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 5.895 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.515 1.785 5.895 1.955 ;
        RECT 3.515 1.955 4.605 1.965 ;
        RECT 3.515 1.965 3.765 2.125 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 4.355 1.965 4.605 2.125 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 5.605 0.255 5.895 0.725 ;
        RECT 5.605 0.905 5.895 1.785 ;
        RECT 5.615 1.955 5.895 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.795 1.665 2.635 ;
      RECT 1.835 1.625 2.085 2.085 ;
      RECT 1.835 2.085 2.925 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.255 1.455 3.345 1.625 ;
      RECT 2.255 1.625 2.505 1.915 ;
      RECT 2.675 1.795 2.925 2.085 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 3.095 1.625 3.345 2.295 ;
      RECT 3.095 2.295 5.025 2.465 ;
      RECT 3.555 0.085 3.725 0.555 ;
      RECT 3.935 2.135 4.185 2.295 ;
      RECT 4.395 0.085 4.565 0.555 ;
      RECT 4.775 2.135 5.025 2.295 ;
      RECT 5.195 2.125 5.445 2.465 ;
      RECT 5.235 0.085 5.405 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.125 2.615 2.295 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.125 5.375 2.295 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 2.385 2.065 2.68 2.14 ;
      RECT 2.385 2.14 5.44 2.28 ;
      RECT 2.385 2.28 2.68 2.335 ;
      RECT 5.145 2.065 5.44 2.14 ;
      RECT 5.145 2.28 5.44 2.335 ;
  END
END sky130_fd_sc_hd__nor3_4
MACRO sky130_fd_sc_hd__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.185 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.075 2.965 1.285 ;
        RECT 2.375 1.285 2.64 1.625 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.595 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.755 0.255 3.085 0.725 ;
        RECT 2.835 1.455 3.595 1.625 ;
        RECT 2.835 1.625 3.045 2.125 ;
        RECT 3.135 0.905 3.595 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.465 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 1.875 0.085 2.585 0.555 ;
      RECT 2.415 1.795 2.625 2.295 ;
      RECT 3.215 1.795 3.465 2.295 ;
      RECT 3.255 0.085 3.545 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__nor3_2
MACRO sky130_fd_sc_hd__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.655 1.755 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.995 0.975 1.325 ;
        RECT 0.595 1.325 0.83 2.005 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.425 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.604500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.385 0.345 0.655 ;
        RECT 0.09 0.655 1.315 0.825 ;
        RECT 0.09 1.495 0.425 2.28 ;
        RECT 0.09 2.28 1.17 2.45 ;
        RECT 1 1.495 1.315 1.665 ;
        RECT 1 1.665 1.17 2.28 ;
        RECT 1.015 0.385 1.185 0.655 ;
        RECT 1.145 0.825 1.315 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 1.355 0.085 1.685 0.485 ;
      RECT 1.435 1.835 1.75 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__nor3_1
MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.24 1.275 ;
        RECT 0.91 1.275 1.08 1.325 ;
      LAYER mcon ;
        RECT 1.07 1.105 1.24 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.23 1.03 2.62 1.36 ;
      LAYER mcon ;
        RECT 2.45 1.105 2.62 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.25 0.955 4.625 1.275 ;
      LAYER mcon ;
        RECT 4.31 1.105 4.48 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.885 1.035 6.325 1.275 ;
      LAYER mcon ;
        RECT 6.15 1.105 6.32 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.01 1.075 1.3 1.12 ;
        RECT 1.01 1.12 6.38 1.26 ;
        RECT 1.01 1.26 1.3 1.305 ;
        RECT 2.39 1.075 2.68 1.12 ;
        RECT 2.39 1.26 2.68 1.305 ;
        RECT 4.25 1.075 4.54 1.12 ;
        RECT 4.25 1.26 4.54 1.305 ;
        RECT 6.09 1.075 6.38 1.12 ;
        RECT 6.09 1.26 6.38 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 1.445 1.7 1.88 ;
      LAYER mcon ;
        RECT 1.53 1.445 1.7 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.2 1.435 3.56 1.765 ;
      LAYER mcon ;
        RECT 3.39 1.445 3.56 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.635 1.445 6.055 1.765 ;
      LAYER mcon ;
        RECT 5.69 1.445 5.86 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.47 1.415 1.76 1.46 ;
        RECT 1.47 1.46 5.92 1.6 ;
        RECT 1.47 1.6 1.76 1.645 ;
        RECT 3.33 1.415 3.62 1.46 ;
        RECT 3.33 1.6 3.62 1.645 ;
        RECT 5.63 1.415 5.92 1.46 ;
        RECT 5.63 1.6 5.92 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.67 1.105 2.04 1.275 ;
        RECT 1.87 1.275 2.04 1.595 ;
        RECT 1.87 1.595 2.96 1.765 ;
        RECT 2.79 0.965 3.955 1.25 ;
        RECT 2.79 1.25 2.96 1.595 ;
        RECT 3.785 1.25 3.955 1.515 ;
        RECT 3.785 1.515 5.405 1.685 ;
        RECT 5.155 1.685 5.405 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.83 ;
        RECT 0.085 0.83 0.26 1.485 ;
        RECT 0.085 1.485 0.345 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.84 0.255 7.24 0.81 ;
        RECT 6.84 1.485 7.24 2.465 ;
        RECT 6.91 0.81 7.24 1.485 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 0.635 1.71 0.805 ;
      RECT 0.515 0.805 0.685 0.995 ;
      RECT 0.515 1.325 0.685 1.625 ;
      RECT 0.515 1.625 1.105 1.945 ;
      RECT 0.515 2.15 0.765 2.635 ;
      RECT 0.935 1.945 1.105 2.065 ;
      RECT 0.935 2.065 1.71 2.465 ;
      RECT 1.11 0.255 1.71 0.635 ;
      RECT 1.47 0.805 1.71 0.935 ;
      RECT 1.96 0.255 2.13 0.615 ;
      RECT 1.96 0.615 2.97 0.785 ;
      RECT 1.96 1.935 3.035 2.105 ;
      RECT 1.96 2.105 2.13 2.465 ;
      RECT 2.3 0.085 2.63 0.445 ;
      RECT 2.3 2.275 2.63 2.635 ;
      RECT 2.8 0.255 2.97 0.615 ;
      RECT 2.8 2.105 3.035 2.465 ;
      RECT 3.24 0.085 3.57 0.49 ;
      RECT 3.24 2.255 3.57 2.635 ;
      RECT 3.74 0.255 3.91 0.615 ;
      RECT 3.74 0.615 4.75 0.785 ;
      RECT 3.74 1.935 4.75 2.105 ;
      RECT 3.74 2.105 3.91 2.465 ;
      RECT 4.08 0.085 4.41 0.445 ;
      RECT 4.08 2.275 4.41 2.635 ;
      RECT 4.58 0.255 4.75 0.615 ;
      RECT 4.58 2.105 4.75 2.465 ;
      RECT 4.795 0.955 5.46 1.125 ;
      RECT 4.965 0.765 5.46 0.955 ;
      RECT 5.085 0.255 6.095 0.505 ;
      RECT 5.085 0.505 5.255 0.595 ;
      RECT 5.085 2.125 6.17 2.465 ;
      RECT 5.925 0.505 6.095 0.615 ;
      RECT 5.925 0.615 6.665 0.785 ;
      RECT 6 1.935 6.665 2.105 ;
      RECT 6 2.105 6.17 2.125 ;
      RECT 6.265 0.085 6.595 0.445 ;
      RECT 6.34 2.275 6.67 2.635 ;
      RECT 6.495 0.785 6.665 0.995 ;
      RECT 6.495 0.995 6.74 1.325 ;
      RECT 6.495 1.325 6.665 1.935 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.23 0.765 5.4 0.935 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 5.46 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 5.17 0.735 5.46 0.78 ;
      RECT 5.17 0.92 5.46 0.965 ;
  END
END sky130_fd_sc_hd__fa_1
MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 0.995 1.755 1.275 ;
        RECT 1.245 1.275 1.505 1.325 ;
      LAYER mcon ;
        RECT 1.525 1.105 1.695 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685 1.03 3.075 1.36 ;
      LAYER mcon ;
        RECT 2.905 1.105 3.075 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.72 0.955 5.08 1.275 ;
      LAYER mcon ;
        RECT 4.765 1.105 4.935 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.105 0.995 6.96 1.275 ;
      LAYER mcon ;
        RECT 6.145 1.105 6.315 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 1.755 1.12 ;
        RECT 1.465 1.12 6.375 1.26 ;
        RECT 1.465 1.26 1.755 1.305 ;
        RECT 2.845 1.075 3.135 1.12 ;
        RECT 2.845 1.26 3.135 1.305 ;
        RECT 4.705 1.075 4.995 1.12 ;
        RECT 4.705 1.26 4.995 1.305 ;
        RECT 6.085 1.075 6.375 1.12 ;
        RECT 6.085 1.26 6.375 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.445 2.155 1.69 ;
      LAYER mcon ;
        RECT 1.985 1.445 2.155 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.655 1.435 4.07 1.745 ;
      LAYER mcon ;
        RECT 3.845 1.445 4.015 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.15 1.445 6.835 1.735 ;
      LAYER mcon ;
        RECT 6.605 1.445 6.775 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.925 1.415 2.215 1.46 ;
        RECT 1.925 1.46 6.835 1.6 ;
        RECT 1.925 1.6 2.215 1.645 ;
        RECT 3.785 1.415 4.075 1.46 ;
        RECT 3.785 1.6 4.075 1.645 ;
        RECT 6.545 1.415 6.835 1.46 ;
        RECT 6.545 1.6 6.835 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.475500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125 1.105 2.495 1.275 ;
        RECT 2.325 1.275 2.495 1.57 ;
        RECT 2.325 1.57 3.415 1.74 ;
        RECT 3.245 0.965 4.465 1.25 ;
        RECT 3.245 1.25 3.415 1.57 ;
        RECT 4.295 1.25 4.465 1.435 ;
        RECT 4.295 1.435 4.655 1.515 ;
        RECT 4.295 1.515 5.92 1.685 ;
        RECT 5.67 1.355 5.92 1.515 ;
        RECT 5.67 1.685 5.92 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.735 0.69 0.905 ;
        RECT 0.085 0.905 0.37 1.415 ;
        RECT 0.085 1.415 0.735 1.585 ;
        RECT 0.52 0.315 0.85 0.485 ;
        RECT 0.52 0.485 0.69 0.735 ;
        RECT 0.565 1.585 0.735 1.78 ;
        RECT 0.565 1.78 0.81 1.95 ;
        RECT 0.6 1.95 0.81 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.523500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.395 0.255 7.725 0.485 ;
        RECT 7.395 1.795 7.645 1.965 ;
        RECT 7.395 1.965 7.565 2.465 ;
        RECT 7.475 0.485 7.725 0.735 ;
        RECT 7.475 0.735 8.195 0.905 ;
        RECT 7.475 1.415 8.195 1.585 ;
        RECT 7.475 1.585 7.645 1.795 ;
        RECT 7.97 0.905 8.195 1.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.18 0.085 0.35 0.565 ;
      RECT 0.18 1.795 0.35 2.635 ;
      RECT 0.54 1.075 1.075 1.245 ;
      RECT 0.905 0.655 2.165 0.825 ;
      RECT 0.905 0.825 1.075 1.075 ;
      RECT 0.905 1.245 1.075 1.43 ;
      RECT 0.905 1.43 1.11 1.495 ;
      RECT 0.905 1.495 1.475 1.6 ;
      RECT 0.94 1.6 1.475 1.665 ;
      RECT 0.98 2.275 1.31 2.635 ;
      RECT 1.02 0.085 1.35 0.465 ;
      RECT 1.305 1.665 1.475 1.91 ;
      RECT 1.305 1.91 2.245 2.08 ;
      RECT 1.535 0.255 2.165 0.655 ;
      RECT 1.9 2.08 2.245 2.465 ;
      RECT 1.925 0.825 2.165 0.935 ;
      RECT 2.415 0.255 2.585 0.615 ;
      RECT 2.415 0.615 3.425 0.785 ;
      RECT 2.415 1.935 3.49 2.105 ;
      RECT 2.415 2.105 2.585 2.465 ;
      RECT 2.755 0.085 3.085 0.445 ;
      RECT 2.755 2.275 3.085 2.635 ;
      RECT 3.255 0.255 3.425 0.615 ;
      RECT 3.255 2.105 3.49 2.465 ;
      RECT 3.695 0.085 4.025 0.49 ;
      RECT 3.695 1.915 4.025 2.635 ;
      RECT 4.195 0.255 4.365 0.615 ;
      RECT 4.195 0.615 5.205 0.785 ;
      RECT 4.195 1.935 5.205 2.105 ;
      RECT 4.195 2.105 4.365 2.465 ;
      RECT 4.535 0.085 4.865 0.445 ;
      RECT 4.535 2.275 4.865 2.635 ;
      RECT 5.035 0.255 5.205 0.615 ;
      RECT 5.035 2.105 5.205 2.465 ;
      RECT 5.25 0.955 5.935 1.125 ;
      RECT 5.42 0.765 5.935 0.955 ;
      RECT 5.485 2.125 6.685 2.465 ;
      RECT 5.54 0.255 6.55 0.505 ;
      RECT 5.54 0.505 5.71 0.595 ;
      RECT 6.38 0.505 6.55 0.655 ;
      RECT 6.38 0.655 7.3 0.825 ;
      RECT 6.515 1.935 7.18 2.105 ;
      RECT 6.515 2.105 6.685 2.125 ;
      RECT 6.78 0.085 7.11 0.445 ;
      RECT 6.89 2.275 7.22 2.635 ;
      RECT 7.01 1.47 7.3 1.64 ;
      RECT 7.01 1.64 7.18 1.935 ;
      RECT 7.13 0.825 7.3 1.075 ;
      RECT 7.13 1.075 7.8 1.245 ;
      RECT 7.13 1.245 7.3 1.47 ;
      RECT 7.815 1.795 7.985 2.635 ;
      RECT 7.895 0.085 8.065 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 0.765 2.155 0.935 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.685 0.765 5.855 0.935 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 1.925 0.735 2.215 0.78 ;
      RECT 1.925 0.78 5.915 0.92 ;
      RECT 1.925 0.92 2.215 0.965 ;
      RECT 5.625 0.735 5.915 0.78 ;
      RECT 5.625 0.92 5.915 0.965 ;
  END
END sky130_fd_sc_hd__fa_2
MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.08 0.995 2.68 1.275 ;
        RECT 2.08 1.275 2.34 1.325 ;
      LAYER mcon ;
        RECT 2.45 1.105 2.62 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.61 1.03 4 1.36 ;
      LAYER mcon ;
        RECT 3.83 1.105 4 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.645 0.955 6.005 1.275 ;
      LAYER mcon ;
        RECT 5.69 1.105 5.86 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.03 0.995 7.885 1.275 ;
      LAYER mcon ;
        RECT 7.07 1.105 7.24 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.39 1.075 2.68 1.12 ;
        RECT 2.39 1.12 7.3 1.26 ;
        RECT 2.39 1.26 2.68 1.305 ;
        RECT 3.77 1.075 4.06 1.12 ;
        RECT 3.77 1.26 4.06 1.305 ;
        RECT 5.63 1.075 5.92 1.12 ;
        RECT 5.63 1.26 5.92 1.305 ;
        RECT 7.01 1.075 7.3 1.12 ;
        RECT 7.01 1.26 7.3 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 1.445 3.08 1.69 ;
      LAYER mcon ;
        RECT 2.91 1.445 3.08 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.58 1.435 4.995 1.745 ;
      LAYER mcon ;
        RECT 4.77 1.445 4.94 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.075 1.445 7.76 1.735 ;
      LAYER mcon ;
        RECT 7.53 1.445 7.7 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.85 1.415 3.14 1.46 ;
        RECT 2.85 1.46 7.76 1.6 ;
        RECT 2.85 1.6 3.14 1.645 ;
        RECT 4.71 1.415 5 1.46 ;
        RECT 4.71 1.6 5 1.645 ;
        RECT 7.47 1.415 7.76 1.46 ;
        RECT 7.47 1.6 7.76 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.105 3.42 1.275 ;
        RECT 3.25 1.275 3.42 1.57 ;
        RECT 3.25 1.57 4.34 1.74 ;
        RECT 4.17 0.965 5.39 1.25 ;
        RECT 4.17 1.25 4.34 1.57 ;
        RECT 5.22 1.25 5.39 1.435 ;
        RECT 5.22 1.435 5.58 1.515 ;
        RECT 5.22 1.515 6.845 1.685 ;
        RECT 6.595 1.355 6.845 1.515 ;
        RECT 6.595 1.685 6.845 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.735 1.525 0.905 ;
        RECT 0.085 0.905 0.435 1.415 ;
        RECT 0.085 1.415 1.57 1.585 ;
        RECT 0.515 0.255 0.845 0.735 ;
        RECT 0.515 1.585 0.845 2.445 ;
        RECT 1.355 0.315 1.685 0.485 ;
        RECT 1.355 0.485 1.525 0.735 ;
        RECT 1.4 1.585 1.57 1.78 ;
        RECT 1.4 1.78 1.645 1.95 ;
        RECT 1.435 1.95 1.645 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.943000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.32 0.255 8.65 0.485 ;
        RECT 8.32 1.795 8.57 1.965 ;
        RECT 8.32 1.965 8.49 2.465 ;
        RECT 8.4 0.485 8.65 0.735 ;
        RECT 8.4 0.735 10.035 0.905 ;
        RECT 8.4 1.415 10.035 1.585 ;
        RECT 8.4 1.585 8.57 1.795 ;
        RECT 9.16 0.27 9.49 0.735 ;
        RECT 9.16 1.585 9.49 2.425 ;
        RECT 9.7 0.905 10.035 1.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.175 0.085 0.345 0.565 ;
      RECT 0.175 1.795 0.345 2.635 ;
      RECT 0.605 1.075 1.91 1.245 ;
      RECT 1.015 0.085 1.185 0.565 ;
      RECT 1.015 1.795 1.185 2.635 ;
      RECT 1.74 0.655 3.09 0.825 ;
      RECT 1.74 0.825 1.91 1.075 ;
      RECT 1.74 1.245 1.91 1.43 ;
      RECT 1.74 1.43 1.945 1.495 ;
      RECT 1.74 1.495 2.31 1.6 ;
      RECT 1.775 1.6 2.31 1.665 ;
      RECT 1.815 2.275 2.145 2.635 ;
      RECT 1.855 0.085 2.185 0.465 ;
      RECT 2.14 1.665 2.31 1.91 ;
      RECT 2.14 1.91 3.17 2.08 ;
      RECT 2.37 0.255 3.09 0.655 ;
      RECT 2.735 2.08 3.17 2.465 ;
      RECT 2.85 0.825 3.09 0.935 ;
      RECT 3.34 0.255 3.51 0.615 ;
      RECT 3.34 0.615 4.35 0.785 ;
      RECT 3.34 1.935 4.415 2.105 ;
      RECT 3.34 2.105 3.51 2.465 ;
      RECT 3.68 0.085 4.01 0.445 ;
      RECT 3.68 2.275 4.01 2.635 ;
      RECT 4.18 0.255 4.35 0.615 ;
      RECT 4.18 2.105 4.415 2.465 ;
      RECT 4.62 0.085 4.95 0.49 ;
      RECT 4.62 1.915 4.95 2.635 ;
      RECT 5.12 0.255 5.29 0.615 ;
      RECT 5.12 0.615 6.13 0.785 ;
      RECT 5.12 1.935 6.13 2.105 ;
      RECT 5.12 2.105 5.29 2.465 ;
      RECT 5.46 0.085 5.79 0.445 ;
      RECT 5.46 2.275 5.79 2.635 ;
      RECT 5.96 0.255 6.13 0.615 ;
      RECT 5.96 2.105 6.13 2.465 ;
      RECT 6.175 0.955 6.86 1.125 ;
      RECT 6.345 0.765 6.86 0.955 ;
      RECT 6.41 2.125 7.61 2.465 ;
      RECT 6.465 0.255 7.475 0.505 ;
      RECT 6.465 0.505 6.635 0.595 ;
      RECT 7.305 0.505 7.475 0.655 ;
      RECT 7.305 0.655 8.225 0.825 ;
      RECT 7.44 1.935 8.105 2.105 ;
      RECT 7.44 2.105 7.61 2.125 ;
      RECT 7.705 0.085 8.035 0.445 ;
      RECT 7.815 2.275 8.145 2.635 ;
      RECT 7.935 1.47 8.225 1.64 ;
      RECT 7.935 1.64 8.105 1.935 ;
      RECT 8.055 0.825 8.225 1.075 ;
      RECT 8.055 1.075 9.445 1.245 ;
      RECT 8.055 1.245 8.225 1.47 ;
      RECT 8.74 1.795 8.91 2.635 ;
      RECT 8.82 0.085 8.99 0.565 ;
      RECT 9.66 0.085 9.83 0.565 ;
      RECT 9.66 1.795 9.83 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.91 0.765 3.08 0.935 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.61 0.765 6.78 0.935 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
    LAYER met1 ;
      RECT 2.85 0.735 3.14 0.78 ;
      RECT 2.85 0.78 6.84 0.92 ;
      RECT 2.85 0.92 3.14 0.965 ;
      RECT 6.55 0.735 6.84 0.78 ;
      RECT 6.55 0.92 6.84 0.965 ;
  END
END sky130_fd_sc_hd__fa_4
MACRO sky130_fd_sc_hd__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.86 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.935 0.255 14.265 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.7 1.065 12.145 1.3 ;
        RECT 11.7 1.3 12.03 2.465 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 15.18 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.885 1.435 ;
        RECT -0.19 1.435 15.37 2.91 ;
        RECT 7.2 1.305 15.37 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 15.18 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 15.18 0.085 ;
      RECT 0 2.635 15.18 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 5.665 2.175 6.01 2.635 ;
      RECT 5.76 0.085 6.01 0.905 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.245 0.085 8.64 0.56 ;
      RECT 8.425 1.835 8.66 2.635 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 9.37 2.105 9.66 2.635 ;
      RECT 9.465 0.085 9.74 0.615 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.19 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.19 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.19 2.165 ;
      RECT 11.36 1.495 11.53 2.635 ;
      RECT 11.395 0.085 11.645 0.9 ;
      RECT 12.2 1.465 12.45 2.635 ;
      RECT 12.315 0.085 12.565 0.9 ;
      RECT 12.62 1.575 12.85 2.01 ;
      RECT 12.735 0.89 13.36 1.22 ;
      RECT 13.02 0.255 13.36 0.89 ;
      RECT 13.02 1.22 13.36 2.465 ;
      RECT 13.53 0.085 13.765 0.9 ;
      RECT 13.53 1.465 13.765 2.635 ;
      RECT 14.435 0.085 14.695 0.9 ;
      RECT 14.435 1.465 14.695 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 10.98 1.785 11.15 1.955 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 12.65 1.785 12.82 1.955 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.11 0.765 13.28 0.935 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 14.405 2.635 14.575 2.805 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.865 2.635 15.035 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 13.34 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 10.92 1.755 11.21 1.8 ;
      RECT 10.92 1.8 12.88 1.94 ;
      RECT 10.92 1.94 11.21 1.985 ;
      RECT 12.59 1.755 12.88 1.8 ;
      RECT 12.59 1.94 12.88 1.985 ;
      RECT 13.05 0.735 13.34 0.78 ;
      RECT 13.05 0.92 13.34 0.965 ;
  END
END sky130_fd_sc_hd__sedfxbp_2
MACRO sky130_fd_sc_hd__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525 0.255 13.855 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.7 1.065 12.145 1.41 ;
        RECT 11.7 1.41 12.03 2.465 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.885 1.435 ;
        RECT -0.19 1.435 14.45 2.91 ;
        RECT 7.2 1.305 14.45 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.26 0.085 ;
      RECT 0 2.635 14.26 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 5.665 2.175 6.01 2.635 ;
      RECT 5.76 0.085 6.01 0.905 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.245 0.085 8.64 0.56 ;
      RECT 8.425 1.835 8.66 2.635 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 9.37 2.105 9.66 2.635 ;
      RECT 9.465 0.085 9.74 0.615 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.19 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.19 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.19 2.165 ;
      RECT 11.36 1.495 11.53 2.635 ;
      RECT 11.395 0.085 11.645 0.9 ;
      RECT 12.2 1.575 12.43 2.01 ;
      RECT 12.315 0.89 12.94 1.22 ;
      RECT 12.6 0.255 12.94 0.89 ;
      RECT 12.6 1.22 12.94 2.465 ;
      RECT 13.11 0.085 13.355 0.9 ;
      RECT 13.11 1.465 13.355 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 10.98 1.785 11.15 1.955 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.23 1.785 12.4 1.955 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 12.69 0.765 12.86 0.935 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.92 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 10.92 1.755 11.21 1.8 ;
      RECT 10.92 1.8 12.46 1.94 ;
      RECT 10.92 1.94 11.21 1.985 ;
      RECT 12.17 1.755 12.46 1.8 ;
      RECT 12.17 1.94 12.46 1.985 ;
      RECT 12.63 0.735 12.92 0.78 ;
      RECT 12.63 0.92 12.92 0.965 ;
  END
END sky130_fd_sc_hd__sedfxbp_1
MACRO sky130_fd_sc_hd__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.015 1.475 1.32 ;
        RECT 0.575 1.32 1.475 1.515 ;
        RECT 0.575 1.515 3.695 1.685 ;
        RECT 3.445 0.99 3.695 1.515 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.07 3.275 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.015 5.255 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 1.855 5.15 2.025 ;
        RECT 3.935 1.445 5.835 1.7 ;
        RECT 3.935 1.7 5.15 1.855 ;
        RECT 4.03 0.615 5.835 0.845 ;
        RECT 4.08 2.025 5.15 2.085 ;
        RECT 4.08 2.085 4.29 2.465 ;
        RECT 4.96 2.085 5.15 2.465 ;
        RECT 5.425 0.845 5.835 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.12 0.615 3.86 0.82 ;
      RECT 0.12 1.82 0.405 2.635 ;
      RECT 0.55 0.085 0.88 0.445 ;
      RECT 0.575 1.915 1.67 2.085 ;
      RECT 0.575 2.085 0.81 2.465 ;
      RECT 0.98 2.255 1.31 2.635 ;
      RECT 1.41 0.085 1.74 0.445 ;
      RECT 1.48 2.085 1.67 2.275 ;
      RECT 1.48 2.275 3.46 2.465 ;
      RECT 2.27 0.085 2.6 0.445 ;
      RECT 3.13 0.085 3.46 0.445 ;
      RECT 3.63 0.255 5.65 0.445 ;
      RECT 3.63 0.445 3.86 0.615 ;
      RECT 3.63 2.195 3.91 2.635 ;
      RECT 4.46 2.255 4.79 2.635 ;
      RECT 5.32 1.88 5.65 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__o21ai_4
MACRO sky130_fd_sc_hd__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.41 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.995 0.975 1.325 ;
        RECT 0.59 1.325 0.785 2.375 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.202500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.295 1.75 1.655 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.517000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.505 1.315 1.785 ;
        RECT 0.965 1.785 1.295 2.465 ;
        RECT 1.145 0.955 1.665 1.125 ;
        RECT 1.145 1.125 1.315 1.505 ;
        RECT 1.495 0.39 1.665 0.955 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.09 0.265 0.38 0.615 ;
      RECT 0.09 0.615 1.305 0.785 ;
      RECT 0.09 1.495 0.41 2.635 ;
      RECT 0.575 0.085 0.905 0.445 ;
      RECT 1.075 0.31 1.305 0.615 ;
      RECT 1.495 1.835 1.75 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__o21ai_1
MACRO sky130_fd_sc_hd__o21ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.415 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.1 1.005 1.34 ;
        RECT 0.605 1.34 0.775 1.645 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.355 1.73 1.685 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.290500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.51 1.345 1.68 ;
        RECT 0.965 1.68 1.3 2.465 ;
        RECT 1.175 0.955 1.74 1.125 ;
        RECT 1.175 1.125 1.345 1.51 ;
        RECT 1.455 0.28 1.74 0.955 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.12 0.28 0.38 0.615 ;
      RECT 0.12 0.615 1.285 0.785 ;
      RECT 0.145 1.825 0.475 2.635 ;
      RECT 0.55 0.085 0.88 0.445 ;
      RECT 1.05 0.28 1.285 0.615 ;
      RECT 1.47 1.855 1.725 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__o21ai_0
MACRO sky130_fd_sc_hd__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 1.055 0.45 1.445 ;
        RECT 0.12 1.445 2.095 1.615 ;
        RECT 1.6 1.075 2.095 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.62 1.075 1.42 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815 0.765 3.13 1.4 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.742000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.785 2.645 1.965 ;
        RECT 0.995 1.965 1.295 2.125 ;
        RECT 2.41 1.965 2.645 2.465 ;
        RECT 2.435 0.595 2.645 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.105 0.255 0.435 0.715 ;
      RECT 0.105 0.715 2.265 0.885 ;
      RECT 0.105 1.785 0.435 2.635 ;
      RECT 0.605 1.785 0.825 2.295 ;
      RECT 0.605 2.295 1.715 2.465 ;
      RECT 0.615 0.085 0.785 0.545 ;
      RECT 0.965 0.255 1.295 0.715 ;
      RECT 1.525 0.085 1.695 0.545 ;
      RECT 1.525 2.135 1.715 2.295 ;
      RECT 1.91 2.175 2.24 2.635 ;
      RECT 1.935 0.255 3.125 0.425 ;
      RECT 1.935 0.425 2.265 0.715 ;
      RECT 2.815 0.425 3.125 0.595 ;
      RECT 2.815 1.57 3.125 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o21ai_2
MACRO sky130_fd_sc_hd__dlrbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.536250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.65 0.415 5.91 0.655 ;
        RECT 5.65 0.655 5.95 0.685 ;
        RECT 5.65 0.685 5.975 0.825 ;
        RECT 5.65 1.495 5.975 1.66 ;
        RECT 5.65 1.66 5.915 2.465 ;
        RECT 5.74 0.825 5.975 0.86 ;
        RECT 5.79 0.86 5.975 0.885 ;
        RECT 5.79 0.885 6.355 1.325 ;
        RECT 5.79 1.325 5.975 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.5 0.255 7.755 0.825 ;
        RECT 7.5 1.445 7.755 2.465 ;
        RECT 7.545 0.825 7.755 1.055 ;
        RECT 7.545 1.055 8.195 1.325 ;
        RECT 7.545 1.325 7.755 1.445 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.39 0.995 5.14 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.78 1.07 ;
      RECT 0.605 1.07 0.84 1.4 ;
      RECT 0.605 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.48 1.165 4.2 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.74 0.085 4.07 0.825 ;
      RECT 3.82 2.135 4.59 2.635 ;
      RECT 3.84 1.495 5.48 1.665 ;
      RECT 3.84 1.665 4.93 1.865 ;
      RECT 4.34 0.415 4.56 0.655 ;
      RECT 4.34 0.655 5.48 0.825 ;
      RECT 4.76 1.865 4.93 2.435 ;
      RECT 5.1 0.085 5.48 0.485 ;
      RECT 5.1 1.855 5.35 2.635 ;
      RECT 5.31 0.825 5.48 0.995 ;
      RECT 5.31 0.995 5.62 1.325 ;
      RECT 5.31 1.325 5.48 1.495 ;
      RECT 6.085 0.085 6.355 0.545 ;
      RECT 6.085 1.83 6.355 2.635 ;
      RECT 6.525 0.255 6.855 0.995 ;
      RECT 6.525 0.995 7.375 1.325 ;
      RECT 6.525 1.325 6.855 2.465 ;
      RECT 7.025 0.085 7.33 0.545 ;
      RECT 7.035 1.835 7.33 2.635 ;
      RECT 7.925 0.085 8.195 0.885 ;
      RECT 7.925 1.495 8.195 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrbn_2
MACRO sky130_fd_sc_hd__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.38 2.465 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475 0.255 7.735 0.595 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.56 0.595 7.735 1.785 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.47 0.995 5.455 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.3 1.165 ;
      RECT 3.48 1.165 4.3 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.74 0.085 4.07 0.53 ;
      RECT 3.82 2.135 4.09 2.635 ;
      RECT 3.84 1.535 5.875 1.765 ;
      RECT 3.84 1.765 4.97 1.865 ;
      RECT 4.24 0.255 4.54 0.655 ;
      RECT 4.24 0.655 5.875 0.825 ;
      RECT 4.26 2.135 4.59 2.635 ;
      RECT 4.76 1.865 4.97 2.435 ;
      RECT 5.135 0.085 5.875 0.485 ;
      RECT 5.15 1.935 5.89 2.635 ;
      RECT 5.625 0.825 5.875 1.535 ;
      RECT 6.58 0.255 6.75 0.985 ;
      RECT 6.58 0.985 6.83 0.995 ;
      RECT 6.58 0.995 7.39 1.325 ;
      RECT 6.58 1.325 6.83 2.465 ;
      RECT 6.975 0.085 7.305 0.465 ;
      RECT 7.01 1.835 7.305 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrbn_1
MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcin_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.34 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.665 1.74 1.325 ;
      LAYER mcon ;
        RECT 1.525 0.765 1.695 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.24 0.645 4.49 1.325 ;
      LAYER mcon ;
        RECT 4.285 0.765 4.455 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 0.735 1.755 0.78 ;
        RECT 1.465 0.78 4.515 0.92 ;
        RECT 1.465 0.92 1.755 0.965 ;
        RECT 4.225 0.735 4.515 0.78 ;
        RECT 4.225 0.92 4.515 0.965 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.52 1.075 10.965 1.275 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.6 0.755 6.925 0.925 ;
        RECT 6.6 0.925 6.87 1.675 ;
        RECT 6.7 1.675 6.87 1.785 ;
        RECT 6.755 0.595 6.925 0.755 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.255 12.335 0.825 ;
        RECT 12 1.785 12.335 2.465 ;
        RECT 12.125 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.61 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.42 0.085 ;
      RECT 0 2.635 12.42 2.805 ;
      RECT 0.085 0.735 0.43 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.44 1.84 ;
      RECT 0.085 1.84 1.11 2.01 ;
      RECT 0.085 2.01 0.43 2.465 ;
      RECT 0.1 0.255 0.43 0.735 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.6 2.18 0.77 2.635 ;
      RECT 0.61 0.735 1.325 0.905 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.5 ;
      RECT 0.61 1.5 1.45 1.67 ;
      RECT 0.63 0.085 0.8 0.545 ;
      RECT 0.94 2.01 1.11 2.215 ;
      RECT 0.94 2.215 1.97 2.295 ;
      RECT 0.94 2.295 3.515 2.385 ;
      RECT 0.995 0.255 3.39 0.425 ;
      RECT 0.995 0.425 2.1 0.465 ;
      RECT 0.995 0.465 1.325 0.735 ;
      RECT 1.28 1.67 1.45 1.785 ;
      RECT 1.28 1.785 2.05 1.955 ;
      RECT 1.28 1.955 1.45 2.045 ;
      RECT 1.715 2.385 3.515 2.465 ;
      RECT 1.985 0.675 2.39 1.35 ;
      RECT 2.22 0.595 2.39 0.675 ;
      RECT 2.22 1.35 2.39 1.785 ;
      RECT 2.515 0.425 3.39 0.465 ;
      RECT 2.565 1.785 2.895 2.045 ;
      RECT 2.62 0.655 3.025 0.735 ;
      RECT 2.62 0.735 3.135 0.755 ;
      RECT 2.62 0.755 3.73 0.905 ;
      RECT 2.64 1.075 2.97 1.095 ;
      RECT 2.64 1.095 3.12 1.245 ;
      RECT 2.8 1.245 3.12 1.265 ;
      RECT 2.95 1.265 3.12 1.615 ;
      RECT 3.055 0.905 3.73 0.925 ;
      RECT 3.215 0.465 3.39 0.585 ;
      RECT 3.245 2.11 3.46 2.295 ;
      RECT 3.29 0.925 3.46 2.11 ;
      RECT 3.56 0.255 4.57 0.425 ;
      RECT 3.56 0.425 3.73 0.755 ;
      RECT 3.71 1.15 4.07 1.32 ;
      RECT 3.71 1.32 3.88 2.29 ;
      RECT 3.71 2.29 5.065 2.46 ;
      RECT 3.9 0.595 4.07 1.15 ;
      RECT 4.08 1.695 4.445 2.12 ;
      RECT 4.24 0.425 4.57 0.475 ;
      RECT 4.69 1.385 5.17 1.725 ;
      RECT 4.815 1.895 5.995 2.065 ;
      RECT 4.815 2.065 5.065 2.29 ;
      RECT 4.83 0.51 5 0.995 ;
      RECT 4.83 0.995 5.63 1.325 ;
      RECT 4.83 1.325 5.17 1.385 ;
      RECT 5.18 0.085 5.51 0.805 ;
      RECT 5.26 2.235 5.59 2.635 ;
      RECT 5.635 1.555 6.37 1.725 ;
      RECT 5.68 0.38 5.97 0.815 ;
      RECT 5.8 0.815 5.97 1.555 ;
      RECT 5.825 2.065 5.995 2.295 ;
      RECT 5.825 2.295 7.95 2.465 ;
      RECT 6.14 0.74 6.425 1.325 ;
      RECT 6.2 1.725 6.37 1.895 ;
      RECT 6.2 1.895 6.53 1.955 ;
      RECT 6.2 1.955 7.21 2.125 ;
      RECT 6.255 0.255 7.695 0.425 ;
      RECT 6.255 0.425 6.585 0.57 ;
      RECT 7.04 1.06 7.27 1.23 ;
      RECT 7.04 1.23 7.21 1.955 ;
      RECT 7.1 0.595 7.35 0.925 ;
      RECT 7.1 0.925 7.27 1.06 ;
      RECT 7.38 1.36 7.61 1.53 ;
      RECT 7.38 1.53 7.55 2.125 ;
      RECT 7.44 1.105 7.695 1.29 ;
      RECT 7.44 1.29 7.61 1.36 ;
      RECT 7.52 0.425 7.695 1.105 ;
      RECT 7.78 1.55 8.035 1.72 ;
      RECT 7.78 1.72 7.95 2.295 ;
      RECT 7.865 0.255 9.98 0.425 ;
      RECT 7.865 0.425 8.035 0.74 ;
      RECT 7.865 0.995 8.035 1.55 ;
      RECT 8.22 1.955 8.39 2.295 ;
      RECT 8.22 2.295 9.41 2.465 ;
      RECT 8.305 0.595 8.555 0.925 ;
      RECT 8.375 0.925 8.555 1.445 ;
      RECT 8.375 1.445 8.67 1.53 ;
      RECT 8.375 1.53 8.89 1.785 ;
      RECT 8.56 1.785 8.89 2.125 ;
      RECT 8.725 0.595 9.41 0.765 ;
      RECT 8.835 0.995 9.07 1.325 ;
      RECT 9.24 0.765 9.41 1.875 ;
      RECT 9.24 1.875 10.885 2.025 ;
      RECT 9.24 2.025 10.145 2.03 ;
      RECT 9.24 2.03 10.13 2.035 ;
      RECT 9.24 2.035 10.12 2.04 ;
      RECT 9.24 2.04 10.105 2.045 ;
      RECT 9.24 2.045 9.41 2.295 ;
      RECT 9.64 0.425 9.98 0.825 ;
      RECT 9.64 0.825 9.81 1.535 ;
      RECT 9.64 1.535 10.01 1.705 ;
      RECT 9.98 0.995 10.35 1.325 ;
      RECT 10.055 1.87 10.885 1.875 ;
      RECT 10.07 1.865 10.885 1.87 ;
      RECT 10.085 1.86 10.885 1.865 ;
      RECT 10.1 1.855 10.885 1.86 ;
      RECT 10.18 0.085 10.35 0.565 ;
      RECT 10.18 0.735 10.91 0.905 ;
      RECT 10.18 0.905 10.35 0.995 ;
      RECT 10.18 1.325 10.35 1.445 ;
      RECT 10.18 1.445 10.885 1.855 ;
      RECT 10.19 2.195 10.36 2.635 ;
      RECT 10.53 0.285 10.91 0.735 ;
      RECT 10.535 2.025 10.885 2.465 ;
      RECT 11.075 1.455 11.405 2.465 ;
      RECT 11.155 0.27 11.325 0.68 ;
      RECT 11.155 0.68 11.405 1.455 ;
      RECT 11.495 0.085 11.825 0.51 ;
      RECT 11.575 1.785 11.83 2.635 ;
      RECT 11.645 0.995 11.955 1.615 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.88 1.785 2.05 1.955 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 1.105 2.155 1.275 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.57 1.785 2.74 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.95 1.445 3.12 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.14 1.785 4.31 1.955 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.76 1.445 4.93 1.615 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.14 1.105 6.31 1.275 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.52 0.765 7.69 0.935 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.44 1.445 8.61 1.615 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.9 1.105 9.07 1.275 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.22 0.765 11.39 0.935 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 11.68 1.445 11.85 1.615 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
    LAYER met1 ;
      RECT 1.82 1.755 2.11 1.8 ;
      RECT 1.82 1.8 4.37 1.94 ;
      RECT 1.82 1.94 2.11 1.985 ;
      RECT 1.925 1.075 2.215 1.12 ;
      RECT 1.925 1.12 9.13 1.26 ;
      RECT 1.925 1.26 2.215 1.305 ;
      RECT 2.51 1.755 2.8 1.8 ;
      RECT 2.51 1.94 2.8 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.46 4.99 1.6 ;
      RECT 2.89 1.6 3.18 1.645 ;
      RECT 4.08 1.755 4.37 1.8 ;
      RECT 4.08 1.94 4.37 1.985 ;
      RECT 4.7 1.415 4.99 1.46 ;
      RECT 4.7 1.6 4.99 1.645 ;
      RECT 6.08 1.075 6.37 1.12 ;
      RECT 6.08 1.26 6.37 1.305 ;
      RECT 7.46 0.735 7.75 0.78 ;
      RECT 7.46 0.78 11.45 0.92 ;
      RECT 7.46 0.92 7.75 0.965 ;
      RECT 8.38 1.415 8.67 1.46 ;
      RECT 8.38 1.46 11.91 1.6 ;
      RECT 8.38 1.6 8.67 1.645 ;
      RECT 8.84 1.075 9.13 1.12 ;
      RECT 8.84 1.26 9.13 1.305 ;
      RECT 11.16 0.735 11.45 0.78 ;
      RECT 11.16 0.92 11.45 0.965 ;
      RECT 11.62 1.415 11.91 1.46 ;
      RECT 11.62 1.6 11.91 1.645 ;
  END
END sky130_fd_sc_hd__fahcin_1
MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.5 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.18 0.825 ;
        RECT 1.645 1.845 2.18 2.465 ;
        RECT 1.865 0.825 2.18 1.845 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.25 0.085 0.49 0.595 ;
      RECT 0.27 1.495 1.695 1.665 ;
      RECT 0.27 1.665 0.66 1.84 ;
      RECT 0.67 0.265 0.95 0.595 ;
      RECT 0.67 0.595 0.84 1.495 ;
      RECT 1.145 1.835 1.475 2.635 ;
      RECT 1.18 0.085 1.395 0.595 ;
      RECT 1.525 0.995 1.695 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__or2_1
MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.765 0.345 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.835 2.215 2.005 ;
        RECT 1.44 2.005 1.77 2.465 ;
        RECT 1.52 0.385 1.69 0.655 ;
        RECT 1.52 0.655 2.215 0.825 ;
        RECT 1.785 0.825 2.215 1.835 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.105 0.085 0.345 0.595 ;
      RECT 0.155 1.495 1.615 1.665 ;
      RECT 0.155 1.665 0.515 1.84 ;
      RECT 0.515 0.255 0.805 0.595 ;
      RECT 0.515 0.595 0.695 1.495 ;
      RECT 1.035 0.085 1.35 0.595 ;
      RECT 1.1 1.835 1.27 2.635 ;
      RECT 1.445 0.995 1.615 1.495 ;
      RECT 1.86 0.085 2.19 0.485 ;
      RECT 1.94 2.175 2.11 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__or2_2
MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.995 1.24 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.765 0.345 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 0.265 1.77 0.735 ;
        RECT 1.44 0.735 3.135 0.905 ;
        RECT 1.44 1.835 2.61 2.005 ;
        RECT 1.44 2.005 1.77 2.465 ;
        RECT 2.28 0.265 2.61 0.735 ;
        RECT 2.28 1.495 3.135 1.665 ;
        RECT 2.28 1.665 2.61 1.835 ;
        RECT 2.28 2.005 2.61 2.465 ;
        RECT 2.79 0.905 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.105 0.085 0.345 0.595 ;
      RECT 0.155 1.495 1.615 1.665 ;
      RECT 0.155 1.665 0.515 2.465 ;
      RECT 0.515 0.29 0.845 0.825 ;
      RECT 0.515 0.825 0.695 1.495 ;
      RECT 1.06 0.085 1.23 0.825 ;
      RECT 1.06 1.835 1.23 2.635 ;
      RECT 1.41 1.075 2.62 1.245 ;
      RECT 1.41 1.245 1.615 1.495 ;
      RECT 1.94 0.085 2.11 0.565 ;
      RECT 1.94 2.175 2.11 2.635 ;
      RECT 2.78 0.085 2.95 0.565 ;
      RECT 2.78 1.835 2.95 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__or2_4
MACRO sky130_fd_sc_hd__or2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.995 1.335 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.5 1.615 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.326800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.525 2.18 0.825 ;
        RECT 1.645 2.135 2.18 2.465 ;
        RECT 1.865 0.825 2.18 2.135 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.25 0.085 0.49 0.825 ;
      RECT 0.27 1.785 1.695 1.955 ;
      RECT 0.27 1.955 0.66 2.13 ;
      RECT 0.67 0.425 0.95 0.825 ;
      RECT 0.67 0.825 0.84 1.785 ;
      RECT 1.145 2.125 1.475 2.635 ;
      RECT 1.18 0.085 1.395 0.825 ;
      RECT 1.525 0.995 1.695 1.785 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__or2_0
MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 1.74 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.915 1.295 2.465 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.275 1.91 0.605 2.635 ;
      RECT 0.775 0.085 1.115 0.745 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__conb_1
MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.275 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.995 1.785 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.995 1.285 1.615 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.795 1.615 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.871000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.655 1.925 0.825 ;
        RECT 0.085 0.825 0.345 2.45 ;
        RECT 0.855 0.3 1.055 0.655 ;
        RECT 1.725 0.31 1.925 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.355 0.085 0.685 0.48 ;
      RECT 0.525 0.995 0.745 1.795 ;
      RECT 0.525 1.795 3.135 2.005 ;
      RECT 1.225 0.085 1.555 0.485 ;
      RECT 2.095 0.085 2.425 0.825 ;
      RECT 2.095 2.185 2.425 2.635 ;
      RECT 2.66 0.405 2.83 0.655 ;
      RECT 2.66 0.655 3.135 0.825 ;
      RECT 2.965 0.825 3.135 1.795 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__nor4b_1
MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.075 1.805 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 3.75 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 5.685 1.285 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.81 1.075 8.655 1.285 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 7.245 0.905 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.195 0.255 2.525 0.725 ;
        RECT 3.035 0.255 3.365 0.725 ;
        RECT 4.395 0.255 4.725 0.725 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.115 0.905 6.465 1.455 ;
        RECT 6.115 1.455 7.205 1.625 ;
        RECT 6.115 1.625 6.365 2.125 ;
        RECT 6.915 0.255 7.245 0.725 ;
        RECT 6.955 1.625 7.205 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.095 1.455 2.065 1.625 ;
      RECT 0.095 1.625 0.425 2.465 ;
      RECT 0.175 0.085 0.345 0.895 ;
      RECT 0.595 1.795 0.805 2.635 ;
      RECT 0.975 1.625 1.225 2.465 ;
      RECT 1.015 0.085 1.185 0.555 ;
      RECT 1.395 1.795 1.645 2.635 ;
      RECT 1.815 1.625 2.065 2.295 ;
      RECT 1.815 2.295 3.745 2.465 ;
      RECT 1.855 0.085 2.025 0.555 ;
      RECT 2.235 1.455 5.525 1.625 ;
      RECT 2.235 1.625 2.485 2.125 ;
      RECT 2.655 1.795 2.905 2.295 ;
      RECT 2.695 0.085 2.865 0.555 ;
      RECT 3.075 1.625 3.325 2.125 ;
      RECT 3.495 1.795 3.745 2.295 ;
      RECT 3.535 0.085 4.225 0.555 ;
      RECT 4.015 1.795 4.265 2.295 ;
      RECT 4.015 2.295 7.625 2.465 ;
      RECT 4.435 1.625 4.685 2.125 ;
      RECT 4.855 1.795 5.105 2.295 ;
      RECT 4.895 0.085 5.065 0.555 ;
      RECT 5.275 1.625 5.525 2.125 ;
      RECT 5.695 1.455 5.945 2.295 ;
      RECT 5.735 0.085 5.905 0.555 ;
      RECT 6.535 1.795 6.785 2.295 ;
      RECT 6.575 0.085 6.745 0.555 ;
      RECT 6.635 1.075 7.64 1.285 ;
      RECT 7.375 1.795 7.625 2.295 ;
      RECT 7.415 0.085 7.585 0.555 ;
      RECT 7.47 0.735 8.185 0.905 ;
      RECT 7.47 0.905 7.64 1.075 ;
      RECT 7.47 1.285 7.64 1.455 ;
      RECT 7.47 1.455 8.185 1.625 ;
      RECT 7.81 0.255 8.185 0.735 ;
      RECT 7.85 1.625 8.185 2.465 ;
      RECT 8.355 0.085 8.585 0.905 ;
      RECT 8.355 1.455 8.585 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
  END
END sky130_fd_sc_hd__nor4b_4
MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 1.24 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 1.075 2.635 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.075 3.535 1.285 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.805 1.075 5.435 1.285 ;
        RECT 5.185 1.285 5.435 1.955 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 3.92 0.905 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.75 0.255 3.08 0.725 ;
        RECT 3.59 0.255 3.92 0.725 ;
        RECT 3.63 1.455 4.035 1.625 ;
        RECT 3.63 1.625 3.88 2.125 ;
        RECT 3.715 0.905 3.92 1.075 ;
        RECT 3.715 1.075 4.035 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.085 0.085 0.345 0.905 ;
      RECT 0.085 1.455 2.105 1.625 ;
      RECT 0.085 1.625 0.425 2.465 ;
      RECT 0.595 1.795 0.805 2.635 ;
      RECT 0.975 1.625 1.225 2.465 ;
      RECT 1.015 0.085 1.185 0.555 ;
      RECT 1.395 1.795 1.605 2.295 ;
      RECT 1.395 2.295 3.04 2.465 ;
      RECT 1.775 1.625 2.105 2.125 ;
      RECT 1.855 0.085 2.58 0.555 ;
      RECT 2.275 1.455 3.46 1.625 ;
      RECT 2.275 1.625 2.66 2.125 ;
      RECT 2.83 1.795 3.04 2.295 ;
      RECT 3.21 1.625 3.46 2.295 ;
      RECT 3.21 2.295 4.295 2.465 ;
      RECT 3.25 0.085 3.42 0.555 ;
      RECT 4.05 1.795 4.295 2.295 ;
      RECT 4.09 0.085 4.295 0.895 ;
      RECT 4.32 1.075 4.635 1.245 ;
      RECT 4.465 0.38 4.82 0.905 ;
      RECT 4.465 0.905 4.635 1.075 ;
      RECT 4.465 1.245 4.635 2.035 ;
      RECT 4.465 2.035 4.82 2.45 ;
      RECT 4.99 0.085 5.24 0.825 ;
      RECT 4.99 2.135 5.24 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__nor4b_2
MACRO sky130_fd_sc_hd__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045 1.075 7.455 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.225 0.995 6.395 1.445 ;
        RECT 6.225 1.445 6.805 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.075 2.18 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.345 0.925 ;
        RECT 0.085 0.925 0.33 1.44 ;
        RECT 0.085 1.44 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.5 0.995 0.705 1.325 ;
      RECT 0.515 0.085 0.765 0.525 ;
      RECT 0.53 0.695 1.105 0.865 ;
      RECT 0.53 0.865 0.705 0.995 ;
      RECT 0.535 1.325 0.705 1.875 ;
      RECT 0.535 1.875 1.22 2.045 ;
      RECT 0.535 2.215 0.87 2.635 ;
      RECT 0.935 0.255 2.505 0.425 ;
      RECT 0.935 0.425 1.105 0.695 ;
      RECT 0.935 1.535 2.52 1.705 ;
      RECT 1.05 2.045 1.22 2.235 ;
      RECT 1.05 2.235 2.52 2.405 ;
      RECT 1.275 0.595 1.445 1.535 ;
      RECT 1.56 1.895 4.06 2.065 ;
      RECT 1.745 0.625 2.965 0.795 ;
      RECT 1.745 0.795 2.125 0.905 ;
      RECT 2.07 0.425 2.505 0.455 ;
      RECT 2.35 0.995 2.625 1.325 ;
      RECT 2.35 1.325 2.52 1.535 ;
      RECT 2.675 0.285 3.305 0.455 ;
      RECT 2.69 1.525 3.075 1.695 ;
      RECT 2.795 0.795 2.965 1.375 ;
      RECT 2.795 1.375 3.075 1.525 ;
      RECT 3.135 0.455 3.305 1.035 ;
      RECT 3.135 1.035 3.415 1.205 ;
      RECT 3.225 2.235 3.555 2.635 ;
      RECT 3.245 1.205 3.415 1.895 ;
      RECT 3.475 0.085 3.645 0.865 ;
      RECT 3.645 1.445 4.065 1.715 ;
      RECT 3.825 0.415 4.065 1.445 ;
      RECT 3.89 2.065 4.06 2.275 ;
      RECT 3.89 2.275 6.985 2.445 ;
      RECT 4.245 0.265 4.655 0.485 ;
      RECT 4.245 0.485 4.455 0.595 ;
      RECT 4.245 0.595 4.415 2.105 ;
      RECT 4.585 0.72 4.995 0.825 ;
      RECT 4.585 0.825 4.795 0.89 ;
      RECT 4.585 0.89 4.755 2.275 ;
      RECT 4.625 0.655 4.995 0.72 ;
      RECT 4.825 0.32 4.995 0.655 ;
      RECT 4.935 1.445 5.715 1.615 ;
      RECT 4.935 1.615 5.35 2.045 ;
      RECT 4.95 0.995 5.375 1.27 ;
      RECT 5.165 0.63 5.375 0.995 ;
      RECT 5.545 0.255 6.69 0.425 ;
      RECT 5.545 0.425 5.715 1.445 ;
      RECT 5.885 0.595 6.055 1.935 ;
      RECT 5.885 1.935 8.195 2.105 ;
      RECT 6.225 0.425 6.69 0.465 ;
      RECT 6.565 0.73 6.77 0.945 ;
      RECT 6.565 0.945 6.875 1.275 ;
      RECT 6.975 1.495 7.795 1.705 ;
      RECT 7.015 0.295 7.305 0.735 ;
      RECT 7.015 0.735 7.795 0.75 ;
      RECT 7.055 0.75 7.795 0.905 ;
      RECT 7.395 2.275 7.73 2.635 ;
      RECT 7.475 0.085 7.645 0.565 ;
      RECT 7.625 0.905 7.795 0.995 ;
      RECT 7.625 0.995 7.855 1.325 ;
      RECT 7.625 1.325 7.795 1.495 ;
      RECT 7.71 1.875 8.195 1.935 ;
      RECT 7.895 0.255 8.195 0.585 ;
      RECT 7.9 2.105 8.195 2.465 ;
      RECT 8.025 0.585 8.195 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.445 3.075 1.615 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 0.765 3.995 0.935 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 0.425 4.455 0.595 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.205 1.445 5.375 1.615 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 0.765 6.755 0.935 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 0.425 7.215 0.595 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 2.845 1.415 3.135 1.46 ;
      RECT 2.845 1.46 5.435 1.6 ;
      RECT 2.845 1.6 3.135 1.645 ;
      RECT 3.765 0.735 4.055 0.78 ;
      RECT 3.765 0.78 6.815 0.92 ;
      RECT 3.765 0.92 4.055 0.965 ;
      RECT 4.225 0.395 4.515 0.44 ;
      RECT 4.225 0.44 7.275 0.58 ;
      RECT 4.225 0.58 4.515 0.625 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.145 1.415 5.435 1.46 ;
      RECT 5.145 1.6 5.435 1.645 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
      RECT 6.985 0.395 7.275 0.44 ;
      RECT 6.985 0.58 7.275 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_1
MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425 1.075 8.835 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605 0.995 7.775 1.445 ;
        RECT 7.605 1.445 8.185 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995 1.075 3.56 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 0.375 0.875 0.995 ;
        RECT 0.625 0.995 1.71 1.325 ;
        RECT 0.625 1.325 0.955 2.425 ;
        RECT 1.465 0.35 1.725 0.925 ;
        RECT 1.465 0.925 1.71 0.995 ;
        RECT 1.465 1.325 1.71 1.44 ;
        RECT 1.465 1.44 1.745 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.285 0.085 0.455 0.735 ;
      RECT 0.285 1.49 0.455 2.635 ;
      RECT 1.125 0.085 1.295 0.735 ;
      RECT 1.125 1.495 1.295 2.635 ;
      RECT 1.88 0.995 2.085 1.325 ;
      RECT 1.895 0.085 2.145 0.525 ;
      RECT 1.91 0.695 2.485 0.865 ;
      RECT 1.91 0.865 2.085 0.995 ;
      RECT 1.915 1.325 2.085 1.875 ;
      RECT 1.915 1.875 2.6 2.045 ;
      RECT 1.915 2.215 2.25 2.635 ;
      RECT 2.315 0.255 3.885 0.425 ;
      RECT 2.315 0.425 2.485 0.695 ;
      RECT 2.315 1.535 3.9 1.705 ;
      RECT 2.43 2.045 2.6 2.235 ;
      RECT 2.43 2.235 3.9 2.405 ;
      RECT 2.655 0.595 2.825 1.535 ;
      RECT 2.94 1.895 5.44 2.065 ;
      RECT 3.125 0.625 4.345 0.795 ;
      RECT 3.125 0.795 3.505 0.905 ;
      RECT 3.45 0.425 3.885 0.455 ;
      RECT 3.73 0.995 4.005 1.325 ;
      RECT 3.73 1.325 3.9 1.535 ;
      RECT 4.055 0.285 4.685 0.455 ;
      RECT 4.07 1.525 4.455 1.695 ;
      RECT 4.175 0.795 4.345 1.375 ;
      RECT 4.175 1.375 4.455 1.525 ;
      RECT 4.515 0.455 4.685 1.035 ;
      RECT 4.515 1.035 4.795 1.205 ;
      RECT 4.605 2.235 4.935 2.635 ;
      RECT 4.625 1.205 4.795 1.895 ;
      RECT 4.855 0.085 5.025 0.865 ;
      RECT 5.025 1.445 5.445 1.715 ;
      RECT 5.205 0.415 5.445 1.445 ;
      RECT 5.27 2.065 5.44 2.275 ;
      RECT 5.27 2.275 8.365 2.445 ;
      RECT 5.625 0.265 6.035 0.485 ;
      RECT 5.625 0.485 5.835 0.595 ;
      RECT 5.625 0.595 5.795 2.105 ;
      RECT 5.965 0.72 6.375 0.825 ;
      RECT 5.965 0.825 6.175 0.89 ;
      RECT 5.965 0.89 6.135 2.275 ;
      RECT 6.005 0.655 6.375 0.72 ;
      RECT 6.205 0.32 6.375 0.655 ;
      RECT 6.315 1.445 7.095 1.615 ;
      RECT 6.315 1.615 6.73 2.045 ;
      RECT 6.33 0.995 6.755 1.27 ;
      RECT 6.545 0.63 6.755 0.995 ;
      RECT 6.925 0.255 8.07 0.425 ;
      RECT 6.925 0.425 7.095 1.445 ;
      RECT 7.265 0.595 7.435 1.935 ;
      RECT 7.265 1.935 9.575 2.105 ;
      RECT 7.605 0.425 8.07 0.465 ;
      RECT 7.945 0.73 8.15 0.945 ;
      RECT 7.945 0.945 8.255 1.275 ;
      RECT 8.355 1.495 9.175 1.705 ;
      RECT 8.395 0.295 8.685 0.735 ;
      RECT 8.395 0.735 9.175 0.75 ;
      RECT 8.435 0.75 9.175 0.905 ;
      RECT 8.775 2.275 9.11 2.635 ;
      RECT 8.855 0.085 9.025 0.565 ;
      RECT 9.005 0.905 9.175 0.995 ;
      RECT 9.005 0.995 9.235 1.325 ;
      RECT 9.005 1.325 9.175 1.495 ;
      RECT 9.09 1.875 9.575 1.935 ;
      RECT 9.275 0.255 9.575 0.585 ;
      RECT 9.28 2.105 9.575 2.465 ;
      RECT 9.405 0.585 9.575 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.445 4.455 1.615 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 0.425 5.835 0.595 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 0.765 6.755 0.935 ;
      RECT 6.585 1.445 6.755 1.615 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 0.765 8.135 0.935 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 0.425 8.595 0.595 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 4.225 1.415 4.515 1.46 ;
      RECT 4.225 1.46 6.815 1.6 ;
      RECT 4.225 1.6 4.515 1.645 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.78 8.195 0.92 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.605 0.395 5.895 0.44 ;
      RECT 5.605 0.44 8.655 0.58 ;
      RECT 5.605 0.58 5.895 0.625 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
      RECT 6.525 1.415 6.815 1.46 ;
      RECT 6.525 1.6 6.815 1.645 ;
      RECT 7.905 0.735 8.195 0.78 ;
      RECT 7.905 0.92 8.195 0.965 ;
      RECT 8.365 0.395 8.655 0.44 ;
      RECT 8.365 0.58 8.655 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_4
MACRO sky130_fd_sc_hd__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685 0.995 6.855 1.445 ;
        RECT 6.685 1.445 7.265 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 2.64 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.35 0.805 0.925 ;
        RECT 0.545 0.925 0.79 1.44 ;
        RECT 0.545 1.44 0.825 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.085 0.085 0.375 0.735 ;
      RECT 0.085 1.49 0.375 2.635 ;
      RECT 0.96 0.995 1.165 1.325 ;
      RECT 0.975 0.085 1.225 0.525 ;
      RECT 0.99 0.695 1.565 0.865 ;
      RECT 0.99 0.865 1.165 0.995 ;
      RECT 0.995 1.325 1.165 1.875 ;
      RECT 0.995 1.875 1.68 2.045 ;
      RECT 0.995 2.215 1.33 2.635 ;
      RECT 1.395 0.255 2.965 0.425 ;
      RECT 1.395 0.425 1.565 0.695 ;
      RECT 1.395 1.535 2.98 1.705 ;
      RECT 1.51 2.045 1.68 2.235 ;
      RECT 1.51 2.235 2.98 2.405 ;
      RECT 1.735 0.595 1.905 1.535 ;
      RECT 2.02 1.895 4.52 2.065 ;
      RECT 2.205 0.625 3.425 0.795 ;
      RECT 2.205 0.795 2.585 0.905 ;
      RECT 2.53 0.425 2.965 0.455 ;
      RECT 2.81 0.995 3.085 1.325 ;
      RECT 2.81 1.325 2.98 1.535 ;
      RECT 3.135 0.285 3.765 0.455 ;
      RECT 3.15 1.525 3.535 1.695 ;
      RECT 3.255 0.795 3.425 1.375 ;
      RECT 3.255 1.375 3.535 1.525 ;
      RECT 3.595 0.455 3.765 1.035 ;
      RECT 3.595 1.035 3.875 1.205 ;
      RECT 3.685 2.235 4.015 2.635 ;
      RECT 3.705 1.205 3.875 1.895 ;
      RECT 3.935 0.085 4.105 0.865 ;
      RECT 4.105 1.445 4.525 1.715 ;
      RECT 4.285 0.415 4.525 1.445 ;
      RECT 4.35 2.065 4.52 2.275 ;
      RECT 4.35 2.275 7.445 2.445 ;
      RECT 4.705 0.265 5.115 0.485 ;
      RECT 4.705 0.485 4.915 0.595 ;
      RECT 4.705 0.595 4.875 2.105 ;
      RECT 5.045 0.72 5.455 0.825 ;
      RECT 5.045 0.825 5.255 0.89 ;
      RECT 5.045 0.89 5.215 2.275 ;
      RECT 5.085 0.655 5.455 0.72 ;
      RECT 5.285 0.32 5.455 0.655 ;
      RECT 5.395 1.445 6.175 1.615 ;
      RECT 5.395 1.615 5.81 2.045 ;
      RECT 5.41 0.995 5.835 1.27 ;
      RECT 5.625 0.63 5.835 0.995 ;
      RECT 6.005 0.255 7.15 0.425 ;
      RECT 6.005 0.425 6.175 1.445 ;
      RECT 6.345 0.595 6.515 1.935 ;
      RECT 6.345 1.935 8.655 2.105 ;
      RECT 6.685 0.425 7.15 0.465 ;
      RECT 7.025 0.73 7.23 0.945 ;
      RECT 7.025 0.945 7.335 1.275 ;
      RECT 7.435 1.495 8.255 1.705 ;
      RECT 7.475 0.295 7.765 0.735 ;
      RECT 7.475 0.735 8.255 0.75 ;
      RECT 7.515 0.75 8.255 0.905 ;
      RECT 7.855 2.275 8.19 2.635 ;
      RECT 7.935 0.085 8.105 0.565 ;
      RECT 8.085 0.905 8.255 0.995 ;
      RECT 8.085 0.995 8.315 1.325 ;
      RECT 8.085 1.325 8.255 1.495 ;
      RECT 8.17 1.875 8.655 1.935 ;
      RECT 8.355 0.255 8.655 0.585 ;
      RECT 8.36 2.105 8.655 2.465 ;
      RECT 8.485 0.585 8.655 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 1.445 3.535 1.615 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 0.765 4.455 0.935 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.425 4.915 0.595 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 0.765 5.835 0.935 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 0.765 7.215 0.935 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 0.425 7.675 0.595 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
    LAYER met1 ;
      RECT 3.305 1.415 3.595 1.46 ;
      RECT 3.305 1.46 5.895 1.6 ;
      RECT 3.305 1.6 3.595 1.645 ;
      RECT 4.225 0.735 4.515 0.78 ;
      RECT 4.225 0.78 7.275 0.92 ;
      RECT 4.225 0.92 4.515 0.965 ;
      RECT 4.685 0.395 4.975 0.44 ;
      RECT 4.685 0.44 7.735 0.58 ;
      RECT 4.685 0.58 4.975 0.625 ;
      RECT 5.605 0.735 5.895 0.78 ;
      RECT 5.605 0.92 5.895 0.965 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.985 0.735 7.275 0.78 ;
      RECT 6.985 0.92 7.275 0.965 ;
      RECT 7.445 0.395 7.735 0.44 ;
      RECT 7.445 0.58 7.735 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_2
MACRO sky130_fd_sc_hd__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.34 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.937500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.71 1.78 1.325 ;
      LAYER mcon ;
        RECT 1.525 0.765 1.695 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.265 0.645 4.515 1.325 ;
      LAYER mcon ;
        RECT 4.31 0.765 4.48 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 0.735 1.755 0.78 ;
        RECT 1.465 0.78 4.54 0.92 ;
        RECT 1.465 0.92 1.755 0.965 ;
        RECT 4.25 0.735 4.54 0.78 ;
        RECT 4.25 0.92 4.54 0.965 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.53 1.075 10.975 1.275 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.61 0.755 6.935 0.925 ;
        RECT 6.61 0.925 6.88 1.675 ;
        RECT 6.71 1.675 6.88 1.785 ;
        RECT 6.765 0.595 6.935 0.755 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.463750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.255 12.335 0.825 ;
        RECT 12.01 1.785 12.335 2.465 ;
        RECT 12.135 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.61 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.42 0.085 ;
      RECT 0 2.635 12.42 2.805 ;
      RECT 0.085 0.735 0.43 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.44 1.84 ;
      RECT 0.085 1.84 1.11 2.01 ;
      RECT 0.085 2.01 0.43 2.465 ;
      RECT 0.1 0.255 0.43 0.735 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.6 2.18 0.77 2.635 ;
      RECT 0.61 0.735 1.325 0.905 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.5 ;
      RECT 0.61 1.5 1.45 1.67 ;
      RECT 0.63 0.085 0.8 0.545 ;
      RECT 0.94 2.01 1.11 2.215 ;
      RECT 0.94 2.215 2.545 2.295 ;
      RECT 0.94 2.295 3.54 2.385 ;
      RECT 0.995 0.255 3.41 0.465 ;
      RECT 0.995 0.465 1.325 0.735 ;
      RECT 1.28 1.67 1.45 1.875 ;
      RECT 1.28 1.875 2.92 2.045 ;
      RECT 1.965 0.635 2.47 1.705 ;
      RECT 2.375 2.385 3.54 2.465 ;
      RECT 2.64 0.655 3.025 0.735 ;
      RECT 2.64 0.735 3.16 0.755 ;
      RECT 2.64 0.755 3.75 0.905 ;
      RECT 2.64 1.075 2.975 1.16 ;
      RECT 2.64 1.16 3.1 1.615 ;
      RECT 3.055 0.905 3.75 0.925 ;
      RECT 3.24 0.465 3.41 0.585 ;
      RECT 3.27 0.925 3.44 2.295 ;
      RECT 3.58 0.255 4.595 0.425 ;
      RECT 3.58 0.425 3.75 0.755 ;
      RECT 3.725 1.15 4.095 1.32 ;
      RECT 3.725 1.32 3.895 2.295 ;
      RECT 3.725 2.295 5.1 2.465 ;
      RECT 3.925 0.595 4.095 1.15 ;
      RECT 4.21 1.755 4.38 2.095 ;
      RECT 4.265 0.425 4.595 0.475 ;
      RECT 4.7 1.385 5.18 1.725 ;
      RECT 4.84 0.51 5.03 0.995 ;
      RECT 4.84 0.995 5.18 1.385 ;
      RECT 4.875 1.895 6.005 2.065 ;
      RECT 4.875 2.065 5.1 2.295 ;
      RECT 5.2 0.085 5.53 0.805 ;
      RECT 5.27 2.235 5.6 2.635 ;
      RECT 5.645 1.555 6.38 1.725 ;
      RECT 5.7 0.38 5.98 0.815 ;
      RECT 5.81 0.815 5.98 1.555 ;
      RECT 5.835 2.065 6.005 2.295 ;
      RECT 5.835 2.295 7.96 2.465 ;
      RECT 6.15 0.74 6.435 1.325 ;
      RECT 6.21 1.725 6.38 1.895 ;
      RECT 6.21 1.895 6.54 1.955 ;
      RECT 6.21 1.955 7.22 2.125 ;
      RECT 6.265 0.255 7.7 0.425 ;
      RECT 6.265 0.425 6.595 0.57 ;
      RECT 7.05 1.06 7.28 1.23 ;
      RECT 7.05 1.23 7.22 1.955 ;
      RECT 7.11 0.595 7.36 0.925 ;
      RECT 7.11 0.925 7.28 1.06 ;
      RECT 7.39 1.36 7.62 1.53 ;
      RECT 7.39 1.53 7.56 2.125 ;
      RECT 7.45 1.105 7.7 1.29 ;
      RECT 7.45 1.29 7.62 1.36 ;
      RECT 7.53 0.425 7.7 1.105 ;
      RECT 7.79 1.55 8.045 1.72 ;
      RECT 7.79 1.72 7.96 2.295 ;
      RECT 7.875 0.995 8.045 1.55 ;
      RECT 7.935 0.255 9.45 0.425 ;
      RECT 7.935 0.425 8.27 0.825 ;
      RECT 8.23 1.785 8.4 2.295 ;
      RECT 8.23 2.295 9.95 2.465 ;
      RECT 8.44 0.595 8.9 0.765 ;
      RECT 8.44 0.765 8.61 1.445 ;
      RECT 8.44 1.445 8.74 1.53 ;
      RECT 8.44 1.53 8.9 1.615 ;
      RECT 8.57 1.615 8.9 2.125 ;
      RECT 8.78 0.995 9.11 1.275 ;
      RECT 9.07 1.53 9.45 2.045 ;
      RECT 9.07 2.045 9.42 2.125 ;
      RECT 9.28 0.425 9.45 1.53 ;
      RECT 9.62 2.215 9.95 2.295 ;
      RECT 9.65 0.255 10.02 0.825 ;
      RECT 9.65 0.825 9.82 1.535 ;
      RECT 9.65 1.535 9.95 2.215 ;
      RECT 9.99 0.995 10.36 1.325 ;
      RECT 10.12 2.275 10.455 2.635 ;
      RECT 10.19 0.735 10.92 0.905 ;
      RECT 10.19 0.905 10.36 0.995 ;
      RECT 10.19 1.325 10.36 1.455 ;
      RECT 10.19 1.455 10.835 2.045 ;
      RECT 10.2 0.085 10.37 0.565 ;
      RECT 10.54 0.285 10.92 0.735 ;
      RECT 10.625 2.045 10.835 2.465 ;
      RECT 11.085 1.455 11.415 2.465 ;
      RECT 11.165 0.27 11.335 0.68 ;
      RECT 11.165 0.68 11.415 1.455 ;
      RECT 11.535 0.085 11.825 0.555 ;
      RECT 11.585 1.785 11.84 2.635 ;
      RECT 11.655 0.995 11.965 1.615 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.28 1.785 1.45 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 1.105 2.155 1.275 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.21 1.785 4.38 1.955 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.77 1.445 4.94 1.615 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.15 1.105 6.32 1.275 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.53 0.765 7.7 0.935 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.45 1.445 8.62 1.615 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.91 1.105 9.08 1.275 ;
      RECT 9.28 1.785 9.45 1.955 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.19 1.785 10.36 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.23 0.765 11.4 0.935 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 11.69 1.445 11.86 1.615 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
    LAYER met1 ;
      RECT 1.195 1.755 1.51 1.8 ;
      RECT 1.195 1.8 4.44 1.94 ;
      RECT 1.195 1.94 1.51 1.985 ;
      RECT 1.925 1.075 2.215 1.12 ;
      RECT 1.925 1.12 9.14 1.26 ;
      RECT 1.925 1.26 2.215 1.305 ;
      RECT 2.845 1.415 3.16 1.46 ;
      RECT 2.845 1.46 5 1.6 ;
      RECT 2.845 1.6 3.16 1.645 ;
      RECT 4.15 1.755 4.44 1.8 ;
      RECT 4.15 1.94 4.44 1.985 ;
      RECT 4.71 1.415 5 1.46 ;
      RECT 4.71 1.6 5 1.645 ;
      RECT 6.09 1.075 6.38 1.12 ;
      RECT 6.09 1.26 6.38 1.305 ;
      RECT 7.47 0.735 7.76 0.78 ;
      RECT 7.47 0.78 11.46 0.92 ;
      RECT 7.47 0.92 7.76 0.965 ;
      RECT 8.39 1.415 8.68 1.46 ;
      RECT 8.39 1.46 11.92 1.6 ;
      RECT 8.39 1.6 8.68 1.645 ;
      RECT 8.85 1.075 9.14 1.12 ;
      RECT 8.85 1.26 9.14 1.305 ;
      RECT 9.195 1.755 9.51 1.8 ;
      RECT 9.195 1.8 10.42 1.94 ;
      RECT 9.195 1.94 9.51 1.985 ;
      RECT 10.13 1.755 10.42 1.8 ;
      RECT 10.13 1.94 10.42 1.985 ;
      RECT 11.17 0.735 11.46 0.78 ;
      RECT 11.17 0.92 11.46 0.965 ;
      RECT 11.63 1.415 11.92 1.46 ;
      RECT 11.63 1.6 11.92 1.645 ;
  END
END sky130_fd_sc_hd__fahcon_1
MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.065 4.97 1.31 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.03 1.065 3.375 1.48 ;
        RECT 3.03 1.48 6.45 1.705 ;
        RECT 5.205 1.075 6.45 1.48 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.65 1.615 ;
        RECT 0.48 0.995 0.65 1.075 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 0.37 1.465 0.615 ;
        RECT 1.275 0.615 2.325 0.695 ;
        RECT 1.275 0.695 4.885 0.865 ;
        RECT 1.56 1.585 2.86 1.705 ;
        RECT 1.56 1.705 2.725 2.035 ;
        RECT 2.135 0.255 2.325 0.615 ;
        RECT 2.57 0.865 4.885 0.895 ;
        RECT 2.57 0.895 2.86 1.585 ;
        RECT 3.255 0.675 4.885 0.695 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.09 0.255 0.445 0.615 ;
      RECT 0.09 0.615 1.105 0.795 ;
      RECT 0.125 1.785 0.99 2.005 ;
      RECT 0.125 2.005 0.455 2.465 ;
      RECT 0.625 2.175 0.885 2.635 ;
      RECT 0.72 0.085 1.105 0.445 ;
      RECT 0.82 0.795 1.105 1.035 ;
      RECT 0.82 1.035 2.4 1.345 ;
      RECT 0.82 1.345 0.99 1.785 ;
      RECT 1.16 1.795 1.355 2.215 ;
      RECT 1.16 2.215 3.095 2.465 ;
      RECT 1.635 0.085 1.965 0.445 ;
      RECT 1.935 2.205 3.095 2.215 ;
      RECT 2.495 0.085 3.085 0.525 ;
      RECT 2.895 1.875 6.605 2.105 ;
      RECT 2.895 2.105 3.095 2.205 ;
      RECT 3.265 0.255 5.315 0.505 ;
      RECT 3.265 2.275 3.595 2.635 ;
      RECT 4.125 2.275 4.455 2.635 ;
      RECT 4.625 2.105 4.815 2.465 ;
      RECT 4.985 2.275 5.315 2.635 ;
      RECT 5.055 0.505 5.315 0.735 ;
      RECT 5.055 0.735 6.175 0.905 ;
      RECT 5.485 0.085 5.675 0.565 ;
      RECT 5.485 2.105 5.665 2.465 ;
      RECT 5.845 0.255 6.175 0.735 ;
      RECT 5.845 2.275 6.175 2.635 ;
      RECT 6.345 0.085 6.605 0.885 ;
      RECT 6.345 2.105 6.605 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
  END
END sky130_fd_sc_hd__a21boi_4
MACRO sky130_fd_sc_hd__a21boi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.765 2.17 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.34 0.765 2.615 1.435 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.47 1.2 0.895 1.955 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.392200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.2 1.61 1.655 ;
        RECT 1.065 1.655 1.305 2.465 ;
        RECT 1.315 0.255 1.61 1.2 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 0.28 0.38 0.78 ;
      RECT 0.095 0.78 1.145 1.03 ;
      RECT 0.095 1.03 0.3 2.085 ;
      RECT 0.095 2.085 0.355 2.465 ;
      RECT 0.525 2.175 0.855 2.635 ;
      RECT 0.55 0.085 1.145 0.61 ;
      RECT 1.475 1.825 2.665 2.005 ;
      RECT 1.475 2.005 1.805 2.465 ;
      RECT 1.975 2.175 2.165 2.635 ;
      RECT 2.335 0.085 2.665 0.595 ;
      RECT 2.335 2.005 2.665 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__a21boi_0
MACRO sky130_fd_sc_hd__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.995 2.155 1.345 ;
        RECT 1.945 0.375 2.155 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 0.995 2.64 1.345 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.975 0.335 1.665 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.045 1.58 1.345 ;
        RECT 1.045 1.345 1.375 2.455 ;
        RECT 1.335 0.265 1.765 0.795 ;
        RECT 1.335 0.795 1.58 1.045 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 1.845 0.855 2.045 ;
      RECT 0.095 2.045 0.355 2.435 ;
      RECT 0.365 0.265 0.745 0.715 ;
      RECT 0.515 0.715 0.745 1.165 ;
      RECT 0.515 1.165 0.855 1.845 ;
      RECT 0.525 2.225 0.855 2.635 ;
      RECT 0.925 0.085 1.155 0.865 ;
      RECT 1.545 1.525 2.585 1.725 ;
      RECT 1.545 1.725 1.735 2.455 ;
      RECT 1.905 1.905 2.235 2.635 ;
      RECT 2.325 0.085 2.655 0.815 ;
      RECT 2.415 1.725 2.585 2.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__a21boi_1
MACRO sky130_fd_sc_hd__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605 0.995 3.215 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 2.425 1.245 ;
        RECT 2.1 1.245 2.425 1.495 ;
        RECT 2.1 1.495 3.675 1.675 ;
        RECT 3.385 1.035 3.795 1.295 ;
        RECT 3.385 1.295 3.675 1.495 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.765 0.425 1.805 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.255 1.72 0.615 ;
        RECT 1.52 0.615 3.06 0.785 ;
        RECT 1.52 0.785 1.715 2.115 ;
        RECT 2.73 0.255 3.06 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.095 2.08 0.425 2.635 ;
      RECT 0.265 0.36 0.795 0.53 ;
      RECT 0.595 0.53 0.795 1.07 ;
      RECT 0.595 1.07 1.325 1.285 ;
      RECT 0.595 1.285 0.855 2.265 ;
      RECT 0.985 0.085 1.225 0.885 ;
      RECT 1.045 1.795 1.35 2.285 ;
      RECT 1.045 2.285 2.215 2.465 ;
      RECT 1.885 1.855 3.92 2.025 ;
      RECT 1.885 2.025 2.215 2.285 ;
      RECT 1.94 0.085 2.27 0.445 ;
      RECT 2.385 2.195 2.555 2.635 ;
      RECT 2.81 2.025 3.92 2.105 ;
      RECT 2.81 2.105 2.98 2.465 ;
      RECT 3.16 2.275 3.49 2.635 ;
      RECT 3.635 0.085 3.93 0.865 ;
      RECT 3.66 2.105 3.92 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a21boi_2
MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s4s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.57 1.7 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.66 0.255 3.105 0.825 ;
        RECT 2.66 1.495 3.565 1.675 ;
        RECT 2.66 1.675 3.105 2.465 ;
        RECT 2.735 0.825 3.105 0.995 ;
        RECT 2.735 0.995 3.565 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.12 -0.085 0.29 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.255 0.52 0.655 ;
      RECT 0.085 0.655 1.075 0.825 ;
      RECT 0.085 1.87 1.075 2.04 ;
      RECT 0.085 2.04 0.52 2.465 ;
      RECT 0.69 0.085 1.075 0.485 ;
      RECT 0.69 2.21 1.075 2.635 ;
      RECT 0.74 0.825 1.075 0.995 ;
      RECT 0.74 0.995 1.15 1.325 ;
      RECT 0.74 1.325 1.075 1.87 ;
      RECT 1.245 0.255 1.515 0.825 ;
      RECT 1.245 1.495 1.97 1.675 ;
      RECT 1.245 1.675 1.515 2.465 ;
      RECT 1.32 0.825 1.515 0.995 ;
      RECT 1.32 0.995 1.97 1.495 ;
      RECT 1.685 0.255 1.935 0.655 ;
      RECT 1.685 0.655 2.49 0.825 ;
      RECT 1.685 1.845 2.49 2.04 ;
      RECT 1.685 2.04 1.935 2.465 ;
      RECT 2.105 0.085 2.49 0.485 ;
      RECT 2.105 2.21 2.49 2.635 ;
      RECT 2.14 0.825 2.49 0.995 ;
      RECT 2.14 0.995 2.565 1.325 ;
      RECT 2.14 1.325 2.49 1.845 ;
      RECT 3.275 0.255 3.53 0.655 ;
      RECT 3.275 0.655 4.085 0.825 ;
      RECT 3.275 1.845 4.085 2.04 ;
      RECT 3.275 2.04 3.53 2.465 ;
      RECT 3.7 0.085 4.085 0.485 ;
      RECT 3.7 2.21 4.085 2.635 ;
      RECT 3.735 0.825 4.085 0.995 ;
      RECT 3.735 0.995 4.16 1.325 ;
      RECT 3.735 1.325 4.085 1.845 ;
      RECT 4.255 0.255 4.515 0.825 ;
      RECT 4.255 1.495 4.515 2.465 ;
      RECT 4.33 0.825 4.515 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1
MACRO sky130_fd_sc_hd__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.365 2.62 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.81 0.75 3.125 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.995 1.79 1.41 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.635 0.955 0.825 ;
        RECT 0.555 0.825 0.785 2.465 ;
        RECT 0.765 0.255 0.955 0.635 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.095 1.665 0.385 2.635 ;
      RECT 0.265 0.085 0.595 0.465 ;
      RECT 0.955 0.995 1.295 1.69 ;
      RECT 0.955 1.69 1.79 1.92 ;
      RECT 0.955 2.22 1.285 2.635 ;
      RECT 1.125 0.085 1.455 0.445 ;
      RECT 1.125 0.655 1.865 0.825 ;
      RECT 1.125 0.825 1.295 0.995 ;
      RECT 1.475 1.92 1.79 2.465 ;
      RECT 1.675 0.255 1.865 0.655 ;
      RECT 1.96 1.67 3.075 1.935 ;
      RECT 1.96 1.935 2.185 2.465 ;
      RECT 2.355 2.125 2.685 2.635 ;
      RECT 2.805 0.085 3.135 0.565 ;
      RECT 2.855 1.935 3.075 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a21o_2
MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.99 1.01 4.515 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425 1.01 3.82 1.275 ;
        RECT 3.645 1.275 3.82 1.51 ;
        RECT 3.645 1.51 4.935 1.68 ;
        RECT 4.685 1.055 5.1 1.29 ;
        RECT 4.685 1.29 4.935 1.51 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.995 2.705 1.525 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.615 1.735 0.785 ;
        RECT 0.145 0.785 0.63 1.585 ;
        RECT 0.145 1.585 1.735 1.755 ;
        RECT 0.625 1.755 0.795 2.185 ;
        RECT 1.485 1.755 1.735 2.185 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.105 0.085 0.445 0.445 ;
      RECT 0.115 1.935 0.445 2.635 ;
      RECT 0.8 0.995 2.205 1.325 ;
      RECT 0.975 0.085 1.305 0.445 ;
      RECT 0.975 1.935 1.305 2.635 ;
      RECT 1.91 0.085 2.685 0.445 ;
      RECT 1.915 1.515 2.165 2.635 ;
      RECT 2.035 0.615 3.045 0.67 ;
      RECT 2.035 0.67 4.365 0.785 ;
      RECT 2.035 0.785 2.205 0.995 ;
      RECT 2.455 1.695 2.625 2.295 ;
      RECT 2.455 2.295 3.465 2.465 ;
      RECT 2.875 0.255 3.045 0.615 ;
      RECT 2.875 0.785 4.365 0.84 ;
      RECT 2.875 0.84 3.045 2.125 ;
      RECT 3.255 0.085 3.585 0.445 ;
      RECT 3.285 1.445 3.465 1.85 ;
      RECT 3.285 1.85 5.36 2.02 ;
      RECT 3.285 2.02 3.465 2.295 ;
      RECT 3.635 2.275 3.965 2.635 ;
      RECT 4.085 0.405 4.365 0.67 ;
      RECT 4.135 2.02 4.305 2.465 ;
      RECT 4.475 2.275 4.805 2.635 ;
      RECT 4.945 0.085 5.225 0.885 ;
      RECT 5.03 2.02 5.36 2.395 ;
      RECT 5.105 1.46 5.36 1.85 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__a21o_4
MACRO sky130_fd_sc_hd__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.66 1.015 2.185 1.325 ;
        RECT 1.955 0.375 2.185 1.015 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 0.995 2.665 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.015 1.48 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.355 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.525 1.905 0.865 2.635 ;
      RECT 0.545 0.635 1.775 0.835 ;
      RECT 0.545 0.835 0.835 1.505 ;
      RECT 0.545 1.505 1.315 1.725 ;
      RECT 0.615 0.085 1.285 0.455 ;
      RECT 1.045 1.725 1.315 2.455 ;
      RECT 1.465 0.265 1.775 0.635 ;
      RECT 1.495 1.505 2.655 1.745 ;
      RECT 1.495 1.745 1.725 2.455 ;
      RECT 1.895 1.925 2.225 2.635 ;
      RECT 2.365 0.085 2.655 0.815 ;
      RECT 2.395 1.745 2.655 2.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__a21o_1
MACRO sky130_fd_sc_hd__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.735 2.415 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.59 0.085 1.325 0.565 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.335 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.99 1.495 2.235 1.665 ;
      RECT 0.99 1.665 1.41 1.915 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.495 0.655 2.235 0.825 ;
      RECT 1.835 0.085 2.215 0.485 ;
      RECT 1.915 1.835 2.195 2.635 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.295 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__or2b_1
MACRO sky130_fd_sc_hd__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.63 1.075 2.32 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.955 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.29 2.655 0.735 ;
        RECT 2.325 0.735 4.055 0.905 ;
        RECT 2.365 1.785 3.455 1.955 ;
        RECT 2.365 1.955 2.615 2.465 ;
        RECT 2.83 1.445 4.055 1.615 ;
        RECT 2.83 1.615 3.455 1.785 ;
        RECT 3.165 0.29 3.495 0.735 ;
        RECT 3.205 1.955 3.455 2.465 ;
        RECT 3.67 0.905 4.055 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 2.125 0.345 2.635 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.59 0.085 1.245 0.565 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.12 1.325 ;
      RECT 0.595 1.325 0.765 2.465 ;
      RECT 0.99 1.495 2.66 1.615 ;
      RECT 0.99 1.615 1.46 2.465 ;
      RECT 1.29 0.735 1.745 0.905 ;
      RECT 1.29 0.905 1.46 1.445 ;
      RECT 1.29 1.445 2.66 1.495 ;
      RECT 1.415 0.305 1.745 0.735 ;
      RECT 1.915 1.835 2.195 2.635 ;
      RECT 1.98 0.085 2.155 0.905 ;
      RECT 2.49 1.075 3.5 1.245 ;
      RECT 2.49 1.245 2.66 1.445 ;
      RECT 2.785 2.135 3.035 2.635 ;
      RECT 2.825 0.085 2.995 0.55 ;
      RECT 3.625 1.795 3.875 2.635 ;
      RECT 3.665 0.085 3.835 0.55 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__or2b_4
MACRO sky130_fd_sc_hd__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.73 2.415 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 0.415 2.63 0.76 ;
        RECT 2.4 1.495 2.63 2.465 ;
        RECT 2.46 0.76 2.63 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 0.105 0.265 0.42 0.735 ;
      RECT 0.105 0.735 0.84 0.905 ;
      RECT 0.59 0.085 1.32 0.565 ;
      RECT 0.595 0.905 0.84 0.995 ;
      RECT 0.595 0.995 1.33 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.985 1.495 2.23 1.665 ;
      RECT 0.985 1.665 1.405 1.915 ;
      RECT 1.49 0.305 1.66 0.655 ;
      RECT 1.49 0.655 2.23 0.825 ;
      RECT 1.83 0.085 2.21 0.485 ;
      RECT 1.91 1.835 2.19 2.635 ;
      RECT 2.06 0.825 2.23 0.995 ;
      RECT 2.06 0.995 2.29 1.325 ;
      RECT 2.06 1.325 2.23 1.495 ;
      RECT 2.8 0.085 3.055 0.925 ;
      RECT 2.8 1.46 3.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__or2b_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075 5.245 0.2 5.395 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.25 1.305 7.405 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 7.36 5.525 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 7.36 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.825 0.085 6.155 0.845 ;
      RECT 5.905 1.61 6.075 2.635 ;
      RECT 6.755 0.085 7.005 0.925 ;
      RECT 6.755 1.61 6.935 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.585 5.355 6.755 5.525 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.045 5.355 7.215 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 7.36 0.24 ;
    LAYER nwell ;
      RECT -0.19 1.305 0.65 4.135 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
MACRO sky130_fd_sc_hd__dlrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.68 0.33 5.85 0.665 ;
        RECT 5.68 0.665 6.15 0.835 ;
        RECT 5.68 1.495 6.065 1.66 ;
        RECT 5.68 1.66 5.93 2.465 ;
        RECT 5.79 0.835 6.15 0.885 ;
        RECT 5.79 0.885 6.36 1.325 ;
        RECT 5.79 1.325 6.065 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515 0.255 7.765 0.825 ;
        RECT 7.515 1.605 7.765 2.465 ;
        RECT 7.595 0.825 7.765 1.055 ;
        RECT 7.595 1.055 8.195 1.325 ;
        RECT 7.595 1.325 7.765 1.605 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.4 0.995 5.15 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.745 2.255 3.585 2.425 ;
      RECT 2.77 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.905 ;
      RECT 2.925 1.905 3.125 1.995 ;
      RECT 3.27 2.125 3.585 2.255 ;
      RECT 3.305 2.075 3.585 2.125 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.395 2.015 3.605 2.045 ;
      RECT 3.395 2.045 3.585 2.075 ;
      RECT 3.415 1.99 3.605 2.015 ;
      RECT 3.42 1.975 3.605 1.99 ;
      RECT 3.43 1.96 3.605 1.975 ;
      RECT 3.435 1.165 4.2 1.325 ;
      RECT 3.435 1.325 3.605 1.96 ;
      RECT 3.74 0.085 4.07 0.53 ;
      RECT 3.755 2.135 4.6 2.635 ;
      RECT 3.84 1.535 5.51 1.705 ;
      RECT 3.84 1.705 4.94 1.865 ;
      RECT 4.27 0.415 4.57 0.655 ;
      RECT 4.27 0.655 5.51 0.825 ;
      RECT 4.77 1.865 4.94 2.435 ;
      RECT 5.11 0.085 5.49 0.485 ;
      RECT 5.11 1.875 5.49 2.635 ;
      RECT 5.32 0.825 5.51 0.995 ;
      RECT 5.32 0.995 5.62 1.325 ;
      RECT 5.32 1.325 5.51 1.535 ;
      RECT 6.02 0.085 6.36 0.465 ;
      RECT 6.1 1.83 6.36 2.635 ;
      RECT 6.535 0.255 6.865 0.995 ;
      RECT 6.535 0.995 7.425 1.325 ;
      RECT 6.535 1.325 6.87 2.465 ;
      RECT 7.035 0.085 7.34 0.545 ;
      RECT 7.045 1.835 7.34 2.635 ;
      RECT 7.935 0.085 8.195 0.885 ;
      RECT 7.935 1.495 8.195 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.785 3.1 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.16 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
  END
END sky130_fd_sc_hd__dlrbp_2
MACRO sky130_fd_sc_hd__dlrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.41 2.465 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475 0.255 7.735 0.595 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.565 0.595 7.735 1.785 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.45 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.6 0.765 3.095 1.035 ;
      RECT 2.745 2.255 3.585 2.425 ;
      RECT 2.77 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.905 ;
      RECT 2.925 1.905 3.13 1.995 ;
      RECT 3.27 2.125 3.585 2.255 ;
      RECT 3.305 2.075 3.585 2.125 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.395 2.015 3.605 2.045 ;
      RECT 3.395 2.045 3.585 2.075 ;
      RECT 3.415 1.99 3.605 2.015 ;
      RECT 3.42 1.975 3.605 1.99 ;
      RECT 3.43 1.96 3.605 1.975 ;
      RECT 3.435 1.165 4.2 1.325 ;
      RECT 3.435 1.325 3.605 1.96 ;
      RECT 3.735 0.085 4.07 0.53 ;
      RECT 3.755 2.135 4.59 2.635 ;
      RECT 3.84 1.535 5.89 1.765 ;
      RECT 3.84 1.765 4.95 1.865 ;
      RECT 4.24 0.255 4.54 0.655 ;
      RECT 4.24 0.655 5.89 0.825 ;
      RECT 4.78 1.865 4.95 2.435 ;
      RECT 5.12 0.085 5.89 0.485 ;
      RECT 5.12 1.935 5.89 2.635 ;
      RECT 5.655 0.825 5.89 1.535 ;
      RECT 6.58 0.255 6.805 0.995 ;
      RECT 6.58 0.995 7.395 1.325 ;
      RECT 6.58 1.325 6.83 2.465 ;
      RECT 6.975 0.085 7.305 0.465 ;
      RECT 7.01 1.835 7.305 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.925 1.785 3.095 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.155 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrbp_1
MACRO sky130_fd_sc_hd__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.995 2.325 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.995 1.82 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.88 0.995 1.24 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.36 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.72 0.255 3.05 0.615 ;
        RECT 2.72 0.615 3.54 0.785 ;
        RECT 2.81 1.905 3.54 2.075 ;
        RECT 2.81 2.075 3 2.465 ;
        RECT 3.345 0.785 3.54 1.905 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 1.51 2.665 1.765 ;
      RECT 0.09 1.765 0.355 2.465 ;
      RECT 0.095 0.255 0.43 0.425 ;
      RECT 0.095 0.425 0.71 0.825 ;
      RECT 0.525 1.935 0.855 2.635 ;
      RECT 0.53 0.825 0.71 1.51 ;
      RECT 0.88 0.635 2.15 0.825 ;
      RECT 1.025 1.765 1.695 2.465 ;
      RECT 1.39 0.085 1.725 0.465 ;
      RECT 2.2 1.935 2.63 2.635 ;
      RECT 2.315 0.085 2.55 0.525 ;
      RECT 2.495 0.995 3.175 1.325 ;
      RECT 2.495 1.325 2.665 1.51 ;
      RECT 3.17 2.255 3.5 2.635 ;
      RECT 3.22 0.085 3.55 0.445 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o211a_2
MACRO sky130_fd_sc_hd__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 1.075 1.72 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 1.075 2.22 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 1.075 2.72 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245 1.075 3.595 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.885 ;
        RECT 0.085 0.885 0.26 1.495 ;
        RECT 0.085 1.495 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.43 1.075 1.125 1.245 ;
      RECT 0.595 0.085 0.845 0.885 ;
      RECT 0.595 1.495 0.765 2.635 ;
      RECT 0.955 1.245 1.125 1.495 ;
      RECT 0.955 1.495 3.39 1.665 ;
      RECT 1.035 0.255 1.365 0.735 ;
      RECT 1.035 0.735 2.26 0.905 ;
      RECT 1.035 1.835 1.285 2.635 ;
      RECT 1.535 0.085 1.76 0.545 ;
      RECT 1.93 0.255 2.26 0.735 ;
      RECT 1.93 1.665 2.26 2.465 ;
      RECT 2.56 1.835 2.89 2.635 ;
      RECT 2.89 0.255 3.39 0.865 ;
      RECT 2.89 0.865 3.06 1.495 ;
      RECT 3.06 1.665 3.39 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o211a_1
MACRO sky130_fd_sc_hd__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.49 1.035 4.845 1.495 ;
        RECT 4.49 1.495 6.29 1.685 ;
        RECT 5.89 1.035 6.29 1.495 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.03 1.035 5.705 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.995 2.83 1.445 ;
        RECT 2.54 1.445 4.28 1.685 ;
        RECT 3.95 1.035 4.28 1.445 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.055 1.035 3.74 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.911000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 1.605 0.805 ;
        RECT 0.085 0.805 0.365 1.435 ;
        RECT 0.085 1.435 2.03 1.7 ;
        RECT 0.595 0.255 0.765 0.615 ;
        RECT 0.595 0.615 1.605 0.635 ;
        RECT 0.98 1.7 1.16 2.465 ;
        RECT 1.435 0.255 1.605 0.615 ;
        RECT 1.84 1.7 2.03 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 0.48 1.87 0.81 2.635 ;
      RECT 0.535 1.065 2.37 1.265 ;
      RECT 0.935 0.085 1.265 0.445 ;
      RECT 1.34 1.87 1.67 2.635 ;
      RECT 1.775 0.085 2.14 0.465 ;
      RECT 2.2 0.635 3.52 0.815 ;
      RECT 2.2 0.815 2.37 1.065 ;
      RECT 2.2 1.265 2.37 1.855 ;
      RECT 2.2 1.855 5.485 2.025 ;
      RECT 2.2 2.2 2.53 2.635 ;
      RECT 2.33 0.255 4.5 0.465 ;
      RECT 2.7 2.025 3.06 2.465 ;
      RECT 3.285 2.195 3.615 2.635 ;
      RECT 3.785 2.025 4.12 2.465 ;
      RECT 4.17 0.465 4.5 0.695 ;
      RECT 4.17 0.695 6.345 0.865 ;
      RECT 4.29 2.195 4.555 2.635 ;
      RECT 4.67 0.085 4.985 0.525 ;
      RECT 5.155 0.255 5.485 0.695 ;
      RECT 5.155 2.025 5.485 2.465 ;
      RECT 5.655 0.085 5.845 0.525 ;
      RECT 6.015 0.255 6.345 0.695 ;
      RECT 6.015 1.915 6.345 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__o211a_4
MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.51 1.56 12.78 2.465 ;
        RECT 12.52 0.255 12.78 0.76 ;
        RECT 12.6 0.76 12.78 1.56 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 13.07 2.91 ;
        RECT 4.405 1.305 13.07 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.88 0.085 ;
      RECT 0 2.635 12.88 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.72 0.085 10.89 0.545 ;
      RECT 10.72 1.495 10.97 2.635 ;
      RECT 11.65 1.535 12.325 1.705 ;
      RECT 11.65 1.705 11.83 2.465 ;
      RECT 11.66 0.255 11.83 0.635 ;
      RECT 11.66 0.635 12.325 0.805 ;
      RECT 12.01 0.085 12.34 0.465 ;
      RECT 12.01 1.875 12.34 2.635 ;
      RECT 12.155 0.805 12.325 1.06 ;
      RECT 12.155 1.06 12.43 1.39 ;
      RECT 12.155 1.39 12.325 1.535 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrbp_1
MACRO sky130_fd_sc_hd__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.575 0.265 11.925 1.695 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.435 1.535 12.825 2.08 ;
        RECT 12.445 0.31 12.825 0.825 ;
        RECT 12.525 2.08 12.825 2.465 ;
        RECT 12.655 0.825 12.825 1.535 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 13.53 2.91 ;
        RECT 4.405 1.305 13.53 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 13.34 0.085 ;
      RECT 0 2.635 13.34 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 1.055 ;
      RECT 10.345 1.055 11.06 1.295 ;
      RECT 10.375 1.295 11.06 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.715 0.345 10.885 0.715 ;
      RECT 10.715 0.715 11.405 0.885 ;
      RECT 10.715 1.795 11.405 1.865 ;
      RECT 10.715 1.865 12.265 2.035 ;
      RECT 10.715 2.035 10.89 2.465 ;
      RECT 11.09 0.085 11.365 0.545 ;
      RECT 11.09 2.205 11.42 2.635 ;
      RECT 11.23 0.885 11.405 1.795 ;
      RECT 11.55 2.035 12.265 2.085 ;
      RECT 12.025 2.255 12.355 2.635 ;
      RECT 12.095 0.995 12.485 1.325 ;
      RECT 12.095 1.325 12.265 1.865 ;
      RECT 12.105 0.085 12.275 0.825 ;
      RECT 12.995 0.085 13.165 0.93 ;
      RECT 12.995 1.495 13.245 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrbp_2
MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.625 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.57 0.255 3.135 0.825 ;
        RECT 2.57 1.495 3.135 2.465 ;
        RECT 2.675 0.825 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.255 0.485 0.715 ;
      RECT 0.085 0.715 1.03 0.885 ;
      RECT 0.085 1.785 1.03 2.005 ;
      RECT 0.085 2.005 0.485 2.465 ;
      RECT 0.655 0.085 0.925 0.545 ;
      RECT 0.655 2.175 0.925 2.635 ;
      RECT 0.795 0.885 1.03 0.995 ;
      RECT 0.795 0.995 1.085 1.325 ;
      RECT 0.795 1.325 1.03 1.785 ;
      RECT 1.155 0.255 1.425 0.585 ;
      RECT 1.155 2.135 1.425 2.465 ;
      RECT 1.255 0.585 1.425 1.055 ;
      RECT 1.255 1.055 2.03 1.615 ;
      RECT 1.255 1.615 1.425 2.135 ;
      RECT 1.615 0.255 1.875 0.715 ;
      RECT 1.615 0.715 2.4 0.885 ;
      RECT 1.615 1.785 2.4 2.005 ;
      RECT 1.615 2.005 1.875 2.465 ;
      RECT 2.075 0.085 2.4 0.545 ;
      RECT 2.075 2.175 2.4 2.635 ;
      RECT 2.2 0.885 2.4 0.995 ;
      RECT 2.2 0.995 2.505 1.325 ;
      RECT 2.2 1.325 2.4 1.785 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1
MACRO sky130_fd_sc_hd__a221o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.675 2.255 1.075 ;
        RECT 1.97 1.075 2.3 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.275 ;
        RECT 1.42 0.675 1.7 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.255 3.575 0.585 ;
        RECT 3.32 1.795 3.575 2.465 ;
        RECT 3.39 0.585 3.575 0.665 ;
        RECT 3.405 0.665 3.575 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.24 0.905 ;
      RECT 0.175 1.455 3.235 1.625 ;
      RECT 0.175 1.625 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.515 1.795 0.845 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.65 2.035 ;
      RECT 1.015 2.035 1.245 2.125 ;
      RECT 1.07 0.255 2.605 0.505 ;
      RECT 1.07 0.505 1.24 0.735 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 1.875 2.215 2.23 2.635 ;
      RECT 2.4 2.035 2.65 2.465 ;
      RECT 2.435 0.505 2.605 0.735 ;
      RECT 2.435 0.735 3.235 0.905 ;
      RECT 2.775 0.085 3.105 0.565 ;
      RECT 2.82 1.875 3.15 2.635 ;
      RECT 3.065 0.905 3.235 1.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a221o_1
MACRO sky130_fd_sc_hd__a221o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.675 2.255 1.075 ;
        RECT 1.97 1.075 2.3 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.275 ;
        RECT 1.42 0.675 1.7 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.44 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.255 3.575 0.585 ;
        RECT 3.32 1.795 3.575 2.465 ;
        RECT 3.39 0.585 3.575 0.665 ;
        RECT 3.405 0.665 3.575 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.24 0.905 ;
      RECT 0.175 1.455 3.235 1.625 ;
      RECT 0.175 1.625 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.515 1.795 0.845 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.65 2.035 ;
      RECT 1.015 2.035 1.245 2.125 ;
      RECT 1.07 0.255 2.605 0.505 ;
      RECT 1.07 0.505 1.24 0.735 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 1.875 2.215 2.23 2.635 ;
      RECT 2.4 2.035 2.65 2.465 ;
      RECT 2.435 0.505 2.605 0.735 ;
      RECT 2.435 0.735 3.235 0.905 ;
      RECT 2.775 0.085 3.105 0.565 ;
      RECT 2.82 1.875 3.15 2.635 ;
      RECT 3.065 0.905 3.235 1.455 ;
      RECT 3.745 0.085 3.915 0.98 ;
      RECT 3.745 1.445 3.915 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a221o_2
MACRO sky130_fd_sc_hd__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.075 3.19 1.105 ;
        RECT 2.855 1.105 4.06 1.285 ;
        RECT 3.71 1.075 4.06 1.105 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.075 2.68 1.285 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 1.075 6.035 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.27 1.075 7.28 1.285 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.23 1.075 4.725 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.735 1.685 0.905 ;
        RECT 0.095 0.905 0.325 1.455 ;
        RECT 0.095 1.455 1.645 1.625 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 1.685 0.735 ;
        RECT 0.555 1.625 0.805 2.465 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 1.395 1.625 1.645 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.085 0.325 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.155 1.795 0.385 2.635 ;
      RECT 0.175 0.085 0.345 0.555 ;
      RECT 0.495 1.075 1.845 1.115 ;
      RECT 0.495 1.115 1.985 1.285 ;
      RECT 0.975 1.795 1.225 2.635 ;
      RECT 1.015 0.085 1.185 0.555 ;
      RECT 1.815 1.285 1.985 1.455 ;
      RECT 1.815 1.455 5.065 1.625 ;
      RECT 1.815 1.795 2.065 2.635 ;
      RECT 1.855 0.085 2.025 0.555 ;
      RECT 1.855 0.735 2.525 0.905 ;
      RECT 1.945 0.905 2.165 0.935 ;
      RECT 2.195 0.255 2.525 0.735 ;
      RECT 2.235 1.795 4.23 1.875 ;
      RECT 2.235 1.875 5.575 1.965 ;
      RECT 2.235 1.965 2.485 2.465 ;
      RECT 2.655 2.135 2.905 2.635 ;
      RECT 2.695 0.085 2.865 0.895 ;
      RECT 3.075 1.965 3.33 2.465 ;
      RECT 3.08 0.305 4.305 0.475 ;
      RECT 3.19 0.735 3.885 0.905 ;
      RECT 3.315 0.905 3.61 0.935 ;
      RECT 3.5 2.135 3.75 2.635 ;
      RECT 3.55 0.645 3.885 0.735 ;
      RECT 3.94 2.215 6.385 2.295 ;
      RECT 3.94 2.295 7.225 2.465 ;
      RECT 4.055 0.475 4.305 0.725 ;
      RECT 4.055 0.725 5.065 0.905 ;
      RECT 4.06 1.965 5.575 2.045 ;
      RECT 4.405 1.625 4.735 1.705 ;
      RECT 4.475 0.085 4.645 0.555 ;
      RECT 4.815 0.255 5.985 0.475 ;
      RECT 4.815 0.475 5.065 0.725 ;
      RECT 4.895 0.905 5.065 1.455 ;
      RECT 5.235 0.645 6.505 0.725 ;
      RECT 5.235 0.725 7.345 0.905 ;
      RECT 5.245 1.455 6.805 1.625 ;
      RECT 5.245 1.625 5.575 1.875 ;
      RECT 5.745 1.795 6.385 2.215 ;
      RECT 6.555 1.625 6.805 2.125 ;
      RECT 6.675 0.085 6.845 0.555 ;
      RECT 6.975 1.785 7.225 2.295 ;
      RECT 7.015 0.255 7.345 0.725 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.995 0.765 2.165 0.935 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.4 0.765 3.57 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 1.935 0.735 2.225 0.78 ;
      RECT 1.935 0.78 3.63 0.92 ;
      RECT 1.935 0.92 2.225 0.965 ;
      RECT 3.34 0.735 3.63 0.78 ;
      RECT 3.34 0.92 3.63 0.965 ;
  END
END sky130_fd_sc_hd__a221o_4
MACRO sky130_fd_sc_hd__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probe_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.25 0.56 4.27 2.16 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.595 1.835 0.765 2.635 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.355 0.085 1.685 0.565 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
      RECT 1.435 1.835 1.605 2.635 ;
      RECT 1.855 0.255 2.025 0.735 ;
      RECT 1.855 0.735 4.545 0.905 ;
      RECT 1.855 1.445 4.545 1.615 ;
      RECT 1.855 1.615 2.025 2.465 ;
      RECT 2.195 0.085 2.525 0.565 ;
      RECT 2.195 1.835 2.525 2.635 ;
      RECT 2.695 0.255 2.865 0.735 ;
      RECT 2.695 1.615 2.865 2.465 ;
      RECT 3.035 0.085 3.365 0.565 ;
      RECT 3.035 1.835 3.365 2.635 ;
      RECT 3.535 0.255 3.705 0.735 ;
      RECT 3.535 1.615 3.705 2.465 ;
      RECT 3.875 0.085 4.205 0.565 ;
      RECT 3.875 1.835 4.205 2.635 ;
      RECT 4.29 0.905 4.545 1.055 ;
      RECT 4.29 1.055 4.885 1.315 ;
      RECT 4.29 1.315 4.545 1.445 ;
      RECT 4.375 0.255 4.545 0.735 ;
      RECT 4.375 1.615 4.545 2.465 ;
      RECT 4.715 0.085 5.045 0.885 ;
      RECT 4.715 1.485 5.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.32 1.105 4.49 1.275 ;
      RECT 4.68 1.105 4.85 1.275 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
    LAYER met1 ;
      RECT 3.465 1.06 4.105 1.075 ;
      RECT 3.465 1.075 4.91 1.305 ;
      RECT 3.465 1.305 4.105 1.32 ;
    LAYER met2 ;
      RECT 3.445 1.005 4.125 1.375 ;
    LAYER met3 ;
      RECT 3.395 1.025 4.175 1.355 ;
    LAYER met4 ;
      RECT 1.37 0.68 4.15 1.86 ;
    LAYER via ;
      RECT 3.495 1.06 3.755 1.32 ;
      RECT 3.815 1.06 4.075 1.32 ;
    LAYER via2 ;
      RECT 3.445 1.05 3.725 1.33 ;
      RECT 3.845 1.05 4.125 1.33 ;
    LAYER via3 ;
      RECT 3.425 1.03 3.745 1.35 ;
      RECT 3.825 1.03 4.145 1.35 ;
    LAYER via4 ;
      RECT 2.97 0.68 4.15 1.86 ;
  END
END sky130_fd_sc_hd__probe_p_8
MACRO sky130_fd_sc_hd__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.675 1.72 1.075 ;
        RECT 1.51 1.075 1.84 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 2.415 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.285 ;
        RECT 1.02 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.575 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.255 3.16 0.585 ;
        RECT 2.9 1.785 3.16 2.465 ;
        RECT 2.99 0.585 3.16 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.095 0.085 0.545 0.85 ;
      RECT 0.095 1.455 2.815 1.625 ;
      RECT 0.095 1.625 0.425 2.295 ;
      RECT 0.095 2.295 1.265 2.465 ;
      RECT 0.595 1.795 2.23 2.035 ;
      RECT 0.595 2.035 0.825 2.125 ;
      RECT 0.82 0.255 2.145 0.505 ;
      RECT 0.935 2.255 1.265 2.295 ;
      RECT 1.455 2.215 1.81 2.635 ;
      RECT 1.975 0.505 2.145 0.735 ;
      RECT 1.975 0.735 2.815 0.905 ;
      RECT 1.98 2.035 2.23 2.465 ;
      RECT 2.355 0.085 2.685 0.565 ;
      RECT 2.4 1.875 2.73 2.635 ;
      RECT 2.645 0.905 2.815 1.455 ;
      RECT 3.33 0.085 3.5 0.985 ;
      RECT 3.33 1.445 3.5 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a22o_2
MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.9 1.075 5.395 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.35 1.075 4.68 1.445 ;
        RECT 4.35 1.445 5.735 1.615 ;
        RECT 5.565 1.075 6.355 1.275 ;
        RECT 5.565 1.275 5.735 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.68 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.42 1.075 2.955 1.445 ;
        RECT 2.42 1.445 4.18 1.615 ;
        RECT 3.85 1.075 4.18 1.445 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.725 1.77 0.905 ;
        RECT 0.085 0.905 0.37 1.445 ;
        RECT 0.085 1.445 1.73 1.615 ;
        RECT 0.6 0.265 0.93 0.725 ;
        RECT 0.64 1.615 0.89 2.465 ;
        RECT 1.44 0.255 1.77 0.725 ;
        RECT 1.48 1.615 1.73 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.22 1.825 0.47 2.635 ;
      RECT 0.26 0.085 0.43 0.555 ;
      RECT 0.54 1.075 2.23 1.275 ;
      RECT 1.06 1.795 1.31 2.635 ;
      RECT 1.1 0.085 1.27 0.555 ;
      RECT 1.9 1.275 2.23 1.785 ;
      RECT 1.9 1.785 3.93 1.955 ;
      RECT 1.9 2.125 2.15 2.635 ;
      RECT 1.94 0.085 2.63 0.555 ;
      RECT 1.94 0.735 5.31 0.905 ;
      RECT 1.94 0.905 2.23 1.075 ;
      RECT 2.42 2.125 2.67 2.295 ;
      RECT 2.42 2.295 4.43 2.465 ;
      RECT 2.8 0.255 3.97 0.475 ;
      RECT 2.84 1.955 3.09 2.125 ;
      RECT 3.17 0.645 3.605 0.735 ;
      RECT 3.26 2.125 3.51 2.295 ;
      RECT 3.68 1.955 3.93 2.125 ;
      RECT 4.1 1.785 6.11 1.955 ;
      RECT 4.1 1.955 4.43 2.295 ;
      RECT 4.185 0.085 4.355 0.555 ;
      RECT 4.56 0.255 5.73 0.475 ;
      RECT 4.6 2.125 4.85 2.635 ;
      RECT 4.935 0.645 5.31 0.735 ;
      RECT 5.02 1.955 5.27 2.465 ;
      RECT 5.44 2.125 5.69 2.635 ;
      RECT 5.48 0.475 5.73 0.895 ;
      RECT 5.9 0.085 6.07 0.895 ;
      RECT 5.905 1.455 6.11 1.785 ;
      RECT 5.905 1.955 6.11 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__a22o_4
MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.675 1.695 1.075 ;
        RECT 1.485 1.075 1.815 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.04 2.395 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.285 ;
        RECT 1.02 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 0.255 3.135 0.585 ;
        RECT 2.875 1.785 3.135 2.465 ;
        RECT 2.965 0.585 3.135 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 0.085 0.545 0.85 ;
      RECT 0.09 1.455 1.265 1.515 ;
      RECT 0.09 1.515 2.795 1.625 ;
      RECT 0.09 1.625 0.345 2.245 ;
      RECT 0.09 2.245 0.425 2.465 ;
      RECT 0.595 1.795 0.78 1.885 ;
      RECT 0.595 1.885 2.205 2.085 ;
      RECT 0.595 2.085 0.825 2.125 ;
      RECT 0.82 0.255 2.12 0.465 ;
      RECT 0.935 1.625 2.735 1.685 ;
      RECT 0.935 1.685 1.265 1.715 ;
      RECT 1.37 1.875 2.205 1.885 ;
      RECT 1.43 2.255 1.785 2.635 ;
      RECT 1.95 0.465 2.12 0.615 ;
      RECT 1.95 0.615 2.705 0.74 ;
      RECT 1.95 0.74 2.795 0.785 ;
      RECT 1.955 2.085 2.205 2.465 ;
      RECT 2.375 0.085 2.705 0.445 ;
      RECT 2.455 1.855 2.705 2.635 ;
      RECT 2.525 0.785 2.795 0.905 ;
      RECT 2.595 1.48 2.795 1.515 ;
      RECT 2.625 0.905 2.795 1.48 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a22o_1
MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvpwrvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvpwrvgnd_1
MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fah_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.44 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 2.495 1.275 ;
        RECT 1.99 1.275 2.19 1.41 ;
        RECT 2.015 1.41 2.19 1.725 ;
      LAYER mcon ;
        RECT 1.99 1.105 2.16 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.675 0.995 5.925 1.325 ;
      LAYER mcon ;
        RECT 5.68 1.105 5.85 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.93 1.075 2.22 1.12 ;
        RECT 1.93 1.12 5.91 1.26 ;
        RECT 1.93 1.26 2.22 1.305 ;
        RECT 5.62 1.075 5.91 1.12 ;
        RECT 5.62 1.26 5.91 1.305 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.475 1.075 9.865 1.325 ;
        RECT 9.69 0.735 10.01 0.935 ;
        RECT 9.69 0.935 9.865 1.075 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.87 0.27 11.31 0.825 ;
        RECT 10.87 0.825 11.04 1.495 ;
        RECT 10.87 1.495 11.39 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.506000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.98 0.255 12.335 0.825 ;
        RECT 11.985 1.785 12.335 2.465 ;
        RECT 12.11 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.61 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.42 0.085 ;
      RECT 0 2.635 12.42 2.805 ;
      RECT 0.085 0.255 0.425 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.445 1.895 ;
      RECT 0.085 1.895 2.805 2.065 ;
      RECT 0.085 2.065 0.395 2.465 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.565 2.26 0.93 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.595 0.735 1.32 0.905 ;
      RECT 0.595 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.38 ;
      RECT 0.61 1.38 0.815 1.445 ;
      RECT 0.61 1.445 1.315 1.455 ;
      RECT 0.615 1.455 1.315 1.615 ;
      RECT 0.985 1.615 1.315 1.715 ;
      RECT 0.99 0.255 1.32 0.735 ;
      RECT 1.49 1.445 1.82 1.5 ;
      RECT 1.49 1.5 1.84 1.725 ;
      RECT 1.5 0.255 1.84 0.715 ;
      RECT 1.5 0.715 2.52 0.885 ;
      RECT 1.5 0.885 1.82 0.905 ;
      RECT 1.615 0.905 1.82 1.445 ;
      RECT 2.01 0.085 2.18 0.545 ;
      RECT 2.065 2.235 2.395 2.635 ;
      RECT 2.35 0.255 4.84 0.425 ;
      RECT 2.35 0.425 2.52 0.715 ;
      RECT 2.36 1.445 2.86 1.715 ;
      RECT 2.635 2.065 2.805 2.295 ;
      RECT 2.635 2.295 4.95 2.465 ;
      RECT 2.69 0.595 2.86 1.445 ;
      RECT 3.03 0.425 4.84 0.465 ;
      RECT 3.03 0.465 3.2 1.955 ;
      RECT 3.03 1.955 4.32 2.125 ;
      RECT 3.37 0.635 3.9 0.805 ;
      RECT 3.37 0.805 3.54 1.455 ;
      RECT 3.37 1.455 3.815 1.785 ;
      RECT 3.985 1.785 4.32 1.955 ;
      RECT 4.07 0.645 4.4 0.735 ;
      RECT 4.07 0.735 4.56 0.755 ;
      RECT 4.07 0.755 5.17 0.78 ;
      RECT 4.07 0.78 5.155 0.805 ;
      RECT 4.07 0.805 5.145 0.905 ;
      RECT 4.07 1.075 4.4 1.16 ;
      RECT 4.07 1.16 4.535 1.615 ;
      RECT 4.48 0.905 5.145 0.925 ;
      RECT 4.65 0.465 4.84 0.585 ;
      RECT 4.705 0.925 4.875 2.295 ;
      RECT 4.925 0.735 5.18 0.74 ;
      RECT 4.925 0.74 5.17 0.755 ;
      RECT 4.95 0.715 5.18 0.735 ;
      RECT 4.98 0.69 5.18 0.715 ;
      RECT 5 0.655 5.18 0.69 ;
      RECT 5.01 0.255 6.1 0.425 ;
      RECT 5.01 0.425 5.18 0.655 ;
      RECT 5.125 1.15 5.505 1.32 ;
      RECT 5.125 1.32 5.295 2.295 ;
      RECT 5.125 2.295 7.56 2.465 ;
      RECT 5.32 0.865 5.52 0.925 ;
      RECT 5.32 0.925 5.505 1.15 ;
      RECT 5.335 0.84 5.52 0.865 ;
      RECT 5.35 0.595 5.52 0.84 ;
      RECT 5.475 1.7 5.875 2.03 ;
      RECT 5.75 0.425 6.1 0.565 ;
      RECT 6.105 0.74 6.435 1.275 ;
      RECT 6.105 1.445 6.46 1.615 ;
      RECT 6.27 0.255 9.735 0.425 ;
      RECT 6.27 0.425 6.6 0.57 ;
      RECT 6.29 1.615 6.46 1.955 ;
      RECT 6.29 1.955 7.22 2.125 ;
      RECT 6.61 0.755 6.94 0.925 ;
      RECT 6.61 0.925 6.88 1.275 ;
      RECT 6.71 1.275 6.88 1.785 ;
      RECT 6.77 0.595 6.94 0.755 ;
      RECT 7.05 1.06 7.28 1.13 ;
      RECT 7.05 1.13 7.245 1.175 ;
      RECT 7.05 1.175 7.22 1.955 ;
      RECT 7.065 1.045 7.28 1.06 ;
      RECT 7.09 1.01 7.28 1.045 ;
      RECT 7.11 0.595 7.445 0.765 ;
      RECT 7.11 0.765 7.28 1.01 ;
      RECT 7.39 1.275 7.62 1.375 ;
      RECT 7.39 1.375 7.595 1.4 ;
      RECT 7.39 1.4 7.575 1.425 ;
      RECT 7.39 1.425 7.56 2.295 ;
      RECT 7.45 0.995 7.62 1.275 ;
      RECT 7.705 0.425 7.96 0.825 ;
      RECT 7.73 1.51 7.96 2.295 ;
      RECT 7.73 2.295 9.655 2.465 ;
      RECT 7.79 0.825 7.96 1.51 ;
      RECT 8.145 1.955 9.25 2.125 ;
      RECT 8.155 0.595 8.405 0.925 ;
      RECT 8.225 0.925 8.405 1.445 ;
      RECT 8.225 1.445 8.91 1.785 ;
      RECT 8.575 0.595 8.745 1.105 ;
      RECT 8.575 1.105 9.25 1.275 ;
      RECT 8.92 0.685 9.3 0.935 ;
      RECT 9.08 1.275 9.25 1.955 ;
      RECT 9.4 0.425 9.735 0.515 ;
      RECT 9.42 1.495 10.35 1.705 ;
      RECT 9.42 1.705 9.655 2.295 ;
      RECT 9.84 2.275 10.175 2.635 ;
      RECT 9.905 0.085 10.075 0.565 ;
      RECT 10.18 0.995 10.35 1.495 ;
      RECT 10.245 0.285 10.69 0.825 ;
      RECT 10.345 1.875 10.69 2.465 ;
      RECT 10.52 0.825 10.69 1.875 ;
      RECT 11.21 0.995 11.46 1.325 ;
      RECT 11.48 0.085 11.81 0.825 ;
      RECT 11.56 1.785 11.815 2.635 ;
      RECT 11.63 0.995 11.94 1.615 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.37 0.765 3.54 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.365 1.445 4.535 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.57 1.785 5.74 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.15 0.765 6.32 0.935 ;
      RECT 6.15 1.445 6.32 1.615 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.61 1.105 6.78 1.275 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.46 1.445 8.63 1.615 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.92 0.765 9.09 0.935 ;
      RECT 9.08 1.785 9.25 1.955 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.785 10.69 1.955 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.22 1.105 11.39 1.275 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 11.68 1.445 11.85 1.615 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
    LAYER met1 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.46 6.38 1.6 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 3.31 0.735 3.6 0.78 ;
      RECT 3.31 0.78 9.15 0.92 ;
      RECT 3.31 0.92 3.6 0.965 ;
      RECT 3.925 1.755 4.215 1.8 ;
      RECT 3.925 1.8 5.8 1.94 ;
      RECT 3.925 1.94 4.215 1.985 ;
      RECT 4.305 1.415 4.595 1.46 ;
      RECT 4.305 1.6 4.595 1.645 ;
      RECT 5.51 1.755 5.8 1.8 ;
      RECT 5.51 1.94 5.8 1.985 ;
      RECT 6.09 0.735 6.38 0.78 ;
      RECT 6.09 0.92 6.38 0.965 ;
      RECT 6.09 1.415 6.38 1.46 ;
      RECT 6.09 1.6 6.38 1.645 ;
      RECT 6.55 1.075 6.84 1.12 ;
      RECT 6.55 1.12 11.45 1.26 ;
      RECT 6.55 1.26 6.84 1.305 ;
      RECT 8.4 1.415 8.69 1.46 ;
      RECT 8.4 1.46 11.91 1.6 ;
      RECT 8.4 1.6 8.69 1.645 ;
      RECT 8.86 0.735 9.15 0.78 ;
      RECT 8.86 0.92 9.15 0.965 ;
      RECT 9.02 1.755 9.31 1.8 ;
      RECT 9.02 1.8 10.75 1.94 ;
      RECT 9.02 1.94 9.31 1.985 ;
      RECT 10.46 1.755 10.75 1.8 ;
      RECT 10.46 1.94 10.75 1.985 ;
      RECT 11.16 1.075 11.45 1.12 ;
      RECT 11.16 1.26 11.45 1.305 ;
      RECT 11.62 1.415 11.91 1.46 ;
      RECT 11.62 1.6 11.91 1.645 ;
  END
END sky130_fd_sc_hd__fah_1
MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.755 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.24 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 0.745 0.33 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.699000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 1.745 0.595 ;
        RECT 0.515 0.595 0.695 1.495 ;
        RECT 0.515 1.495 1.745 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.415 0.595 1.745 0.825 ;
        RECT 1.415 1.665 1.745 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.09 0.085 0.345 0.575 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 1.015 1.835 1.245 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__nand3_1
MACRO sky130_fd_sc_hd__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.33 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 2.16 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 3.595 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 0.845 1.445 ;
        RECT 0.515 1.445 3.045 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.715 1.665 3.045 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 0.295 2.105 0.465 ;
      RECT 0.09 0.465 0.345 0.785 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.355 0.635 3.045 0.905 ;
      RECT 1.855 1.835 2.545 2.635 ;
      RECT 2.295 0.085 2.625 0.465 ;
      RECT 3.215 0.085 3.595 0.885 ;
      RECT 3.215 1.445 3.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__nand3_2
MACRO sky130_fd_sc_hd__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.85 1.075 5.565 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.54 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.7 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 6.355 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 0.655 6.355 0.905 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 6.125 0.905 6.355 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 3.785 0.905 ;
      RECT 0.09 1.445 0.345 2.635 ;
      RECT 0.595 0.085 0.765 0.565 ;
      RECT 0.935 0.255 1.265 0.735 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.435 0.085 1.605 0.565 ;
      RECT 1.775 0.655 2.105 0.735 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.195 0.255 6 0.485 ;
      RECT 2.615 0.655 2.945 0.735 ;
      RECT 2.695 1.835 2.865 2.635 ;
      RECT 3.455 0.655 3.785 0.735 ;
      RECT 3.535 1.835 4.225 2.635 ;
      RECT 4.895 1.835 5.065 2.635 ;
      RECT 5.735 1.835 6 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__nand3_4
MACRO sky130_fd_sc_hd__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.995 2.06 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.995 1.305 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.995 2.675 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.125 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.265 0.425 1.685 ;
        RECT 0.09 1.685 0.355 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135 -0.085 0.305 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.525 1.915 0.855 2.635 ;
      RECT 0.6 0.625 3.085 0.815 ;
      RECT 0.6 0.815 0.825 1.505 ;
      RECT 0.6 1.505 3.095 1.685 ;
      RECT 0.605 0.085 1.35 0.455 ;
      RECT 1.045 1.865 2.235 2.095 ;
      RECT 1.045 2.095 1.305 2.455 ;
      RECT 1.475 2.265 1.805 2.635 ;
      RECT 1.915 0.265 2.17 0.625 ;
      RECT 1.975 2.095 2.235 2.455 ;
      RECT 2.35 0.085 2.68 0.455 ;
      RECT 2.805 1.685 3.095 2.455 ;
      RECT 2.86 0.265 3.085 0.625 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a211o_1
MACRO sky130_fd_sc_hd__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.035 1.02 5.38 1.33 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.495 1.02 4.825 1.51 ;
        RECT 4.495 1.51 5.845 1.7 ;
        RECT 5.635 1.02 6.225 1.32 ;
        RECT 5.635 1.32 5.845 1.51 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.985 2.805 1.325 ;
        RECT 2.625 1.325 2.805 1.445 ;
        RECT 2.625 1.445 4.175 1.7 ;
        RECT 3.845 0.985 4.175 1.445 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975 0.985 3.645 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.933750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 2.025 0.875 ;
        RECT 0.085 0.875 0.34 1.495 ;
        RECT 0.085 1.495 1.64 1.705 ;
        RECT 0.595 1.705 0.78 2.465 ;
        RECT 0.985 0.255 1.175 0.615 ;
        RECT 0.985 0.615 2.025 0.635 ;
        RECT 1.45 1.705 1.64 2.465 ;
        RECT 1.845 0.255 2.025 0.615 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.09 1.875 0.425 2.635 ;
      RECT 0.485 0.085 0.815 0.465 ;
      RECT 0.525 1.045 2.37 1.325 ;
      RECT 0.95 1.875 1.28 2.635 ;
      RECT 1.345 0.085 1.675 0.445 ;
      RECT 1.81 1.835 2.06 2.635 ;
      RECT 2.185 1.325 2.37 1.505 ;
      RECT 2.185 1.505 2.455 1.675 ;
      RECT 2.195 0.615 5.49 0.805 ;
      RECT 2.195 0.805 2.37 1.045 ;
      RECT 2.22 0.085 2.555 0.445 ;
      RECT 2.28 1.675 2.455 1.87 ;
      RECT 2.28 1.87 3.51 2.04 ;
      RECT 2.32 2.21 4.45 2.465 ;
      RECT 2.725 0.255 2.97 0.615 ;
      RECT 3.14 0.085 3.47 0.445 ;
      RECT 3.64 0.255 4.02 0.615 ;
      RECT 4.12 1.88 6.345 2.105 ;
      RECT 4.12 2.105 4.45 2.21 ;
      RECT 4.19 0.085 4.56 0.445 ;
      RECT 4.62 2.275 4.95 2.635 ;
      RECT 5.16 0.275 5.49 0.615 ;
      RECT 5.16 2.105 5.42 2.465 ;
      RECT 5.59 2.275 5.92 2.635 ;
      RECT 6.015 0.085 6.345 0.805 ;
      RECT 6.015 1.535 6.345 1.88 ;
      RECT 6.09 2.105 6.345 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__a211o_4
MACRO sky130_fd_sc_hd__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.045 2.45 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.045 1.81 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.62 1.045 3.07 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.045 3.595 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.452000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.255 0.775 0.635 ;
        RECT 0.555 0.635 0.785 2.335 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 0.085 0.385 0.905 ;
      RECT 0.09 1.49 0.385 2.635 ;
      RECT 0.945 0.085 1.795 0.445 ;
      RECT 1 0.695 3.585 0.875 ;
      RECT 1 0.875 1.31 1.49 ;
      RECT 1 1.49 3.585 1.66 ;
      RECT 1 1.83 1.255 2.635 ;
      RECT 1.455 1.84 2.795 2.02 ;
      RECT 1.455 2.02 1.785 2.465 ;
      RECT 1.955 2.19 2.23 2.635 ;
      RECT 2.275 0.275 2.605 0.695 ;
      RECT 2.465 2.02 2.795 2.465 ;
      RECT 2.81 0.085 3.085 0.525 ;
      RECT 3.255 0.275 3.585 0.695 ;
      RECT 3.255 1.66 3.585 2.325 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a211o_2
MACRO sky130_fd_sc_hd__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.93 1.075 1.625 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.67 1.445 ;
        RECT 0.425 1.445 1.965 1.615 ;
        RECT 1.795 1.075 2.395 1.245 ;
        RECT 1.795 1.245 1.965 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.525000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 2.125 2.645 2.295 ;
        RECT 2.475 1.755 3.135 1.955 ;
        RECT 2.475 1.955 2.645 2.125 ;
        RECT 2.815 0.345 3.135 0.825 ;
        RECT 2.965 0.825 3.135 1.755 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.28 0.55 0.825 ;
      RECT 0.085 0.825 0.255 1.785 ;
      RECT 0.085 1.785 2.305 1.955 ;
      RECT 0.085 2.125 0.385 2.635 ;
      RECT 0.555 1.955 0.885 2.465 ;
      RECT 1.055 0.085 1.225 0.905 ;
      RECT 1.055 2.125 1.685 2.635 ;
      RECT 1.395 0.255 1.725 0.735 ;
      RECT 1.395 0.735 2.645 0.825 ;
      RECT 1.395 0.825 2.305 0.905 ;
      RECT 1.895 0.085 2.245 0.475 ;
      RECT 2.135 0.655 2.645 0.735 ;
      RECT 2.135 1.415 2.795 1.585 ;
      RECT 2.135 1.585 2.305 1.785 ;
      RECT 2.415 0.255 2.645 0.655 ;
      RECT 2.625 0.995 2.795 1.415 ;
      RECT 2.815 2.125 3.115 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__xnor2_1
MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.255 1.075 2.705 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485 1.075 0.96 1.285 ;
        RECT 0.79 1.285 0.96 1.445 ;
        RECT 0.79 1.445 3.1 1.615 ;
        RECT 2.93 1.075 3.955 1.285 ;
        RECT 2.93 1.285 3.1 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.913000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.795 5.295 1.965 ;
        RECT 3.725 1.965 3.935 2.125 ;
        RECT 4.585 0.305 5.895 0.475 ;
        RECT 5.045 1.415 5.895 1.625 ;
        RECT 5.045 1.625 5.295 1.795 ;
        RECT 5.045 1.965 5.295 2.125 ;
        RECT 5.505 0.475 5.895 1.415 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.645 0.86 0.895 ;
      RECT 0.085 0.895 0.315 1.785 ;
      RECT 0.085 1.785 3.48 1.955 ;
      RECT 0.085 1.955 2.08 1.965 ;
      RECT 0.085 1.965 0.4 2.465 ;
      RECT 0.105 0.255 1.28 0.475 ;
      RECT 0.57 2.135 0.82 2.635 ;
      RECT 0.99 1.965 1.24 2.465 ;
      RECT 1.03 0.475 1.28 0.725 ;
      RECT 1.03 0.725 2.12 0.905 ;
      RECT 1.41 2.135 1.66 2.635 ;
      RECT 1.45 0.085 1.62 0.555 ;
      RECT 1.79 0.255 2.12 0.725 ;
      RECT 1.83 1.965 2.08 2.465 ;
      RECT 2.39 2.125 2.64 2.465 ;
      RECT 2.43 0.085 2.6 0.905 ;
      RECT 2.77 0.255 3.1 0.725 ;
      RECT 2.77 0.725 5.335 0.905 ;
      RECT 2.81 2.135 3.06 2.635 ;
      RECT 3.23 2.125 3.555 2.295 ;
      RECT 3.23 2.295 4.355 2.465 ;
      RECT 3.27 0.085 3.44 0.555 ;
      RECT 3.31 1.455 4.805 1.625 ;
      RECT 3.31 1.625 3.48 1.785 ;
      RECT 3.61 0.255 3.975 0.725 ;
      RECT 4.105 2.135 4.355 2.295 ;
      RECT 4.145 0.085 4.315 0.555 ;
      RECT 4.625 2.135 4.875 2.635 ;
      RECT 4.635 1.075 5.295 1.245 ;
      RECT 4.635 1.245 4.805 1.455 ;
      RECT 5.005 0.645 5.335 0.725 ;
      RECT 5.465 1.795 5.895 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.465 2.125 2.635 2.295 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.385 2.125 3.555 2.295 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 2.405 2.095 2.695 2.14 ;
      RECT 2.405 2.14 3.615 2.28 ;
      RECT 2.405 2.28 2.695 2.325 ;
      RECT 3.325 2.095 3.615 2.14 ;
      RECT 3.325 2.28 3.615 2.325 ;
  END
END sky130_fd_sc_hd__xnor2_2
MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175 1.075 5.39 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 1.075 1.855 1.275 ;
        RECT 1.685 1.275 1.855 1.445 ;
        RECT 1.685 1.445 5.73 1.615 ;
        RECT 5.56 1.075 7.43 1.275 ;
        RECT 5.56 1.275 5.73 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.721000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.16 1.785 8.25 2.045 ;
        RECT 7.96 1.445 10.035 1.665 ;
        RECT 7.96 1.665 8.25 1.785 ;
        RECT 7.96 2.045 8.25 2.465 ;
        RECT 8.38 0.645 10.035 0.905 ;
        RECT 8.84 1.665 9.09 2.465 ;
        RECT 9.68 1.665 10.035 2.465 ;
        RECT 9.815 0.905 10.035 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.085 0.645 1.76 0.905 ;
      RECT 0.085 0.905 0.32 1.445 ;
      RECT 0.085 1.445 1.3 1.615 ;
      RECT 0.085 1.615 0.46 2.465 ;
      RECT 0.17 0.255 2.18 0.475 ;
      RECT 0.63 1.835 0.88 2.635 ;
      RECT 1.05 1.615 1.3 1.785 ;
      RECT 1.05 1.785 3.82 2.005 ;
      RECT 1.05 2.005 1.3 2.465 ;
      RECT 1.47 2.175 1.72 2.635 ;
      RECT 1.89 2.005 2.14 2.465 ;
      RECT 1.93 0.475 2.18 0.725 ;
      RECT 1.93 0.725 3.86 0.905 ;
      RECT 2.31 2.175 2.56 2.635 ;
      RECT 2.35 0.085 2.52 0.555 ;
      RECT 2.69 0.255 3.02 0.725 ;
      RECT 2.73 2.005 2.98 2.465 ;
      RECT 3.15 2.175 3.4 2.635 ;
      RECT 3.19 0.085 3.36 0.555 ;
      RECT 3.53 0.255 3.86 0.725 ;
      RECT 3.57 2.005 3.82 2.465 ;
      RECT 4.035 0.085 4.31 0.905 ;
      RECT 4.035 1.785 5.99 2.005 ;
      RECT 4.035 2.005 4.35 2.465 ;
      RECT 4.48 0.255 4.81 0.725 ;
      RECT 4.48 0.725 7.43 0.735 ;
      RECT 4.48 0.735 8.21 0.905 ;
      RECT 4.52 2.175 4.77 2.635 ;
      RECT 4.94 2.005 5.19 2.465 ;
      RECT 4.98 0.085 5.15 0.555 ;
      RECT 5.32 0.255 5.65 0.725 ;
      RECT 5.36 2.175 5.61 2.635 ;
      RECT 5.78 2.005 5.99 2.215 ;
      RECT 5.78 2.215 7.75 2.465 ;
      RECT 5.82 0.085 5.99 0.555 ;
      RECT 5.9 1.445 7.77 1.615 ;
      RECT 6.16 0.255 6.49 0.725 ;
      RECT 6.66 0.085 6.83 0.555 ;
      RECT 7 0.255 7.33 0.725 ;
      RECT 7.5 0.085 7.77 0.555 ;
      RECT 7.6 1.075 9.645 1.275 ;
      RECT 7.6 1.275 7.77 1.445 ;
      RECT 7.96 0.305 9.97 0.475 ;
      RECT 7.96 0.475 8.21 0.735 ;
      RECT 8.42 1.835 8.67 2.635 ;
      RECT 9.26 1.835 9.51 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 1.445 1.235 1.615 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 1.445 6.295 1.615 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
    LAYER met1 ;
      RECT 1.005 1.415 1.295 1.46 ;
      RECT 1.005 1.46 6.355 1.6 ;
      RECT 1.005 1.6 1.295 1.645 ;
      RECT 6.065 1.415 6.355 1.46 ;
      RECT 6.065 1.6 6.355 1.645 ;
  END
END sky130_fd_sc_hd__xnor2_4
MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.465 0.305 10.795 2.42 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.795 1.125 4.98 1.72 ;
      RECT 4.815 0.735 5.32 0.955 ;
      RECT 4.915 2.175 5.955 2.375 ;
      RECT 5.005 0.255 5.68 0.565 ;
      RECT 5.15 0.955 5.32 1.655 ;
      RECT 5.15 1.655 5.615 2.005 ;
      RECT 5.51 0.565 5.68 1.315 ;
      RECT 5.51 1.315 6.36 1.485 ;
      RECT 5.785 1.485 6.36 1.575 ;
      RECT 5.785 1.575 5.955 2.175 ;
      RECT 5.87 0.765 6.935 1.045 ;
      RECT 5.87 1.045 7.445 1.065 ;
      RECT 5.87 1.065 6.07 1.095 ;
      RECT 5.945 0.085 6.34 0.56 ;
      RECT 6.125 1.835 6.36 2.635 ;
      RECT 6.19 1.245 6.36 1.315 ;
      RECT 6.53 0.255 6.935 0.765 ;
      RECT 6.53 1.065 7.445 1.375 ;
      RECT 6.53 1.375 6.86 2.465 ;
      RECT 7.07 2.105 7.36 2.635 ;
      RECT 7.165 0.085 7.44 0.615 ;
      RECT 7.79 1.245 7.98 1.965 ;
      RECT 7.925 2.165 8.81 2.355 ;
      RECT 8.005 0.705 8.47 1.035 ;
      RECT 8.025 0.33 8.81 0.535 ;
      RECT 8.15 1.035 8.47 1.995 ;
      RECT 8.64 0.535 8.81 0.995 ;
      RECT 8.64 0.995 9.51 1.325 ;
      RECT 8.64 1.325 8.81 2.165 ;
      RECT 8.98 1.53 9.88 1.905 ;
      RECT 8.98 2.135 9.24 2.635 ;
      RECT 9.05 0.085 9.365 0.615 ;
      RECT 9.54 1.905 9.88 2.465 ;
      RECT 9.55 0.3 9.88 0.825 ;
      RECT 9.69 0.825 9.88 1.53 ;
      RECT 10.05 0.085 10.295 0.9 ;
      RECT 10.05 1.465 10.295 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.21 1.785 5.38 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.8 1.785 7.97 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.22 1.445 8.39 1.615 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.7 0.765 9.87 0.935 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 8.03 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 8.45 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 9.93 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.15 1.755 5.44 1.8 ;
      RECT 5.15 1.94 5.44 1.985 ;
      RECT 7.74 1.755 8.03 1.8 ;
      RECT 7.74 1.94 8.03 1.985 ;
      RECT 8.16 1.415 8.45 1.46 ;
      RECT 8.16 1.6 8.45 1.645 ;
      RECT 9.64 0.735 9.93 0.78 ;
      RECT 9.64 0.92 9.93 0.965 ;
  END
END sky130_fd_sc_hd__edfxtp_1
MACRO sky130_fd_sc_hd__diode_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__diode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 4.6 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  0.434700 ;
    ANTENNAGATEAREA  0.434700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.835 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 0.92 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.11 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.92 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.92 0.085 ;
      RECT 0 2.635 0.92 2.805 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
  END
END sky130_fd_sc_hd__diode_2
MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.48 1.285 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.390500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.185 0.27 3.625 0.64 ;
        RECT 3.185 1.53 3.625 2.465 ;
        RECT 3.345 0.64 3.625 1.53 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.27 0.415 0.735 ;
      RECT 0.085 0.735 1.27 0.905 ;
      RECT 0.085 1.455 1.27 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.585 0.085 0.915 0.565 ;
      RECT 0.6 1.8 0.93 2.635 ;
      RECT 0.765 1.075 1.435 1.245 ;
      RECT 0.85 0.905 1.27 1.075 ;
      RECT 0.85 1.245 1.27 1.455 ;
      RECT 1.39 1.785 1.795 2.465 ;
      RECT 1.44 0.27 1.795 0.9 ;
      RECT 1.625 0.9 1.795 1.075 ;
      RECT 1.625 1.075 2.305 1.245 ;
      RECT 1.625 1.245 1.795 1.785 ;
      RECT 1.985 0.27 2.235 0.735 ;
      RECT 1.985 0.735 2.645 0.905 ;
      RECT 1.985 1.46 2.645 1.63 ;
      RECT 1.985 1.63 2.235 2.465 ;
      RECT 2.475 0.905 2.645 0.995 ;
      RECT 2.475 0.995 3.175 1.325 ;
      RECT 2.475 1.325 2.645 1.46 ;
      RECT 2.685 0.085 3.015 0.565 ;
      RECT 2.685 1.8 3.015 2.635 ;
      RECT 3.795 0.085 4.055 0.635 ;
      RECT 3.795 1.8 4.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2
MACRO sky130_fd_sc_hd__clkdlybuf4s50_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.535 1.29 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.255 3.595 0.64 ;
        RECT 3.19 1.69 3.595 2.465 ;
        RECT 3.345 0.64 3.595 1.69 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.255 0.415 0.735 ;
      RECT 0.085 0.735 1.055 0.905 ;
      RECT 0.085 1.46 1.055 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.585 0.085 0.915 0.565 ;
      RECT 0.6 1.8 0.93 2.635 ;
      RECT 0.705 0.905 1.055 1.025 ;
      RECT 0.705 1.025 1.135 1.315 ;
      RECT 0.705 1.315 1.055 1.46 ;
      RECT 1.38 0.255 1.73 1.07 ;
      RECT 1.38 1.07 2.24 1.32 ;
      RECT 1.38 1.32 1.73 2.465 ;
      RECT 1.99 0.255 2.24 0.73 ;
      RECT 1.99 0.73 2.58 0.9 ;
      RECT 1.99 1.495 2.58 1.665 ;
      RECT 1.99 1.665 2.24 2.465 ;
      RECT 2.41 0.9 2.58 0.995 ;
      RECT 2.41 0.995 3.175 1.325 ;
      RECT 2.41 1.325 2.58 1.495 ;
      RECT 2.69 0.085 3.02 0.6 ;
      RECT 2.69 1.835 3.02 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_1
MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.075 3.22 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.075 4.48 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.715 1.075 5.86 1.625 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.08 1.725 1.285 ;
        RECT 1.175 1.075 1.505 1.08 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.825 1.285 ;
        RECT 0.145 1.285 0.325 1.625 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.955 0.845 2.125 ;
        RECT 0.595 1.455 2.18 1.625 ;
        RECT 0.595 1.625 0.765 1.955 ;
        RECT 1.355 0.655 3.1 0.825 ;
        RECT 1.435 1.625 1.605 2.125 ;
        RECT 1.965 0.825 2.18 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.095 0.295 0.425 0.465 ;
      RECT 0.175 0.465 0.345 0.715 ;
      RECT 0.175 0.715 1.185 0.885 ;
      RECT 0.175 1.795 0.345 2.295 ;
      RECT 0.175 2.295 2.025 2.465 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.935 0.295 2.115 0.465 ;
      RECT 1.015 0.465 1.185 0.715 ;
      RECT 1.015 1.795 1.185 2.295 ;
      RECT 1.855 1.795 2.025 1.915 ;
      RECT 1.855 1.915 5.805 2.085 ;
      RECT 1.855 2.085 2.025 2.295 ;
      RECT 2.27 2.255 2.94 2.635 ;
      RECT 2.35 0.295 4.37 0.465 ;
      RECT 3.18 1.795 3.35 1.915 ;
      RECT 3.18 2.085 3.35 2.465 ;
      RECT 3.55 2.255 4.22 2.635 ;
      RECT 3.62 0.635 5.39 0.805 ;
      RECT 4.39 1.795 4.56 1.915 ;
      RECT 4.39 2.085 4.56 2.465 ;
      RECT 4.555 0.085 4.89 0.465 ;
      RECT 4.765 2.255 5.435 2.635 ;
      RECT 5.06 0.275 5.39 0.635 ;
      RECT 5.56 0.085 5.885 0.885 ;
      RECT 5.635 1.795 5.805 1.915 ;
      RECT 5.635 2.085 5.805 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__a32oi_2
MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.23 1.075 1.595 1.255 ;
        RECT 1.405 0.345 1.705 0.765 ;
        RECT 1.405 0.765 1.595 1.075 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.995 2.165 1.325 ;
        RECT 1.965 0.415 2.165 0.995 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.015 2.75 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.995 1.025 1.425 ;
        RECT 0.855 1.425 1.255 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.575500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 1.165 0.805 ;
        RECT 0.515 0.805 0.685 1.785 ;
        RECT 0.515 1.785 0.865 2.085 ;
        RECT 0.915 0.295 1.165 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.835 0.345 2.255 ;
      RECT 0.085 2.255 1.345 2.465 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 1.095 1.785 2.185 1.955 ;
      RECT 1.095 1.955 1.345 2.255 ;
      RECT 1.555 2.135 1.805 2.635 ;
      RECT 2.015 1.745 2.185 1.785 ;
      RECT 2.015 1.955 2.185 2.465 ;
      RECT 2.355 0.085 2.695 0.805 ;
      RECT 2.355 1.495 2.695 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a32oi_1
MACRO sky130_fd_sc_hd__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 5.465 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.075 7.695 1.3 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.295 1.075 9.985 1.28 ;
        RECT 9.805 0.755 9.985 1.075 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.585 0.995 3.555 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.75 1.305 ;
        RECT 0.11 1.305 0.33 1.965 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.575 3.365 1.745 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 1.355 1.745 1.685 2.085 ;
        RECT 1.975 0.99 2.365 1.575 ;
        RECT 1.975 1.745 2.525 2.085 ;
        RECT 2.195 0.635 5.565 0.805 ;
        RECT 2.195 0.805 2.365 0.99 ;
        RECT 3.035 1.745 3.365 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.095 2.255 3.705 2.425 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 2.025 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.355 0.085 1.685 0.465 ;
      RECT 1.855 0.295 3.785 0.465 ;
      RECT 1.855 0.465 2.025 0.635 ;
      RECT 3.535 1.575 9.925 1.745 ;
      RECT 3.535 1.745 3.705 2.255 ;
      RECT 3.895 1.915 4.225 2.635 ;
      RECT 3.975 0.295 7.805 0.465 ;
      RECT 4.395 1.745 4.565 2.465 ;
      RECT 4.77 1.915 5.44 2.635 ;
      RECT 5.64 1.745 5.81 2.465 ;
      RECT 6.215 0.635 9.505 0.805 ;
      RECT 6.215 1.915 6.545 2.635 ;
      RECT 6.715 1.745 6.885 2.465 ;
      RECT 7.055 1.915 7.385 2.635 ;
      RECT 7.555 1.745 7.725 2.465 ;
      RECT 7.995 0.085 8.325 0.465 ;
      RECT 8.415 1.915 8.745 2.635 ;
      RECT 8.495 0.255 8.665 0.635 ;
      RECT 8.835 0.085 9.165 0.465 ;
      RECT 8.915 1.745 9.085 2.465 ;
      RECT 9.255 1.915 9.585 2.635 ;
      RECT 9.335 0.255 9.505 0.635 ;
      RECT 9.685 0.085 10.025 0.465 ;
      RECT 9.755 1.745 9.925 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__a32oi_4
MACRO sky130_fd_sc_hd__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.865 0.255 10.125 0.825 ;
        RECT 9.865 1.445 10.125 2.465 ;
        RECT 9.91 0.825 10.125 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.37 0.255 8.7 2.465 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
      LAYER mcon ;
        RECT 3.825 0.765 3.995 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
      LAYER mcon ;
        RECT 7.045 0.765 7.215 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.77 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.58 0.085 ;
      RECT 0 2.635 10.58 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.43 2.255 3.81 2.635 ;
      RECT 3.61 0.085 4.02 0.525 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.33 2.255 4.66 2.635 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.74 0.085 5.08 0.545 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.47 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.78 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.83 1.745 ;
      RECT 5.93 2.255 6.34 2.635 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 6.67 0.085 7.33 0.565 ;
      RECT 7.01 1.945 7.34 2.635 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.83 0.68 ;
      RECT 7.51 1.745 7.83 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.83 1.575 ;
      RECT 8.02 0.085 8.2 0.905 ;
      RECT 8.02 1.48 8.2 2.635 ;
      RECT 8.89 0.255 9.22 0.995 ;
      RECT 8.89 0.995 9.74 1.325 ;
      RECT 8.89 1.325 9.22 2.465 ;
      RECT 9.445 0.085 9.615 0.585 ;
      RECT 9.445 1.825 9.615 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.245 1.105 5.415 1.275 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 5.435 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.475 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.185 1.075 5.475 1.12 ;
      RECT 5.185 1.26 5.475 1.305 ;
  END
END sky130_fd_sc_hd__dfsbp_1
MACRO sky130_fd_sc_hd__dfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.15 1.495 10.915 1.665 ;
        RECT 10.15 1.665 10.48 2.465 ;
        RECT 10.23 0.255 10.48 0.72 ;
        RECT 10.23 0.72 10.915 0.825 ;
        RECT 10.345 0.825 10.915 0.845 ;
        RECT 10.36 0.845 10.915 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.37 0.255 8.7 2.465 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
      LAYER mcon ;
        RECT 3.825 0.765 3.995 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
      LAYER mcon ;
        RECT 7.045 0.765 7.215 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.43 2.255 3.81 2.635 ;
      RECT 3.61 0.085 4.02 0.525 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.33 2.255 4.66 2.635 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.74 0.085 5.08 0.545 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.47 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.78 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.83 1.745 ;
      RECT 5.93 2.255 6.34 2.635 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 6.67 0.085 7.33 0.565 ;
      RECT 7.01 1.945 7.34 2.635 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.83 0.68 ;
      RECT 7.51 1.745 7.83 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.83 1.575 ;
      RECT 8.02 0.085 8.2 0.905 ;
      RECT 8.02 1.48 8.2 2.635 ;
      RECT 8.87 0.085 9.12 0.905 ;
      RECT 8.87 1.48 9.12 2.635 ;
      RECT 9.31 0.255 9.56 0.995 ;
      RECT 9.31 0.995 10.19 1.325 ;
      RECT 9.31 1.325 9.64 2.465 ;
      RECT 9.73 0.085 10.06 0.825 ;
      RECT 9.81 1.495 9.98 2.635 ;
      RECT 10.65 0.085 10.915 0.55 ;
      RECT 10.65 1.835 10.915 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.245 1.105 5.415 1.275 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 5.435 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.475 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.185 1.075 5.475 1.12 ;
      RECT 5.185 1.26 5.475 1.305 ;
  END
END sky130_fd_sc_hd__dfsbp_2
MACRO sky130_fd_sc_hd__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.225 0.255 11.555 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.4 1.065 9.845 1.41 ;
        RECT 9.4 1.41 9.73 2.465 ;
        RECT 9.515 0.255 9.845 1.065 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.15 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.795 1.125 4.98 1.72 ;
      RECT 4.815 0.735 5.32 0.955 ;
      RECT 4.915 2.175 5.955 2.375 ;
      RECT 5.005 0.255 5.68 0.565 ;
      RECT 5.15 0.955 5.32 1.655 ;
      RECT 5.15 1.655 5.615 2.005 ;
      RECT 5.51 0.565 5.68 1.315 ;
      RECT 5.51 1.315 6.36 1.485 ;
      RECT 5.785 1.485 6.36 1.575 ;
      RECT 5.785 1.575 5.955 2.175 ;
      RECT 5.87 0.765 6.935 1.045 ;
      RECT 5.87 1.045 7.445 1.065 ;
      RECT 5.87 1.065 6.07 1.095 ;
      RECT 5.945 0.085 6.34 0.56 ;
      RECT 6.125 1.835 6.36 2.635 ;
      RECT 6.19 1.245 6.36 1.315 ;
      RECT 6.53 0.255 6.935 0.765 ;
      RECT 6.53 1.065 7.445 1.375 ;
      RECT 6.53 1.375 6.86 2.465 ;
      RECT 7.07 2.105 7.36 2.635 ;
      RECT 7.165 0.085 7.44 0.615 ;
      RECT 7.79 1.245 7.98 1.965 ;
      RECT 7.925 2.165 8.89 2.355 ;
      RECT 8.005 0.705 8.47 1.035 ;
      RECT 8.025 0.33 8.89 0.535 ;
      RECT 8.15 1.035 8.47 1.995 ;
      RECT 8.64 0.535 8.89 2.165 ;
      RECT 9.06 1.495 9.23 2.635 ;
      RECT 9.095 0.085 9.345 0.9 ;
      RECT 9.9 1.575 10.13 2.01 ;
      RECT 10.015 0.89 10.64 1.22 ;
      RECT 10.3 0.255 10.64 0.89 ;
      RECT 10.3 1.22 10.64 2.465 ;
      RECT 10.81 0.085 11.055 0.9 ;
      RECT 10.81 1.465 11.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.21 1.785 5.38 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.8 1.785 7.97 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.22 1.445 8.39 1.615 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.68 1.785 8.85 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 9.93 1.785 10.1 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.39 0.765 10.56 0.935 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 8.03 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 8.45 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 10.62 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.15 1.755 5.44 1.8 ;
      RECT 5.15 1.94 5.44 1.985 ;
      RECT 7.74 1.755 8.03 1.8 ;
      RECT 7.74 1.94 8.03 1.985 ;
      RECT 8.16 1.415 8.45 1.46 ;
      RECT 8.16 1.6 8.45 1.645 ;
      RECT 8.62 1.755 8.91 1.8 ;
      RECT 8.62 1.8 10.16 1.94 ;
      RECT 8.62 1.94 8.91 1.985 ;
      RECT 9.87 1.755 10.16 1.8 ;
      RECT 9.87 1.94 10.16 1.985 ;
      RECT 10.33 0.735 10.62 0.78 ;
      RECT 10.33 0.92 10.62 0.965 ;
  END
END sky130_fd_sc_hd__edfxbp_1
MACRO sky130_fd_sc_hd__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.67 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165 1.075 2.495 1.325 ;
        RECT 2.315 1.325 2.495 1.445 ;
        RECT 2.315 1.445 2.645 1.615 ;
        RECT 2.445 1.615 2.645 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 1.075 1.335 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 1.075 1.995 1.325 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.535 0.715 1.785 0.895 ;
      RECT 0.535 0.895 0.81 1.495 ;
      RECT 0.535 1.495 2.145 1.705 ;
      RECT 0.555 1.875 1.34 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 1.035 0.295 2.285 0.475 ;
      RECT 1.42 0.645 1.785 0.715 ;
      RECT 1.735 1.705 2.145 1.805 ;
      RECT 1.735 1.805 2.12 2.465 ;
      RECT 1.955 0.475 2.285 0.695 ;
      RECT 1.955 0.695 3.135 0.865 ;
      RECT 2.455 0.085 2.625 0.525 ;
      RECT 2.795 0.28 3.135 0.695 ;
      RECT 2.815 1.455 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o22a_1
MACRO sky130_fd_sc_hd__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.075 3.59 1.275 ;
        RECT 3.27 1.275 3.59 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595 1.075 2.925 1.325 ;
        RECT 2.745 1.325 2.925 1.445 ;
        RECT 2.745 1.445 3.1 1.615 ;
        RECT 2.9 1.615 3.1 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.075 1.79 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 1.075 2.425 1.325 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.365 0.805 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.13 -0.085 0.3 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.115 1.445 0.365 2.635 ;
      RECT 0.185 0.085 0.355 0.885 ;
      RECT 0.975 0.715 2.215 0.895 ;
      RECT 0.975 0.895 1.255 1.495 ;
      RECT 0.975 1.495 2.575 1.705 ;
      RECT 0.995 1.875 1.795 2.635 ;
      RECT 1.025 0.085 1.205 0.545 ;
      RECT 1.465 0.295 2.73 0.475 ;
      RECT 1.85 0.645 2.215 0.715 ;
      RECT 2.19 1.705 2.575 2.465 ;
      RECT 2.39 0.475 2.73 0.695 ;
      RECT 2.39 0.695 3.59 0.825 ;
      RECT 2.56 0.825 3.59 0.865 ;
      RECT 2.915 0.085 3.085 0.525 ;
      RECT 3.255 0.28 3.59 0.695 ;
      RECT 3.27 1.795 3.59 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o22a_2
MACRO sky130_fd_sc_hd__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.35 1.075 4.68 1.445 ;
        RECT 4.35 1.445 5.735 1.615 ;
        RECT 5.565 1.075 6.355 1.275 ;
        RECT 5.565 1.275 5.735 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.9 1.075 5.395 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.42 1.075 2.955 1.445 ;
        RECT 2.42 1.445 4.18 1.615 ;
        RECT 3.85 1.075 4.18 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.68 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.725 1.77 0.905 ;
        RECT 0.085 0.905 0.37 1.445 ;
        RECT 0.085 1.445 1.73 1.615 ;
        RECT 0.6 0.265 0.93 0.725 ;
        RECT 0.64 1.615 0.89 2.465 ;
        RECT 1.44 0.255 1.77 0.725 ;
        RECT 1.48 1.615 1.73 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.22 1.825 0.47 2.635 ;
      RECT 0.26 0.085 0.43 0.555 ;
      RECT 0.54 1.075 2.23 1.275 ;
      RECT 1.06 1.795 1.31 2.635 ;
      RECT 1.1 0.085 1.27 0.555 ;
      RECT 1.9 1.275 2.23 1.785 ;
      RECT 1.9 1.785 5.27 1.955 ;
      RECT 1.9 2.125 2.67 2.635 ;
      RECT 1.94 0.085 2.11 0.555 ;
      RECT 1.94 0.735 3.97 0.905 ;
      RECT 1.94 0.905 2.23 1.075 ;
      RECT 2.38 0.255 4.47 0.475 ;
      RECT 2.415 0.645 3.97 0.735 ;
      RECT 2.84 2.125 3.09 2.295 ;
      RECT 2.84 2.295 3.93 2.465 ;
      RECT 3.26 1.955 3.51 2.125 ;
      RECT 3.68 2.125 3.93 2.295 ;
      RECT 4.1 2.125 4.43 2.635 ;
      RECT 4.14 0.475 4.47 0.735 ;
      RECT 4.14 0.735 6.15 0.905 ;
      RECT 4.6 2.125 4.85 2.295 ;
      RECT 4.6 2.295 5.69 2.465 ;
      RECT 4.64 0.085 4.81 0.555 ;
      RECT 4.98 0.255 5.31 0.725 ;
      RECT 4.98 0.725 6.15 0.735 ;
      RECT 5.02 1.955 5.27 2.125 ;
      RECT 5.44 1.785 5.69 2.295 ;
      RECT 5.48 0.085 5.65 0.555 ;
      RECT 5.82 0.255 6.15 0.725 ;
      RECT 5.905 1.455 6.11 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__o22a_4
MACRO sky130_fd_sc_hd__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT -1.14 0.77 0.04 1.95 ;
        RECT 1.46 0.77 2.64 1.95 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.26 0.56 2.76 2.16 ;
        RECT 1.16 -1.105 2.76 0.56 ;
        RECT 1.16 2.16 2.76 3.825 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 4.36 -1.17 6.675 0.56 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 4.36 2.16 6.675 3.89 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.595 1.835 0.765 2.635 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.355 0.085 1.685 0.565 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
      RECT 1.435 1.835 1.605 2.635 ;
      RECT 1.855 0.255 2.025 0.735 ;
      RECT 1.855 0.735 4.545 0.905 ;
      RECT 1.855 1.445 4.545 1.615 ;
      RECT 1.855 1.615 2.025 2.465 ;
      RECT 2.195 0.085 2.525 0.565 ;
      RECT 2.195 1.835 2.525 2.635 ;
      RECT 2.695 0.255 2.865 0.735 ;
      RECT 2.695 1.615 2.865 2.465 ;
      RECT 3.035 0.085 3.365 0.565 ;
      RECT 3.035 1.835 3.365 2.635 ;
      RECT 3.535 0.255 3.705 0.735 ;
      RECT 3.535 1.615 3.705 2.465 ;
      RECT 3.875 0.085 4.205 0.565 ;
      RECT 3.875 1.835 4.205 2.635 ;
      RECT 4.29 0.905 4.545 1.055 ;
      RECT 4.29 1.055 4.87 1.315 ;
      RECT 4.29 1.315 4.545 1.445 ;
      RECT 4.375 0.255 4.545 0.735 ;
      RECT 4.375 1.615 4.545 2.465 ;
      RECT 4.715 0.085 5.045 0.885 ;
      RECT 4.715 1.485 5.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.305 1.105 4.475 1.275 ;
      RECT 4.665 1.105 4.835 1.275 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
    LAYER met1 ;
      RECT 0 -0.24 5.52 -0.13 ;
      RECT 0 -0.13 5.84 0.13 ;
      RECT 0 0.13 5.52 0.24 ;
      RECT 0 2.48 5.52 2.59 ;
      RECT 0 2.59 5.84 2.85 ;
      RECT 0 2.85 5.52 2.96 ;
      RECT 2.02 1.06 2.66 1.12 ;
      RECT 2.02 1.12 4.895 1.26 ;
      RECT 2.02 1.26 2.66 1.32 ;
      RECT 4.245 1.075 4.895 1.12 ;
      RECT 4.245 1.26 4.895 1.305 ;
    LAYER met2 ;
      RECT 1.89 1.05 2.66 1.33 ;
      RECT 5.135 -0.14 5.905 0.14 ;
      RECT 5.135 2.58 5.905 2.86 ;
    LAYER met3 ;
      RECT -0.715 1.03 0.065 1.35 ;
      RECT 1.885 1.025 2.665 1.355 ;
      RECT 5.13 -0.165 5.91 0.165 ;
      RECT 5.13 2.555 5.91 2.885 ;
    LAYER met4 ;
      RECT 4.93 -0.895 6.11 0.285 ;
      RECT 4.93 2.435 6.11 3.615 ;
    LAYER via ;
      RECT 2.05 1.06 2.31 1.32 ;
      RECT 2.37 1.06 2.63 1.32 ;
      RECT 5.23 -0.13 5.49 0.13 ;
      RECT 5.23 2.59 5.49 2.85 ;
      RECT 5.55 -0.13 5.81 0.13 ;
      RECT 5.55 2.59 5.81 2.85 ;
    LAYER via2 ;
      RECT 1.935 1.05 2.215 1.33 ;
      RECT 2.335 1.05 2.615 1.33 ;
      RECT 5.18 -0.14 5.46 0.14 ;
      RECT 5.18 2.58 5.46 2.86 ;
      RECT 5.58 -0.14 5.86 0.14 ;
      RECT 5.58 2.58 5.86 2.86 ;
    LAYER via3 ;
      RECT -0.685 1.03 -0.365 1.35 ;
      RECT -0.285 1.03 0.035 1.35 ;
      RECT 1.915 1.03 2.235 1.35 ;
      RECT 2.315 1.03 2.635 1.35 ;
      RECT 5.16 -0.16 5.48 0.16 ;
      RECT 5.16 2.56 5.48 2.88 ;
      RECT 5.56 -0.16 5.88 0.16 ;
      RECT 5.56 2.56 5.88 2.88 ;
  END
END sky130_fd_sc_hd__probec_p_8
MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.1 1.075 3.595 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 2.93 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
        RECT 0.595 1.325 0.775 1.695 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.255 1.24 0.595 ;
        RECT 0.945 0.595 1.115 1.495 ;
        RECT 0.945 1.495 1.35 1.695 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.43 0.345 0.825 ;
      RECT 0.085 0.825 0.255 1.495 ;
      RECT 0.085 1.495 0.395 1.865 ;
      RECT 0.085 1.865 1.935 2.035 ;
      RECT 0.52 2.205 0.91 2.635 ;
      RECT 0.595 0.085 0.775 0.825 ;
      RECT 1.285 0.89 1.595 1.06 ;
      RECT 1.285 1.06 1.455 1.325 ;
      RECT 1.41 0.085 1.77 0.485 ;
      RECT 1.415 2.205 2.23 2.635 ;
      RECT 1.425 0.655 2.275 0.825 ;
      RECT 1.425 0.825 1.595 0.89 ;
      RECT 1.765 0.995 1.935 1.865 ;
      RECT 1.94 0.255 2.275 0.655 ;
      RECT 2.105 0.825 2.275 1.455 ;
      RECT 2.105 1.455 2.725 2.035 ;
      RECT 2.4 2.035 2.725 2.465 ;
      RECT 2.445 0.365 2.745 0.735 ;
      RECT 2.445 0.735 3.59 0.905 ;
      RECT 2.915 0.085 3.085 0.555 ;
      RECT 3.2 1.875 3.53 2.635 ;
      RECT 3.255 0.27 3.59 0.735 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o21ba_2
MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.99 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 1.075 4.82 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.885 1.285 ;
        RECT 0.605 1.285 0.885 1.705 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.255 1.385 0.725 ;
        RECT 1.055 0.725 2.225 0.905 ;
        RECT 1.055 0.905 1.455 1.445 ;
        RECT 1.055 1.445 2.225 1.705 ;
        RECT 1.895 0.255 2.225 0.725 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.265 0.545 0.855 ;
      RECT 0.085 0.855 0.255 1.455 ;
      RECT 0.085 1.455 0.435 1.875 ;
      RECT 0.085 1.875 2.565 2.045 ;
      RECT 0.085 2.045 0.435 2.465 ;
      RECT 0.635 2.215 0.965 2.635 ;
      RECT 0.715 0.085 0.885 0.905 ;
      RECT 1.475 2.215 1.805 2.635 ;
      RECT 1.555 0.085 1.725 0.555 ;
      RECT 1.625 1.075 2.565 1.275 ;
      RECT 2.315 2.215 2.645 2.635 ;
      RECT 2.395 0.085 2.565 0.555 ;
      RECT 2.395 0.725 3.585 0.895 ;
      RECT 2.395 0.895 2.565 1.075 ;
      RECT 2.395 1.445 2.905 1.615 ;
      RECT 2.395 1.615 2.565 1.875 ;
      RECT 2.735 1.075 3.135 1.245 ;
      RECT 2.735 1.245 2.905 1.445 ;
      RECT 2.805 0.255 4.005 0.475 ;
      RECT 2.815 1.795 4.38 1.965 ;
      RECT 2.815 1.965 2.985 2.465 ;
      RECT 3.2 2.135 3.45 2.635 ;
      RECT 3.235 0.645 3.585 0.725 ;
      RECT 3.395 0.895 3.585 1.795 ;
      RECT 3.685 2.135 3.925 2.295 ;
      RECT 3.685 2.295 4.765 2.465 ;
      RECT 3.755 0.475 4.005 0.725 ;
      RECT 3.755 0.725 5.71 0.905 ;
      RECT 4.135 1.445 4.38 1.795 ;
      RECT 4.135 1.965 4.38 2.125 ;
      RECT 4.175 0.085 4.345 0.555 ;
      RECT 4.515 0.255 4.845 0.725 ;
      RECT 4.595 1.455 5.71 1.665 ;
      RECT 4.595 1.665 4.765 2.295 ;
      RECT 4.935 1.835 5.265 2.635 ;
      RECT 5.015 0.085 5.185 0.555 ;
      RECT 5.355 0.265 5.71 0.725 ;
      RECT 5.435 1.665 5.71 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__o21ba_4
MACRO sky130_fd_sc_hd__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.95 1.075 3.595 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 2.78 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.03 0.995 1.36 1.325 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.45 0.445 0.825 ;
        RECT 0.085 0.825 0.34 1.48 ;
        RECT 0.085 1.48 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.51 0.995 0.86 1.325 ;
      RECT 0.595 1.325 0.86 1.865 ;
      RECT 0.595 1.865 2.575 2.035 ;
      RECT 0.595 2.205 1.005 2.635 ;
      RECT 0.71 0.085 0.88 0.825 ;
      RECT 1.075 1.525 1.7 1.695 ;
      RECT 1.16 0.45 1.33 0.655 ;
      RECT 1.16 0.655 1.7 0.825 ;
      RECT 1.53 0.825 1.7 1.525 ;
      RECT 1.75 2.215 2.08 2.635 ;
      RECT 1.87 0.255 2.04 1.455 ;
      RECT 1.87 1.455 2.575 1.865 ;
      RECT 2.25 2.035 2.575 2.465 ;
      RECT 2.27 0.255 2.6 0.735 ;
      RECT 2.27 0.735 3.44 0.905 ;
      RECT 2.77 0.085 2.94 0.555 ;
      RECT 3.05 1.535 3.38 2.635 ;
      RECT 3.11 0.27 3.44 0.735 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o21ba_1
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.24 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.255 1.245 0.655 ;
        RECT 1.04 0.655 1.725 0.825 ;
        RECT 1.06 1.75 1.725 1.97 ;
        RECT 1.06 1.97 1.245 2.435 ;
        RECT 1.385 0.825 1.725 1.75 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.855 0.855 2.465 ;
      LAYER mcon ;
        RECT 0.61 2.125 0.78 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.415 2.14 1.75 2.465 ;
      LAYER mcon ;
        RECT 1.495 2.14 1.665 2.31 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
        RECT 1.435 2.08 1.725 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.41 ;
      RECT 0.085 1.41 1.215 1.58 ;
      RECT 0.085 1.58 0.355 2.435 ;
      RECT 0.555 0.085 0.83 0.565 ;
      RECT 0.965 0.995 1.215 1.41 ;
      RECT 1.415 0.085 1.75 0.485 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.28 1.68 0.735 ;
        RECT 1.42 0.735 4.73 0.905 ;
        RECT 1.42 1.495 4.73 1.735 ;
        RECT 1.42 1.735 1.68 2.46 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 3.76 0.905 4.73 1.495 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.525 0.39 2.465 ;
      LAYER mcon ;
        RECT 0.175 2.125 0.345 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.99 1.525 1.25 2.465 ;
      LAYER mcon ;
        RECT 1.035 2.125 1.205 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.85 1.905 2.11 2.465 ;
      LAYER mcon ;
        RECT 1.89 2.125 2.06 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.71 1.905 2.97 2.465 ;
      LAYER mcon ;
        RECT 2.74 2.125 2.91 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.57 1.905 3.83 2.465 ;
      LAYER mcon ;
        RECT 3.62 2.125 3.79 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.43 1.905 4.725 2.465 ;
      LAYER mcon ;
        RECT 4.48 2.125 4.65 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 4.99 2.34 ;
        RECT 0.115 2.08 0.405 2.14 ;
        RECT 0.975 2.08 1.265 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.68 2.08 2.97 2.14 ;
        RECT 3.56 2.08 3.85 2.14 ;
        RECT 4.42 2.08 4.71 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.145 0.085 0.39 0.545 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 3.59 1.325 ;
      RECT 0.57 1.325 0.82 2.46 ;
      RECT 0.99 0.085 1.25 0.61 ;
      RECT 1.85 0.085 2.11 0.565 ;
      RECT 2.71 0.085 2.97 0.565 ;
      RECT 3.57 0.085 3.83 0.565 ;
      RECT 4.43 0.085 4.73 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 0.735 9.025 0.905 ;
        RECT 2.315 1.495 9.025 1.72 ;
        RECT 2.315 1.72 7.685 1.735 ;
        RECT 2.315 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
        RECT 4.845 0.28 5.12 0.735 ;
        RECT 4.86 1.735 5.12 2.46 ;
        RECT 5.705 0.28 5.965 0.735 ;
        RECT 5.705 1.735 5.965 2.46 ;
        RECT 6.565 0.28 6.825 0.735 ;
        RECT 6.565 1.735 6.825 2.46 ;
        RECT 7.425 0.28 7.685 0.735 ;
        RECT 7.425 1.735 7.685 2.46 ;
        RECT 7.86 0.905 9.025 1.495 ;
        RECT 8.295 0.28 8.555 0.735 ;
        RECT 8.295 1.72 8.585 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.425 2.465 ;
      LAYER mcon ;
        RECT 0.175 2.125 0.345 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.955 1.495 1.285 2.465 ;
      LAYER mcon ;
        RECT 1.035 2.125 1.205 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.815 1.495 2.145 2.465 ;
      LAYER mcon ;
        RECT 1.89 2.125 2.06 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.71 1.905 2.97 2.465 ;
      LAYER mcon ;
        RECT 2.74 2.125 2.91 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.57 1.905 3.83 2.465 ;
      LAYER mcon ;
        RECT 3.62 2.125 3.79 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.43 1.905 4.69 2.465 ;
      LAYER mcon ;
        RECT 4.48 2.125 4.65 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.29 1.905 5.535 2.465 ;
      LAYER mcon ;
        RECT 5.335 2.125 5.505 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.15 1.905 6.395 2.465 ;
      LAYER mcon ;
        RECT 6.195 2.125 6.365 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.01 1.905 7.255 2.465 ;
      LAYER mcon ;
        RECT 7.05 2.125 7.22 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.87 1.905 8.125 2.465 ;
      LAYER mcon ;
        RECT 7.9 2.125 8.07 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.755 1.89 9.025 2.465 ;
      LAYER mcon ;
        RECT 8.78 2.125 8.95 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 9.13 2.34 ;
        RECT 0.115 2.08 0.405 2.14 ;
        RECT 0.975 2.08 1.265 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.68 2.08 2.97 2.14 ;
        RECT 3.56 2.08 3.85 2.14 ;
        RECT 4.42 2.08 4.71 2.14 ;
        RECT 5.275 2.08 5.565 2.14 ;
        RECT 6.135 2.08 6.425 2.14 ;
        RECT 6.99 2.08 7.28 2.14 ;
        RECT 7.84 2.08 8.13 2.14 ;
        RECT 8.72 2.08 9.01 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.085 0.085 0.39 0.595 ;
      RECT 0.595 0.265 0.82 1.075 ;
      RECT 0.595 1.075 7.69 1.325 ;
      RECT 0.595 1.325 0.785 2.465 ;
      RECT 0.99 0.085 1.25 0.61 ;
      RECT 1.43 0.265 1.68 1.075 ;
      RECT 1.455 1.325 1.645 2.46 ;
      RECT 1.85 0.085 2.11 0.645 ;
      RECT 2.71 0.085 2.97 0.565 ;
      RECT 3.57 0.085 3.83 0.565 ;
      RECT 4.43 0.085 4.675 0.565 ;
      RECT 5.29 0.085 5.535 0.565 ;
      RECT 6.145 0.085 6.395 0.565 ;
      RECT 7.005 0.085 7.255 0.565 ;
      RECT 7.865 0.085 8.125 0.565 ;
      RECT 8.725 0.085 9.025 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.345 1.305 0.735 ;
        RECT 1.01 0.735 2.66 0.905 ;
        RECT 1.025 1.835 2.165 1.965 ;
        RECT 1.025 1.965 1.39 1.97 ;
        RECT 1.025 1.97 1.385 1.975 ;
        RECT 1.025 1.975 1.37 1.98 ;
        RECT 1.025 1.98 1.33 2 ;
        RECT 1.025 2 1.325 2.005 ;
        RECT 1.025 2.005 1.265 2.465 ;
        RECT 1.185 1.825 2.165 1.835 ;
        RECT 1.195 1.82 2.165 1.825 ;
        RECT 1.205 1.815 2.165 1.82 ;
        RECT 1.215 1.805 2.165 1.815 ;
        RECT 1.245 1.785 2.165 1.805 ;
        RECT 1.27 1.75 2.165 1.785 ;
        RECT 1.905 0.345 2.165 0.735 ;
        RECT 1.905 1.415 2.66 1.585 ;
        RECT 1.905 1.585 2.165 1.75 ;
        RECT 1.935 1.965 2.165 2.465 ;
        RECT 2.255 0.905 2.66 1.415 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.835 0.855 2.465 ;
      LAYER mcon ;
        RECT 0.61 2.125 0.78 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.435 2.14 1.765 2.465 ;
        RECT 2.335 1.765 2.62 2.465 ;
      LAYER mcon ;
        RECT 1.495 2.14 1.665 2.31 ;
        RECT 2.375 2.125 2.545 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 2.69 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
        RECT 1.435 2.08 1.725 2.14 ;
        RECT 2.315 2.08 2.605 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.255 0.385 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.115 1.665 ;
      RECT 0.085 1.665 0.355 2.465 ;
      RECT 0.555 0.085 0.83 0.565 ;
      RECT 0.945 1.075 2.085 1.245 ;
      RECT 0.945 1.245 1.115 1.495 ;
      RECT 1.475 0.085 1.73 0.565 ;
      RECT 2.335 0.085 2.615 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.76 ;
        RECT 0.085 0.76 0.255 1.56 ;
        RECT 0.085 1.56 0.355 2.465 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.875 0.855 2.465 ;
      LAYER mcon ;
        RECT 0.61 2.125 0.78 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065 -0.085 1.235 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.425 1.06 0.71 1.39 ;
      RECT 0.525 0.085 0.855 0.465 ;
      RECT 0.54 0.635 1.205 0.805 ;
      RECT 0.54 0.805 0.71 1.06 ;
      RECT 0.54 1.39 0.71 1.535 ;
      RECT 0.54 1.535 1.205 1.705 ;
      RECT 1.035 0.255 1.205 0.635 ;
      RECT 1.035 1.705 1.205 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_1
MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.495 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.497000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.77 0.285 3.095 0.615 ;
        RECT 2.77 1.625 3.095 2.46 ;
        RECT 2.865 0.615 3.095 0.765 ;
        RECT 2.865 0.765 3.595 1.275 ;
        RECT 2.865 1.275 3.095 1.625 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.095 0.305 0.345 0.64 ;
      RECT 0.095 0.64 0.84 0.81 ;
      RECT 0.095 1.785 0.835 1.955 ;
      RECT 0.095 1.955 0.345 2.465 ;
      RECT 0.575 0.085 0.905 0.47 ;
      RECT 0.575 2.125 0.905 2.635 ;
      RECT 0.665 0.81 0.84 0.995 ;
      RECT 0.665 0.995 1.035 1.325 ;
      RECT 0.665 1.325 1.005 1.75 ;
      RECT 0.665 1.75 0.835 1.785 ;
      RECT 1.095 0.255 1.425 0.78 ;
      RECT 1.175 1.425 1.44 2.465 ;
      RECT 1.205 0.78 1.425 0.995 ;
      RECT 1.205 0.995 2.165 1.325 ;
      RECT 1.205 1.325 1.44 1.425 ;
      RECT 1.615 0.255 1.945 0.635 ;
      RECT 1.615 0.635 2.595 0.805 ;
      RECT 1.695 1.5 2.595 1.745 ;
      RECT 1.695 1.745 1.945 2.465 ;
      RECT 2.135 0.085 2.465 0.465 ;
      RECT 2.135 1.915 2.465 2.635 ;
      RECT 2.335 0.805 2.595 1.5 ;
      RECT 3.265 0.085 3.595 0.55 ;
      RECT 3.265 1.635 3.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2
MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.485 1.32 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.702900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015 0.255 3.595 0.64 ;
        RECT 3.035 1.565 3.595 2.465 ;
        RECT 3.23 0.64 3.595 1.565 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.255 0.41 0.735 ;
      RECT 0.085 0.735 1.005 0.905 ;
      RECT 0.085 1.49 1.005 1.66 ;
      RECT 0.085 1.66 0.43 2.465 ;
      RECT 0.58 0.085 0.91 0.565 ;
      RECT 0.6 1.83 0.925 2.635 ;
      RECT 0.655 0.905 1.005 1.025 ;
      RECT 0.655 1.025 1.105 1.295 ;
      RECT 0.655 1.295 1.005 1.49 ;
      RECT 1.175 0.255 1.645 0.855 ;
      RECT 1.195 1.79 1.645 2.465 ;
      RECT 1.47 0.855 1.645 1.075 ;
      RECT 1.47 1.075 2.42 1.25 ;
      RECT 1.47 1.25 1.645 1.79 ;
      RECT 1.815 0.255 2.065 0.735 ;
      RECT 1.815 0.735 2.765 0.905 ;
      RECT 1.815 1.495 2.765 1.665 ;
      RECT 1.815 1.665 2.065 2.465 ;
      RECT 2.235 1.835 2.845 2.635 ;
      RECT 2.24 0.085 2.845 0.565 ;
      RECT 2.595 0.905 2.765 0.99 ;
      RECT 2.595 0.99 3.05 1.325 ;
      RECT 2.595 1.325 2.765 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1
MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputisolatch_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 0.765 2.125 1.095 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.69 0.415 4.975 0.745 ;
        RECT 4.69 1.67 4.975 2.455 ;
        RECT 4.805 0.745 4.975 1.67 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.145500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.13 ;
      RECT 0.61 1.13 0.81 1.46 ;
      RECT 0.61 1.46 0.78 1.795 ;
      RECT 0.98 0.74 1.185 0.91 ;
      RECT 0.98 0.91 1.15 1.825 ;
      RECT 0.98 1.825 1.185 1.915 ;
      RECT 0.98 1.915 2.845 1.965 ;
      RECT 1.015 0.345 1.185 0.74 ;
      RECT 1.015 1.965 2.845 2.085 ;
      RECT 1.015 2.085 1.185 2.465 ;
      RECT 1.32 1.24 1.49 1.525 ;
      RECT 1.32 1.525 2.335 1.695 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.255 1.85 2.635 ;
      RECT 2.05 1.355 2.335 1.525 ;
      RECT 2.295 0.705 2.675 1.035 ;
      RECT 2.31 2.255 3.185 2.425 ;
      RECT 2.38 0.365 3.04 0.535 ;
      RECT 2.505 1.035 2.675 1.575 ;
      RECT 2.505 1.575 2.845 1.915 ;
      RECT 2.87 0.535 3.04 0.995 ;
      RECT 2.87 0.995 3.78 1.165 ;
      RECT 3.015 1.165 3.78 1.325 ;
      RECT 3.015 1.325 3.185 2.255 ;
      RECT 3.265 0.085 3.595 0.53 ;
      RECT 3.355 2.135 3.525 2.635 ;
      RECT 3.42 1.535 4.125 1.865 ;
      RECT 3.835 0.415 4.125 0.745 ;
      RECT 3.835 1.865 4.125 2.435 ;
      RECT 3.95 0.745 4.125 1.535 ;
      RECT 4.295 0.085 4.465 0.715 ;
      RECT 4.295 1.57 4.465 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1
MACRO sky130_fd_sc_hd__o2111a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.83 1.005 4.515 1.315 ;
        RECT 4.31 1.315 4.515 2.355 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.3 0.995 3.66 1.325 ;
        RECT 3.37 1.325 3.66 2.37 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 1.075 3.1 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.255 2.39 1.615 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 1.835 1.615 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.855 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.135 0.085 0.345 0.885 ;
      RECT 0.135 1.495 0.345 2.635 ;
      RECT 1.03 0.715 1.805 0.885 ;
      RECT 1.03 0.885 1.305 1.785 ;
      RECT 1.03 1.785 3.195 2.025 ;
      RECT 1.035 0.085 1.285 0.545 ;
      RECT 1.035 2.195 1.655 2.635 ;
      RECT 1.475 0.255 1.805 0.715 ;
      RECT 1.86 2.025 2.14 2.465 ;
      RECT 2.325 2.255 2.655 2.635 ;
      RECT 2.865 0.255 3.195 0.625 ;
      RECT 2.865 0.625 4.215 0.825 ;
      RECT 2.865 2.025 3.195 2.465 ;
      RECT 3.385 0.085 3.715 0.455 ;
      RECT 3.885 0.255 4.215 0.625 ;
      RECT 3.885 1.495 4.14 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__o2111a_2
MACRO sky130_fd_sc_hd__o2111a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.075 4.035 1.66 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.075 3.535 1.325 ;
        RECT 3.35 1.325 3.535 2.415 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.39 2.69 0.995 ;
        RECT 2.445 0.995 2.705 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.39 2.195 1.325 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265 1.075 1.745 1.325 ;
        RECT 1.535 0.39 1.745 1.075 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.255 0.355 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.525 0.995 0.865 1.325 ;
      RECT 0.525 1.835 1.335 2.635 ;
      RECT 0.535 0.085 0.845 0.565 ;
      RECT 0.695 0.735 1.365 0.905 ;
      RECT 0.695 0.905 0.865 0.995 ;
      RECT 0.695 1.325 0.865 1.495 ;
      RECT 0.695 1.495 3.18 1.665 ;
      RECT 1.025 0.255 1.365 0.735 ;
      RECT 1.505 1.665 1.835 2.465 ;
      RECT 2.02 1.835 2.76 2.635 ;
      RECT 2.87 0.255 3.16 0.705 ;
      RECT 2.87 0.705 4.055 0.875 ;
      RECT 2.93 1.665 3.18 2.465 ;
      RECT 3.33 0.085 3.62 0.535 ;
      RECT 3.73 1.835 4.055 2.635 ;
      RECT 3.79 0.255 4.055 0.705 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o2111a_1
MACRO sky130_fd_sc_hd__o2111a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.89 1.075 4.485 1.245 ;
        RECT 4.13 1.245 4.485 1.32 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135 1.075 3.6 1.245 ;
        RECT 3.145 1.245 3.6 1.32 ;
        RECT 3.305 1.32 3.6 1.49 ;
        RECT 3.305 1.49 4.825 1.66 ;
        RECT 4.655 1.075 4.985 1.32 ;
        RECT 4.655 1.32 4.825 1.49 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.215 1.32 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.15 0.995 1.395 1.49 ;
        RECT 1.15 1.49 2.66 1.66 ;
        RECT 2.445 1.08 2.82 1.32 ;
        RECT 2.445 1.32 2.66 1.49 ;
        RECT 2.49 1.075 2.82 1.08 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 0.34 1.655 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.962500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.65 0.255 5.875 0.695 ;
        RECT 5.65 0.695 7.275 0.865 ;
        RECT 5.755 1.495 7.275 1.665 ;
        RECT 5.755 1.665 5.925 2.465 ;
        RECT 6.545 0.255 6.745 0.695 ;
        RECT 6.585 1.665 6.775 2.465 ;
        RECT 7.005 0.865 7.275 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.09 1.835 5.55 2 ;
      RECT 0.09 2 5.065 2.005 ;
      RECT 0.09 2.005 0.345 2.465 ;
      RECT 0.1 0.255 2.94 0.485 ;
      RECT 0.1 0.485 0.345 0.825 ;
      RECT 0.515 0.655 0.86 1.83 ;
      RECT 0.515 1.83 5.55 1.835 ;
      RECT 0.515 2.175 0.845 2.635 ;
      RECT 1.015 2.005 1.23 2.465 ;
      RECT 1.4 2.175 1.625 2.635 ;
      RECT 1.72 0.655 4.795 0.885 ;
      RECT 1.795 2.005 2.025 2.465 ;
      RECT 2.195 2.175 2.525 2.635 ;
      RECT 2.695 2.005 3.285 2.465 ;
      RECT 3.11 0.085 3.44 0.485 ;
      RECT 3.61 0.255 3.825 0.655 ;
      RECT 3.805 2.18 4.135 2.635 ;
      RECT 3.995 0.085 4.365 0.485 ;
      RECT 4.535 0.255 4.795 0.655 ;
      RECT 4.775 2.005 5.065 2.465 ;
      RECT 5.035 0.085 5.3 0.545 ;
      RECT 5.245 2.17 5.585 2.635 ;
      RECT 5.38 1.075 6.76 1.32 ;
      RECT 5.38 1.32 5.55 1.83 ;
      RECT 6.075 0.085 6.375 0.525 ;
      RECT 6.095 1.835 6.415 2.635 ;
      RECT 6.915 0.085 7.275 0.525 ;
      RECT 6.945 1.835 7.27 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__o2111a_4
MACRO sky130_fd_sc_hd__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.275 12.335 0.825 ;
        RECT 11.995 1.495 12.335 2.45 ;
        RECT 12.145 0.825 12.335 1.495 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
      LAYER mcon ;
        RECT 0.605 1.105 0.775 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
      LAYER mcon ;
        RECT 2.445 1.105 2.615 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
      LAYER mcon ;
        RECT 8.94 1.445 9.11 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.61 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.42 0.085 ;
      RECT 0 2.635 12.42 2.805 ;
      RECT 0.085 0.085 0.7 0.595 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.515 2.195 0.785 2.635 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.825 0.085 2.09 0.545 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 2.69 0.085 3.1 0.555 ;
      RECT 2.69 2.14 2.985 2.635 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.595 2.275 3.925 2.635 ;
      RECT 3.625 0.085 3.955 0.545 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.61 0.085 6.095 0.465 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 5.945 2.275 6.33 2.635 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 6.705 0.085 7.715 0.805 ;
      RECT 7.06 2.125 8.015 2.635 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.16 2.235 9.49 2.635 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.115 0.085 10.365 0.545 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.155 2.235 10.485 2.635 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
      RECT 11.515 0.085 11.825 0.825 ;
      RECT 11.515 1.79 11.825 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.48 1.105 8.65 1.275 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_1
MACRO sky130_fd_sc_hd__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035 0.255 12.365 0.825 ;
        RECT 12.035 1.495 12.365 2.45 ;
        RECT 12.145 0.825 12.365 1.495 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
      LAYER mcon ;
        RECT 0.605 1.105 0.775 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
      LAYER mcon ;
        RECT 2.445 1.105 2.615 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
      LAYER mcon ;
        RECT 8.94 1.445 9.11 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 13.07 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.88 0.085 ;
      RECT 0 2.635 12.88 2.805 ;
      RECT 0.085 0.085 0.7 0.595 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.515 2.195 0.785 2.635 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.825 0.085 2.09 0.545 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 2.69 0.085 3.1 0.555 ;
      RECT 2.69 2.14 2.985 2.635 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.595 2.275 3.925 2.635 ;
      RECT 3.625 0.085 3.955 0.545 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.61 0.085 6.095 0.465 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 5.945 2.275 6.33 2.635 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 6.705 0.085 7.715 0.805 ;
      RECT 7.06 2.125 8.015 2.635 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.16 2.235 9.49 2.635 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.115 0.085 10.365 0.545 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.155 2.235 10.485 2.635 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
      RECT 11.57 0.085 11.865 0.825 ;
      RECT 11.57 1.79 11.82 2.635 ;
      RECT 12.535 0.085 12.795 0.885 ;
      RECT 12.535 1.495 12.795 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.48 1.105 8.65 1.275 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_2
MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.48 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.04 0.275 12.37 0.825 ;
        RECT 12.04 1.495 12.37 2.45 ;
        RECT 12.145 0.825 12.37 1.055 ;
        RECT 12.145 1.055 13.21 1.325 ;
        RECT 12.145 1.325 12.37 1.495 ;
        RECT 12.88 0.255 13.21 1.055 ;
        RECT 12.88 1.325 13.21 2.465 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
      LAYER mcon ;
        RECT 0.605 1.105 0.775 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
      LAYER mcon ;
        RECT 2.445 1.105 2.615 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
      LAYER mcon ;
        RECT 8.94 1.445 9.11 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.8 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 13.99 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.8 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 13.8 0.085 ;
      RECT 0 2.635 13.8 2.805 ;
      RECT 0.085 0.085 0.7 0.595 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.515 2.195 0.785 2.635 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.825 0.085 2.09 0.545 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 2.69 0.085 3.1 0.555 ;
      RECT 2.69 2.14 2.985 2.635 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.595 2.275 3.925 2.635 ;
      RECT 3.625 0.085 3.955 0.545 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.61 0.085 6.095 0.465 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 5.945 2.275 6.33 2.635 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 6.705 0.085 7.715 0.805 ;
      RECT 7.06 2.125 8.015 2.635 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.16 2.235 9.49 2.635 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.115 0.085 10.365 0.545 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.155 2.235 10.485 2.635 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
      RECT 11.515 0.085 11.87 0.825 ;
      RECT 11.515 1.495 11.87 2.635 ;
      RECT 12.54 0.085 12.71 0.885 ;
      RECT 12.54 1.495 12.71 2.635 ;
      RECT 13.38 0.085 13.715 0.885 ;
      RECT 13.38 1.495 13.715 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.48 1.105 8.65 1.275 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_4
MACRO sky130_fd_sc_hd__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.33 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 3.1 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.36 1.075 4.45 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.62 1.075 5.43 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 1.785 0.825 ;
        RECT 1.455 1.445 4.865 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 1.55 0.825 1.785 1.445 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 3.605 1.665 3.935 2.465 ;
        RECT 4.535 1.665 4.865 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.09 0.255 0.345 0.635 ;
      RECT 0.09 0.635 0.67 0.805 ;
      RECT 0.09 1.915 0.67 2.085 ;
      RECT 0.09 2.085 0.345 2.465 ;
      RECT 0.5 0.805 0.67 1.075 ;
      RECT 0.5 1.075 1.38 1.245 ;
      RECT 0.5 1.245 0.67 1.915 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.255 1.285 2.635 ;
      RECT 1.035 0.255 2.125 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 1.035 1.445 1.285 2.255 ;
      RECT 1.955 0.465 2.125 0.635 ;
      RECT 1.955 0.635 3.045 0.905 ;
      RECT 1.955 1.835 2.125 2.635 ;
      RECT 2.295 0.255 3.985 0.465 ;
      RECT 2.795 1.835 3.435 2.635 ;
      RECT 3.235 0.635 4.455 0.715 ;
      RECT 3.235 0.715 5.34 0.905 ;
      RECT 4.105 1.835 4.365 2.635 ;
      RECT 4.155 0.255 4.415 0.615 ;
      RECT 4.155 0.615 4.455 0.635 ;
      RECT 4.665 0.085 4.835 0.545 ;
      RECT 5.005 0.255 5.34 0.715 ;
      RECT 5.035 1.495 5.43 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__nand4b_2
MACRO sky130_fd_sc_hd__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.765 2.185 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 0.765 1.755 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.887500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.13 1.495 3.135 1.665 ;
        RECT 1.13 1.665 1.46 2.465 ;
        RECT 2.085 1.665 2.415 2.465 ;
        RECT 2.695 0.255 3.135 0.825 ;
        RECT 2.925 0.825 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.445 0.475 0.655 ;
      RECT 0.085 0.655 1.335 0.825 ;
      RECT 0.085 0.825 0.255 1.595 ;
      RECT 0.085 1.595 0.51 1.925 ;
      RECT 0.655 0.085 0.985 0.485 ;
      RECT 0.71 1.495 0.96 2.635 ;
      RECT 1.155 0.425 2.525 0.595 ;
      RECT 1.155 0.595 1.335 0.655 ;
      RECT 1.63 1.835 1.915 2.635 ;
      RECT 2.355 0.595 2.525 0.995 ;
      RECT 2.355 0.995 2.755 1.325 ;
      RECT 2.705 1.835 2.92 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__nand4b_1
MACRO sky130_fd_sc_hd__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.93 1.075 4.59 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 6.51 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.015 1.075 8.655 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.64 0.905 ;
        RECT 1.455 1.445 8.185 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 2.375 0.905 2.64 1.445 ;
        RECT 3.135 1.665 3.465 2.465 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
        RECT 7.015 1.665 7.345 2.465 ;
        RECT 7.855 1.665 8.185 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 0.805 0.905 ;
      RECT 0.09 1.495 0.805 1.665 ;
      RECT 0.09 1.665 0.425 2.465 ;
      RECT 0.595 0.085 0.845 0.545 ;
      RECT 0.595 1.835 1.285 2.635 ;
      RECT 0.61 0.905 0.805 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.805 1.495 ;
      RECT 0.995 1.495 1.285 1.835 ;
      RECT 1.035 0.255 4.725 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 1.955 1.835 2.125 2.635 ;
      RECT 2.795 1.835 2.965 2.635 ;
      RECT 3.135 0.635 6.505 0.905 ;
      RECT 3.635 1.835 3.805 2.635 ;
      RECT 4.475 1.835 5.165 2.635 ;
      RECT 4.915 0.255 6.925 0.465 ;
      RECT 5.835 1.835 6.005 2.635 ;
      RECT 6.675 0.465 6.925 0.735 ;
      RECT 6.675 0.735 8.61 0.905 ;
      RECT 6.675 1.835 6.845 2.635 ;
      RECT 7.095 0.085 7.265 0.545 ;
      RECT 7.435 0.255 7.765 0.735 ;
      RECT 7.515 1.835 7.685 2.635 ;
      RECT 7.935 0.085 8.105 0.545 ;
      RECT 8.275 0.255 8.61 0.735 ;
      RECT 8.355 1.445 8.61 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
  END
END sky130_fd_sc_hd__nand4b_4
MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.32 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 2.125 2.67 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.55 1.075 3.55 1.275 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.435 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.675 1.25 0.68 ;
        RECT 0.935 0.68 1.245 0.79 ;
        RECT 0.935 0.79 1.105 1.495 ;
        RECT 0.935 1.495 1.25 1.825 ;
        RECT 0.97 0.26 1.25 0.675 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.325 0.35 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.605 0.765 1.89 ;
      RECT 0.51 1.89 0.765 1.995 ;
      RECT 0.51 1.995 1.715 2.165 ;
      RECT 0.515 2.335 0.845 2.635 ;
      RECT 0.595 0.905 0.765 1.605 ;
      RECT 0.63 0.085 0.8 0.565 ;
      RECT 1.29 0.995 1.585 1.325 ;
      RECT 1.415 0.735 3.055 0.905 ;
      RECT 1.415 0.905 1.585 0.995 ;
      RECT 1.415 1.325 1.585 1.355 ;
      RECT 1.415 1.355 1.6 1.37 ;
      RECT 1.415 1.37 1.61 1.38 ;
      RECT 1.415 1.38 1.62 1.39 ;
      RECT 1.415 1.39 1.625 1.4 ;
      RECT 1.415 1.4 1.63 1.41 ;
      RECT 1.415 1.41 1.645 1.42 ;
      RECT 1.415 1.42 1.655 1.425 ;
      RECT 1.415 1.425 1.665 1.445 ;
      RECT 1.415 1.445 3.56 1.45 ;
      RECT 1.42 1.45 3.56 1.615 ;
      RECT 1.435 0.085 1.815 0.485 ;
      RECT 1.44 1.785 3.03 1.955 ;
      RECT 1.44 1.955 1.715 1.995 ;
      RECT 1.48 2.335 1.815 2.635 ;
      RECT 1.985 0.305 2.155 0.735 ;
      RECT 2.385 0.085 2.715 0.485 ;
      RECT 2.86 1.955 3.03 2.215 ;
      RECT 2.86 2.215 3.345 2.385 ;
      RECT 2.885 0.305 3.055 0.735 ;
      RECT 3.225 0.085 3.555 0.585 ;
      RECT 3.225 1.615 3.56 1.815 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__or4b_2
MACRO sky130_fd_sc_hd__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755 0.995 2.925 1.445 ;
        RECT 2.755 1.445 3.19 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 0.995 2.525 1.45 ;
        RECT 2.335 1.45 2.525 1.785 ;
        RECT 2.335 1.785 2.635 2.375 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 0.995 1.965 1.62 ;
        RECT 1.795 1.62 2.155 2.375 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.995 0.445 1.955 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.455 4.965 1.625 ;
        RECT 3.395 1.625 3.645 2.465 ;
        RECT 3.435 0.255 3.685 0.725 ;
        RECT 3.435 0.725 4.965 0.905 ;
        RECT 4.195 0.255 4.525 0.725 ;
        RECT 4.235 1.625 4.485 2.465 ;
        RECT 4.725 0.905 4.965 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.085 0.345 0.825 ;
      RECT 0.085 2.135 0.365 2.635 ;
      RECT 0.595 0.435 0.785 0.905 ;
      RECT 0.595 2.065 0.785 2.455 ;
      RECT 0.615 0.905 0.785 0.995 ;
      RECT 0.615 0.995 1.215 1.325 ;
      RECT 0.615 1.325 0.785 2.065 ;
      RECT 1.035 0.085 1.285 0.585 ;
      RECT 1.035 1.575 1.625 1.745 ;
      RECT 1.035 1.745 1.365 2.45 ;
      RECT 1.455 0.655 3.265 0.825 ;
      RECT 1.455 0.825 1.625 1.575 ;
      RECT 1.615 0.305 1.785 0.655 ;
      RECT 1.985 0.085 2.315 0.485 ;
      RECT 2.485 0.305 2.655 0.655 ;
      RECT 2.875 0.085 3.255 0.485 ;
      RECT 2.92 1.795 3.17 2.635 ;
      RECT 3.095 0.825 3.265 1.075 ;
      RECT 3.095 1.075 4.555 1.245 ;
      RECT 3.815 1.795 4.065 2.635 ;
      RECT 3.855 0.085 4.025 0.555 ;
      RECT 4.655 1.795 4.905 2.635 ;
      RECT 4.695 0.085 4.865 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__or4b_4
MACRO sky130_fd_sc_hd__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.43 0.995 2.81 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 2.125 2.66 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.995 2.26 1.615 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.425 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.415 3.595 0.76 ;
        RECT 3.32 1.495 3.595 2.465 ;
        RECT 3.425 0.76 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.085 0.425 0.585 ;
      RECT 0.085 1.56 0.425 2.635 ;
      RECT 0.595 0.305 0.84 0.995 ;
      RECT 0.595 0.995 1.25 1.325 ;
      RECT 0.595 1.325 0.835 1.92 ;
      RECT 1.03 1.495 1.35 1.785 ;
      RECT 1.03 1.785 2.66 1.955 ;
      RECT 1.035 0.085 1.365 0.585 ;
      RECT 1.565 0.305 1.735 0.655 ;
      RECT 1.565 0.655 3.15 0.825 ;
      RECT 1.91 0.085 2.24 0.485 ;
      RECT 2.41 0.305 2.58 0.655 ;
      RECT 2.49 1.495 3.15 1.665 ;
      RECT 2.49 1.665 2.66 1.785 ;
      RECT 2.75 0.085 3.13 0.485 ;
      RECT 2.83 1.835 3.11 2.635 ;
      RECT 2.98 0.825 3.15 0.995 ;
      RECT 2.98 0.995 3.255 1.325 ;
      RECT 2.98 1.325 3.15 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__or4b_1
MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.79 1.055 4.045 1.225 ;
        RECT 3.82 1.225 4.045 1.675 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.31 1.005 2.615 1.395 ;
        RECT 2.31 1.395 3.595 1.675 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635 0.315 4.965 0.825 ;
        RECT 4.715 1.545 4.965 2.415 ;
        RECT 4.79 0.825 4.965 1.545 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.315 0.885 0.825 ;
        RECT 0.555 0.825 0.78 1.565 ;
        RECT 0.555 1.565 0.885 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.135 0.085 0.375 0.885 ;
      RECT 0.135 1.495 0.375 2.635 ;
      RECT 0.95 1.075 1.59 1.245 ;
      RECT 1.055 0.085 1.25 0.885 ;
      RECT 1.055 1.515 1.25 2.635 ;
      RECT 1.42 0.345 1.745 0.675 ;
      RECT 1.42 0.675 1.59 1.075 ;
      RECT 1.42 1.245 1.59 2.205 ;
      RECT 1.42 2.205 2.22 2.375 ;
      RECT 1.76 0.995 1.93 1.855 ;
      RECT 1.76 1.855 4.465 2.025 ;
      RECT 1.995 0.345 2.165 0.635 ;
      RECT 1.995 0.635 3.005 0.805 ;
      RECT 2.335 0.085 2.665 0.465 ;
      RECT 2.835 0.345 3.005 0.635 ;
      RECT 2.85 2.205 3.64 2.635 ;
      RECT 3.46 0.345 3.63 0.715 ;
      RECT 3.46 0.715 4.465 0.885 ;
      RECT 3.81 2.025 3.98 2.355 ;
      RECT 4.215 0.085 4.465 0.545 ;
      RECT 4.215 2.205 4.545 2.635 ;
      RECT 4.295 0.885 4.465 0.995 ;
      RECT 4.295 0.995 4.62 1.325 ;
      RECT 4.295 1.325 4.465 1.855 ;
      RECT 5.145 0.085 5.385 0.885 ;
      RECT 5.145 1.495 5.385 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__ha_2
MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 1.075 4.38 1.245 ;
        RECT 4.21 1.245 4.38 1.505 ;
        RECT 4.21 1.505 6.81 1.675 ;
        RECT 5.625 0.995 5.795 1.505 ;
        RECT 6.58 0.995 7.055 1.325 ;
        RECT 6.58 1.325 6.81 1.505 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.55 0.995 5.455 1.165 ;
        RECT 4.55 1.165 4.72 1.325 ;
        RECT 5.285 0.73 6.315 0.825 ;
        RECT 5.285 0.825 5.535 0.845 ;
        RECT 5.285 0.845 5.495 0.875 ;
        RECT 5.285 0.875 5.455 0.995 ;
        RECT 5.295 0.72 6.315 0.73 ;
        RECT 5.31 0.71 6.315 0.72 ;
        RECT 5.32 0.695 6.315 0.71 ;
        RECT 5.335 0.675 6.315 0.695 ;
        RECT 5.345 0.655 6.315 0.675 ;
        RECT 6.085 0.825 6.315 1.325 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595 0.315 7.845 0.735 ;
        RECT 7.595 0.735 8.685 0.905 ;
        RECT 7.595 1.415 8.685 1.585 ;
        RECT 7.595 1.585 7.765 2.415 ;
        RECT 8.405 0.315 8.685 0.735 ;
        RECT 8.405 0.905 8.685 1.415 ;
        RECT 8.405 1.585 8.685 2.415 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.315 0.845 1.065 ;
        RECT 0.515 1.065 1.55 1.335 ;
        RECT 0.515 1.335 0.845 2.415 ;
        RECT 1.355 0.315 1.685 0.825 ;
        RECT 1.355 0.825 1.55 1.065 ;
        RECT 1.355 1.335 1.55 1.565 ;
        RECT 1.355 1.565 1.685 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.135 0.085 0.345 0.885 ;
      RECT 0.135 1.495 0.345 2.635 ;
      RECT 1.015 0.085 1.185 0.885 ;
      RECT 1.015 1.515 1.185 2.635 ;
      RECT 1.72 1.075 2.75 1.245 ;
      RECT 1.855 0.085 2.095 0.885 ;
      RECT 1.855 1.495 2.365 2.635 ;
      RECT 2.27 0.305 3.385 0.475 ;
      RECT 2.58 0.645 3.045 0.815 ;
      RECT 2.58 0.815 2.75 1.075 ;
      RECT 2.58 1.245 2.75 1.765 ;
      RECT 2.58 1.765 3.7 1.935 ;
      RECT 2.77 1.935 2.94 2.355 ;
      RECT 2.92 0.995 3.09 1.425 ;
      RECT 2.92 1.425 4.04 1.595 ;
      RECT 3.19 2.105 3.36 2.635 ;
      RECT 3.215 0.475 3.385 0.645 ;
      RECT 3.215 0.645 5.115 0.815 ;
      RECT 3.53 1.935 3.7 2.205 ;
      RECT 3.53 2.205 4.33 2.375 ;
      RECT 3.555 0.085 3.91 0.465 ;
      RECT 3.87 1.595 4.04 1.855 ;
      RECT 3.87 1.855 7.395 2.025 ;
      RECT 4.08 0.345 4.25 0.645 ;
      RECT 4.42 0.085 4.75 0.465 ;
      RECT 4.92 0.255 5.19 0.585 ;
      RECT 4.92 0.585 5.115 0.645 ;
      RECT 5.24 2.205 5.57 2.635 ;
      RECT 5.385 0.085 5.715 0.465 ;
      RECT 5.835 2.025 6.005 2.355 ;
      RECT 6.175 0.295 6.875 0.465 ;
      RECT 6.175 2.205 6.505 2.635 ;
      RECT 6.675 2.025 6.845 2.355 ;
      RECT 6.705 0.465 6.875 0.645 ;
      RECT 6.705 0.645 7.395 0.815 ;
      RECT 7.055 0.085 7.385 0.465 ;
      RECT 7.055 2.205 7.385 2.635 ;
      RECT 7.225 0.815 7.395 1.075 ;
      RECT 7.225 1.075 8.225 1.245 ;
      RECT 7.225 1.245 7.395 1.855 ;
      RECT 7.935 1.755 8.225 2.635 ;
      RECT 8.015 0.085 8.225 0.565 ;
      RECT 8.855 0.085 9.065 0.885 ;
      RECT 8.855 1.495 9.065 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
  END
END sky130_fd_sc_hd__ha_4
MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.315 3.585 1.485 ;
        RECT 3.36 1.055 3.585 1.315 ;
        RECT 3.36 1.485 3.585 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.85 1.345 2.155 1.655 ;
        RECT 1.85 1.655 3.165 1.825 ;
        RECT 1.85 1.825 2.155 2.375 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.315 4.515 0.825 ;
        RECT 4.175 1.565 4.515 2.415 ;
        RECT 4.33 0.825 4.515 1.565 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.315 0.425 0.825 ;
        RECT 0.09 0.825 0.32 1.565 ;
        RECT 0.09 1.565 0.425 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.49 1.075 1.13 1.245 ;
      RECT 0.595 0.085 0.79 0.885 ;
      RECT 0.595 1.515 0.79 2.275 ;
      RECT 0.595 2.275 1.26 2.635 ;
      RECT 0.96 0.345 1.285 0.675 ;
      RECT 0.96 0.675 1.13 1.075 ;
      RECT 0.96 1.245 1.13 1.935 ;
      RECT 0.96 1.935 1.68 2.105 ;
      RECT 1.3 0.975 3.17 1.145 ;
      RECT 1.3 1.145 1.47 1.325 ;
      RECT 1.51 2.105 1.68 2.355 ;
      RECT 1.535 0.345 1.705 0.635 ;
      RECT 1.535 0.635 2.545 0.805 ;
      RECT 1.875 0.085 2.205 0.465 ;
      RECT 2.375 0.345 2.545 0.635 ;
      RECT 2.45 2.275 3.12 2.635 ;
      RECT 3 0.345 3.17 0.715 ;
      RECT 3 0.715 4.005 0.885 ;
      RECT 3 0.885 3.17 0.975 ;
      RECT 3.35 1.785 4.005 1.955 ;
      RECT 3.35 1.955 3.52 2.355 ;
      RECT 3.755 0.085 4.005 0.545 ;
      RECT 3.755 2.125 4.005 2.635 ;
      RECT 3.835 0.885 4.005 0.995 ;
      RECT 3.835 0.995 4.16 1.325 ;
      RECT 3.835 1.325 4.005 1.785 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__ha_1
MACRO sky130_fd_sc_hd__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.945 0.265 9.2 0.795 ;
        RECT 8.945 1.655 9.2 2.325 ;
        RECT 9.02 0.795 9.2 1.655 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
      LAYER mcon ;
        RECT 3.85 0.765 4.02 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.68 0.735 7.34 1.005 ;
        RECT 6.68 1.005 7.01 1.065 ;
      LAYER mcon ;
        RECT 7.11 0.765 7.28 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.79 0.735 4.08 0.78 ;
        RECT 3.79 0.78 7.34 0.92 ;
        RECT 3.79 0.92 4.08 0.965 ;
        RECT 7.05 0.735 7.34 0.78 ;
        RECT 7.05 0.92 7.34 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.73 2.085 ;
      RECT 3.43 2.255 3.81 2.635 ;
      RECT 3.61 0.085 4.02 0.525 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.73 1.065 ;
      RECT 4.33 2.255 4.66 2.635 ;
      RECT 4.54 1.065 4.73 1.835 ;
      RECT 4.76 0.085 5.08 0.545 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.42 1.965 ;
      RECT 5.13 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.49 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.8 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.85 1.745 ;
      RECT 5.94 2.255 6.36 2.635 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.56 2.085 6.8 2.375 ;
      RECT 6.69 0.085 7.35 0.565 ;
      RECT 7.03 1.945 7.36 2.635 ;
      RECT 7.16 1.175 7.49 1.235 ;
      RECT 7.53 0.35 7.85 0.68 ;
      RECT 7.53 1.745 7.85 1.765 ;
      RECT 7.53 1.765 7.7 2.375 ;
      RECT 7.66 0.68 7.85 1.575 ;
      RECT 7.97 1.915 8.3 2.425 ;
      RECT 8.05 0.345 8.3 0.995 ;
      RECT 8.05 0.995 8.85 1.325 ;
      RECT 8.05 1.325 8.3 1.915 ;
      RECT 8.48 0.085 8.765 0.545 ;
      RECT 8.48 1.835 8.765 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 0.765 3.1 0.935 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.25 1.105 5.42 1.275 ;
      RECT 5.25 1.785 5.42 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 5.48 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 3.16 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 0.735 3.16 0.78 ;
      RECT 2.87 0.92 3.16 0.965 ;
      RECT 2.945 0.965 3.16 1.12 ;
      RECT 2.945 1.12 5.48 1.26 ;
      RECT 5.19 1.075 5.48 1.12 ;
      RECT 5.19 1.26 5.48 1.305 ;
      RECT 5.19 1.755 5.48 1.8 ;
      RECT 5.19 1.94 5.48 1.985 ;
  END
END sky130_fd_sc_hd__dfstp_1
MACRO sky130_fd_sc_hd__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.320000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.925 0.265 9.17 0.715 ;
        RECT 8.925 0.715 10.955 0.885 ;
        RECT 8.925 1.47 10.955 1.64 ;
        RECT 8.925 1.64 9.17 2.465 ;
        RECT 9.765 0.265 9.935 0.715 ;
        RECT 9.765 1.64 9.935 2.465 ;
        RECT 10.605 0.265 10.955 0.715 ;
        RECT 10.605 1.64 10.955 2.465 ;
        RECT 10.725 0.885 10.955 1.47 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
      LAYER mcon ;
        RECT 3.825 0.765 3.995 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
      LAYER mcon ;
        RECT 7.045 0.765 7.215 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.43 2.255 3.81 2.635 ;
      RECT 3.61 0.085 4.02 0.525 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.33 2.255 4.66 2.635 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.74 0.085 5.08 0.545 ;
      RECT 4.88 0.725 6.15 0.895 ;
      RECT 4.88 0.895 5.05 1.655 ;
      RECT 4.88 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.74 2.415 ;
      RECT 5.22 1.065 5.4 1.475 ;
      RECT 5.57 1.235 7.47 1.405 ;
      RECT 5.57 1.405 5.74 1.915 ;
      RECT 5.57 1.915 6.78 2.085 ;
      RECT 5.57 2.085 5.74 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.91 1.575 7.85 1.745 ;
      RECT 5.92 2.255 6.34 2.635 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 6.67 0.085 7.33 0.565 ;
      RECT 7.01 1.945 7.34 2.635 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.85 0.68 ;
      RECT 7.51 1.745 7.85 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.85 1.575 ;
      RECT 7.95 1.915 8.28 2.425 ;
      RECT 8.03 0.345 8.28 1.055 ;
      RECT 8.03 1.055 10.555 1.275 ;
      RECT 8.03 1.275 8.28 1.915 ;
      RECT 8.46 0.085 8.745 0.545 ;
      RECT 8.46 1.835 8.745 2.635 ;
      RECT 9.34 0.085 9.595 0.545 ;
      RECT 9.34 1.81 9.595 2.635 ;
      RECT 10.105 0.085 10.435 0.545 ;
      RECT 10.105 1.81 10.435 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.615 1.785 0.785 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.225 1.105 5.395 1.275 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.555 1.755 0.845 1.8 ;
      RECT 0.555 1.8 5.435 1.94 ;
      RECT 0.555 1.94 0.845 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.455 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.165 1.075 5.455 1.12 ;
      RECT 5.165 1.26 5.455 1.305 ;
  END
END sky130_fd_sc_hd__dfstp_4
MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.81 1.495 9.575 1.615 ;
        RECT 8.81 1.615 9.14 2.46 ;
        RECT 8.89 0.265 9.135 0.765 ;
        RECT 8.89 0.765 9.575 0.825 ;
        RECT 8.975 0.825 9.575 0.855 ;
        RECT 8.975 1.445 9.575 1.495 ;
        RECT 8.99 0.855 9.575 0.895 ;
        RECT 9.02 0.895 9.575 1.445 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
      LAYER mcon ;
        RECT 3.825 0.765 3.995 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.34 1.005 ;
        RECT 6.66 1.005 7.01 1.065 ;
      LAYER mcon ;
        RECT 7.045 0.765 7.215 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.835 0.805 ;
      RECT 0.085 1.795 0.835 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.005 0.565 1.235 2.045 ;
      RECT 1.015 0.345 1.235 0.565 ;
      RECT 1.015 2.045 1.235 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.455 0.085 1.785 0.465 ;
      RECT 1.455 2.135 1.785 2.635 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.43 2.255 3.81 2.635 ;
      RECT 3.61 0.085 4.02 0.525 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.33 2.255 4.66 2.635 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.76 0.085 5.08 0.545 ;
      RECT 4.88 0.725 6.15 0.895 ;
      RECT 4.88 0.895 5.05 1.655 ;
      RECT 4.88 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.74 2.415 ;
      RECT 5.22 1.065 5.4 1.475 ;
      RECT 5.57 1.235 7.49 1.405 ;
      RECT 5.57 1.405 5.74 1.915 ;
      RECT 5.57 1.915 6.78 2.085 ;
      RECT 5.57 2.085 5.74 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.8 0.895 6.15 1.015 ;
      RECT 5.91 1.575 7.88 1.745 ;
      RECT 5.92 2.255 6.34 2.635 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 6.69 0.085 7.33 0.565 ;
      RECT 7.01 1.945 7.34 2.635 ;
      RECT 7.14 1.175 7.49 1.235 ;
      RECT 7.51 1.745 7.88 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.53 0.35 7.88 0.68 ;
      RECT 7.69 0.68 7.88 1.575 ;
      RECT 7.97 1.915 8.3 2.425 ;
      RECT 8.05 0.345 8.22 0.995 ;
      RECT 8.05 0.995 8.85 1.325 ;
      RECT 8.05 1.325 8.3 1.915 ;
      RECT 8.39 0.085 8.72 0.825 ;
      RECT 8.47 1.495 8.64 2.635 ;
      RECT 9.305 0.085 9.575 0.595 ;
      RECT 9.31 1.785 9.575 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 1.785 0.775 1.955 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.225 1.105 5.395 1.275 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.545 1.755 0.835 1.8 ;
      RECT 0.545 1.8 5.435 1.94 ;
      RECT 0.545 1.94 0.835 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.455 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.165 1.075 5.455 1.12 ;
      RECT 5.165 1.26 5.455 1.305 ;
  END
END sky130_fd_sc_hd__dfstp_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 6.125 4.595 6.295 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 6.3 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 6.01 3.455 6.3 3.5 ;
        RECT 6.01 3.64 6.3 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 6.63 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.37 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 6.44 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 6.44 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.825 0.085 6.155 0.9 ;
      RECT 5.905 1.61 6.075 2.635 ;
      RECT 6.065 2.985 6.355 3.955 ;
      RECT 6.065 4.63 6.355 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 6.07 3.485 6.24 3.655 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 6.44 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 7.045 4.595 7.215 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 7.29 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 6.93 3.455 7.22 3.5 ;
        RECT 6.93 3.64 7.22 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 7.405 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 7.36 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 7.36 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.825 0.085 6.155 0.845 ;
      RECT 5.905 1.61 6.075 2.635 ;
      RECT 6.755 0.085 7.005 0.925 ;
      RECT 6.755 1.61 6.935 2.635 ;
      RECT 6.985 2.985 7.275 3.955 ;
      RECT 6.985 4.63 7.275 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.585 5.355 6.755 5.525 ;
      RECT 6.99 3.485 7.16 3.655 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.045 5.355 7.215 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 7.36 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.29 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 5.925 4.595 6.095 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 6.17 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 5.87 3.455 6.16 3.5 ;
        RECT 5.87 3.64 6.16 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 6.63 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.17 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 6.44 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.29 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.29 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 6.44 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.865 0.085 6.155 0.81 ;
      RECT 5.865 2.985 6.155 3.955 ;
      RECT 5.865 4.63 6.155 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 5.93 3.485 6.1 3.655 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 6.44 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
      RECT 5.925 0.32 6.095 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.050000 0.315000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_2
MACRO sky130_fd_sc_hd__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130000 -0.120000 0.350000 0.050000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_8
MACRO sky130_fd_sc_hd__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.055000 0.260000 0.055000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_1
MACRO sky130_fd_sc_hd__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175000 -0.060000 0.285000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_4
MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.56 1.29 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705 0.27 3.15 0.64 ;
        RECT 2.715 1.42 3.18 1.525 ;
        RECT 2.715 1.525 3.15 2.465 ;
        RECT 2.965 0.64 3.15 0.78 ;
        RECT 2.965 0.78 3.18 0.945 ;
        RECT 3.01 0.945 3.18 1.42 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.27 0.415 0.735 ;
      RECT 0.085 0.735 1.055 0.905 ;
      RECT 0.085 1.46 1.055 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.585 0.085 0.915 0.565 ;
      RECT 0.6 1.8 0.93 2.635 ;
      RECT 0.73 0.905 1.055 1.46 ;
      RECT 1.11 1.8 1.44 2.465 ;
      RECT 1.16 0.27 1.44 0.6 ;
      RECT 1.27 0.6 1.44 1.075 ;
      RECT 1.27 1.075 2.205 1.255 ;
      RECT 1.27 1.255 1.44 1.8 ;
      RECT 1.63 0.27 1.96 0.735 ;
      RECT 1.63 0.735 2.545 0.905 ;
      RECT 1.63 1.46 2.545 1.63 ;
      RECT 1.63 1.63 1.96 2.465 ;
      RECT 2.13 1.8 2.545 2.635 ;
      RECT 2.165 0.085 2.535 0.565 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 2.84 1.245 ;
      RECT 2.375 1.245 2.545 1.46 ;
      RECT 3.32 0.085 3.595 0.645 ;
      RECT 3.32 1.625 3.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2
MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.055 0.55 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.255 3.59 0.545 ;
        RECT 3.22 1.76 3.59 2.465 ;
        RECT 3.365 0.545 3.59 1.76 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.095 0.255 0.425 0.715 ;
      RECT 0.095 0.715 1.215 0.885 ;
      RECT 0.095 1.495 1.215 1.665 ;
      RECT 0.095 1.665 0.425 2.465 ;
      RECT 0.595 0.085 0.91 0.545 ;
      RECT 0.595 1.835 0.925 2.635 ;
      RECT 0.72 0.885 1.215 1.495 ;
      RECT 1.385 0.255 1.76 0.825 ;
      RECT 1.385 1.835 1.76 2.465 ;
      RECT 1.59 0.825 1.76 1.055 ;
      RECT 1.59 1.055 2.685 1.25 ;
      RECT 1.59 1.25 1.76 1.835 ;
      RECT 1.93 0.255 2.26 0.715 ;
      RECT 1.93 0.715 3.195 0.885 ;
      RECT 1.93 1.42 3.195 1.59 ;
      RECT 1.93 1.59 2.26 2.465 ;
      RECT 2.71 0.085 3.04 0.545 ;
      RECT 2.71 1.76 3.04 2.635 ;
      RECT 2.855 0.885 3.195 1.42 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1
MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.075 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.43 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.865 2.465 ;
        RECT 0.6 0.255 1.295 0.885 ;
        RECT 0.6 0.885 0.77 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.085 0.085 0.395 0.885 ;
      RECT 0.085 1.495 0.365 2.635 ;
      RECT 1.035 1.495 1.295 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__nand2_1
MACRO sky130_fd_sc_hd__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.29 1.075 6.305 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.51 1.075 3.365 1.295 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.465 6.725 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 3.64 1.075 4.12 1.465 ;
        RECT 3.875 0.655 6.725 0.905 ;
        RECT 3.875 0.905 4.12 1.075 ;
        RECT 3.875 1.665 4.205 2.465 ;
        RECT 4.715 1.665 5.045 2.465 ;
        RECT 5.555 1.665 5.885 2.465 ;
        RECT 6.395 1.665 6.725 2.465 ;
        RECT 6.475 0.905 6.725 1.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 3.705 0.905 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.595 0.085 0.765 0.565 ;
      RECT 0.935 0.255 1.265 0.735 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.435 0.085 1.605 0.565 ;
      RECT 1.775 0.255 2.105 0.735 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.275 0.085 2.445 0.565 ;
      RECT 2.615 0.255 2.945 0.735 ;
      RECT 2.695 1.835 2.865 2.635 ;
      RECT 3.115 0.085 3.285 0.565 ;
      RECT 3.455 0.255 7.27 0.485 ;
      RECT 3.455 0.485 3.705 0.735 ;
      RECT 3.535 1.835 3.705 2.635 ;
      RECT 4.375 1.835 4.545 2.635 ;
      RECT 5.215 1.835 5.385 2.635 ;
      RECT 6.055 1.835 6.225 2.635 ;
      RECT 6.895 0.485 7.27 0.905 ;
      RECT 6.915 1.495 7.27 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__nand2_8
MACRO sky130_fd_sc_hd__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.055 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.73 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 3.365 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 1.91 1.075 2.445 1.495 ;
        RECT 2.195 0.635 3.365 0.805 ;
        RECT 2.195 0.805 2.445 1.075 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.255 0.425 0.715 ;
      RECT 0.09 0.715 2.025 0.905 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.935 0.255 1.265 0.715 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.435 0.085 1.605 0.545 ;
      RECT 1.775 0.255 3.785 0.465 ;
      RECT 1.775 0.465 2.025 0.715 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.695 1.835 2.865 2.635 ;
      RECT 3.535 0.465 3.785 0.885 ;
      RECT 3.535 1.835 3.785 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__nand2_4
MACRO sky130_fd_sc_hd__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.765 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.845 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 2.215 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 0.655 2.215 0.905 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 1.935 0.905 2.215 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.185 0.885 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 0.595 0.085 0.765 0.545 ;
      RECT 0.935 0.255 2.105 0.465 ;
      RECT 0.935 0.465 1.185 0.715 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.775 0.465 2.105 0.485 ;
      RECT 1.855 1.835 2.11 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nand2_2
MACRO sky130_fd_sc_hd__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2 0.995 3.115 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.805 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.995 0.8 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 0.995 4.055 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.73 1.075 5.41 1.295 ;
        RECT 5.175 1.295 5.41 1.625 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295 0.655 5.345 0.825 ;
        RECT 3.235 0.255 3.405 0.655 ;
        RECT 4.085 0.255 4.255 0.655 ;
        RECT 4.26 0.825 4.475 1.51 ;
        RECT 4.26 1.51 4.99 1.575 ;
        RECT 4.26 1.575 5.005 1.68 ;
        RECT 4.66 1.68 5.005 1.745 ;
        RECT 4.66 1.745 4.99 1.915 ;
        RECT 4.66 1.915 5.005 2.085 ;
        RECT 5.175 0.255 5.345 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.095 1.495 0.345 2.635 ;
      RECT 0.175 0.255 0.345 0.655 ;
      RECT 0.175 0.655 2.105 0.825 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.595 1.575 3.915 1.745 ;
      RECT 0.595 1.745 0.765 2.465 ;
      RECT 0.935 1.915 1.265 2.635 ;
      RECT 1.015 0.255 1.185 0.655 ;
      RECT 1.355 0.305 3.045 0.475 ;
      RECT 1.435 1.745 1.605 2.465 ;
      RECT 1.785 1.915 2.135 2.635 ;
      RECT 2.305 1.745 2.475 2.465 ;
      RECT 2.645 1.915 2.975 2.635 ;
      RECT 3.145 2.255 5.345 2.425 ;
      RECT 3.585 0.085 3.915 0.465 ;
      RECT 3.585 1.745 3.915 2.085 ;
      RECT 4.11 1.915 4.44 2.255 ;
      RECT 4.11 2.425 4.44 2.465 ;
      RECT 4.675 0.085 5.005 0.465 ;
      RECT 5.175 1.795 5.345 2.255 ;
      RECT 5.175 2.425 5.345 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__a311oi_2
MACRO sky130_fd_sc_hd__a311oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.265 1.365 0.66 ;
        RECT 1.195 0.66 1.365 0.995 ;
        RECT 1.195 0.995 1.455 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.6 0.265 0.795 0.995 ;
        RECT 0.6 0.995 1.025 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.42 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.71 0.995 1.935 1.835 ;
        RECT 1.71 1.835 2.23 2.005 ;
        RECT 1.95 2.005 2.23 2.355 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.685 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.659750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 0.255 1.705 0.655 ;
        RECT 1.535 0.655 2.65 0.825 ;
        RECT 2.105 0.825 2.275 1.495 ;
        RECT 2.105 1.495 2.65 1.665 ;
        RECT 2.405 0.295 2.65 0.655 ;
        RECT 2.41 1.665 2.65 2.335 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.085 0.325 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.095 0.085 0.425 0.805 ;
      RECT 0.095 1.495 0.425 2.635 ;
      RECT 0.6 1.575 1.54 1.745 ;
      RECT 0.6 1.745 0.77 2.305 ;
      RECT 0.94 1.915 1.2 2.635 ;
      RECT 1.37 1.745 1.54 2.175 ;
      RECT 1.37 2.175 1.7 2.345 ;
      RECT 1.905 0.085 2.235 0.485 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a311oi_1
MACRO sky130_fd_sc_hd__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.995 5.42 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.55 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.67 0.995 6.855 1.63 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.935 0.995 9.53 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.898500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.635 9.485 0.805 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.415 0.255 7.585 0.635 ;
        RECT 7.415 0.805 7.735 1.545 ;
        RECT 7.415 1.545 9.145 1.715 ;
        RECT 7.415 1.715 7.735 1.975 ;
        RECT 7.975 1.53 8.305 1.545 ;
        RECT 7.975 1.715 8.305 2.085 ;
        RECT 8.475 0.255 8.645 0.635 ;
        RECT 8.815 1.715 9.145 2.085 ;
        RECT 9.315 0.255 9.485 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.095 1.575 0.425 2.635 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 3.785 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.595 1.495 4.965 1.665 ;
      RECT 0.595 1.665 0.765 2.465 ;
      RECT 0.935 1.915 1.265 2.635 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.355 0.085 1.685 0.465 ;
      RECT 1.435 1.665 1.605 2.465 ;
      RECT 1.775 1.915 2.105 2.635 ;
      RECT 1.855 0.255 2.025 0.635 ;
      RECT 2.195 0.295 5.565 0.465 ;
      RECT 2.275 1.665 2.445 2.465 ;
      RECT 2.615 1.915 2.945 2.635 ;
      RECT 3.115 1.665 3.285 2.465 ;
      RECT 3.455 1.915 3.785 2.635 ;
      RECT 3.955 1.665 4.125 2.465 ;
      RECT 4.295 1.915 4.625 2.635 ;
      RECT 4.795 1.665 4.965 1.915 ;
      RECT 4.795 1.915 7.245 2.085 ;
      RECT 4.795 2.085 4.965 2.465 ;
      RECT 5.135 2.255 5.465 2.635 ;
      RECT 5.655 2.255 9.565 2.425 ;
      RECT 6.075 0.085 6.405 0.465 ;
      RECT 6.915 0.085 7.245 0.465 ;
      RECT 7.975 0.085 8.305 0.465 ;
      RECT 8.815 0.085 9.145 0.465 ;
      RECT 9.315 1.835 9.565 2.255 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__a311oi_4
MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.555 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.41 0.255 2.7 0.825 ;
        RECT 2.44 1.495 2.7 2.465 ;
        RECT 2.53 0.825 2.7 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.785 0.895 2.005 ;
      RECT 0.085 2.005 0.38 2.465 ;
      RECT 0.095 0.255 0.38 0.715 ;
      RECT 0.095 0.715 0.895 0.885 ;
      RECT 0.55 0.085 0.765 0.545 ;
      RECT 0.55 2.175 0.765 2.635 ;
      RECT 0.725 0.885 0.895 0.995 ;
      RECT 0.725 0.995 0.98 1.325 ;
      RECT 0.725 1.325 0.895 1.785 ;
      RECT 0.935 0.255 1.32 0.545 ;
      RECT 0.935 2.175 1.32 2.465 ;
      RECT 1.15 0.545 1.32 1.075 ;
      RECT 1.15 1.075 1.9 1.275 ;
      RECT 1.15 1.275 1.32 2.175 ;
      RECT 1.515 0.255 1.74 0.735 ;
      RECT 1.515 0.735 2.24 0.905 ;
      RECT 1.515 1.575 2.24 1.745 ;
      RECT 1.515 1.745 1.74 2.43 ;
      RECT 1.91 0.085 2.24 0.565 ;
      RECT 1.91 1.915 2.27 2.635 ;
      RECT 2.07 0.905 2.24 0.995 ;
      RECT 2.07 0.995 2.36 1.325 ;
      RECT 2.07 1.325 2.24 1.575 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1
MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 0.635 1.02 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 2.125 1.345 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.145 0.305 1.365 0.79 ;
        RECT 1.145 0.79 1.475 1.215 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.765 2.215 2.465 ;
        RECT 1.955 0.255 2.215 0.735 ;
        RECT 2.045 0.735 2.215 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.295 0.975 0.465 ;
      RECT 0.085 1.19 0.975 1.26 ;
      RECT 0.085 1.26 0.98 1.285 ;
      RECT 0.085 1.285 0.99 1.3 ;
      RECT 0.085 1.3 0.995 1.315 ;
      RECT 0.085 1.315 1.005 1.32 ;
      RECT 0.085 1.32 1.01 1.33 ;
      RECT 0.085 1.33 1.015 1.34 ;
      RECT 0.085 1.34 1.025 1.345 ;
      RECT 0.085 1.345 1.035 1.355 ;
      RECT 0.085 1.355 1.045 1.36 ;
      RECT 0.085 1.36 0.345 1.81 ;
      RECT 0.085 1.98 0.7 2.08 ;
      RECT 0.085 2.08 0.69 2.635 ;
      RECT 0.515 1.71 0.845 1.955 ;
      RECT 0.515 1.955 0.7 1.98 ;
      RECT 0.71 1.36 1.045 1.365 ;
      RECT 0.71 1.365 1.06 1.37 ;
      RECT 0.71 1.37 1.075 1.38 ;
      RECT 0.71 1.38 1.1 1.385 ;
      RECT 0.71 1.385 1.875 1.39 ;
      RECT 0.74 1.39 1.875 1.425 ;
      RECT 0.775 1.425 1.875 1.45 ;
      RECT 0.805 0.465 0.975 1.19 ;
      RECT 0.805 1.45 1.875 1.48 ;
      RECT 0.825 1.48 1.875 1.51 ;
      RECT 0.845 1.51 1.875 1.54 ;
      RECT 0.915 1.54 1.875 1.55 ;
      RECT 0.94 1.55 1.875 1.56 ;
      RECT 0.96 1.56 1.875 1.575 ;
      RECT 0.98 1.575 1.875 1.59 ;
      RECT 0.985 1.59 1.77 1.6 ;
      RECT 1 1.6 1.77 1.635 ;
      RECT 1.015 1.635 1.77 1.885 ;
      RECT 1.515 2.09 1.77 2.635 ;
      RECT 1.535 0.085 1.785 0.625 ;
      RECT 1.645 0.99 1.875 1.385 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__and3_1
MACRO sky130_fd_sc_hd__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.995 0.875 1.34 ;
        RECT 0.115 1.34 0.365 2.335 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.745 1.355 1.34 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.9 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.515 2.64 0.615 ;
        RECT 2.45 0.615 4.055 0.845 ;
        RECT 2.45 1.535 4.055 1.76 ;
        RECT 2.45 1.76 2.64 2.465 ;
        RECT 3.31 0.255 3.5 0.615 ;
        RECT 3.31 1.76 4.055 1.765 ;
        RECT 3.31 1.765 3.5 2.465 ;
        RECT 3.775 0.845 4.055 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.465 0.255 0.8 0.375 ;
      RECT 0.465 0.375 1.725 0.565 ;
      RECT 0.465 0.565 0.8 0.805 ;
      RECT 0.545 1.58 2.28 1.75 ;
      RECT 0.545 1.75 0.725 2.465 ;
      RECT 0.895 1.935 1.345 2.635 ;
      RECT 1.52 1.75 1.7 2.465 ;
      RECT 1.535 0.565 1.725 0.615 ;
      RECT 1.535 0.615 2.28 0.805 ;
      RECT 1.905 0.085 2.235 0.445 ;
      RECT 1.91 1.935 2.24 2.635 ;
      RECT 2.07 0.805 2.28 1.02 ;
      RECT 2.07 1.02 3.605 1.355 ;
      RECT 2.07 1.355 2.28 1.58 ;
      RECT 2.81 0.085 3.14 0.445 ;
      RECT 2.81 1.935 3.14 2.635 ;
      RECT 3.67 0.085 4 0.445 ;
      RECT 3.67 1.935 4 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__and3_4
MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.47 1.245 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895 2.125 1.37 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.305 1.295 0.75 ;
        RECT 1.065 0.75 1.475 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 1.795 2.245 2.465 ;
        RECT 1.98 0.255 2.23 0.715 ;
        RECT 2.06 0.715 2.23 0.925 ;
        RECT 2.06 0.925 2.675 1.445 ;
        RECT 2.075 1.445 2.245 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 2.13 0.715 2.635 ;
      RECT 0.1 1.425 1.89 1.595 ;
      RECT 0.1 1.595 0.355 1.96 ;
      RECT 0.105 0.305 0.895 0.57 ;
      RECT 0.525 1.765 0.855 1.955 ;
      RECT 0.525 1.955 0.715 2.13 ;
      RECT 0.64 0.57 0.895 1.425 ;
      RECT 1.08 1.595 1.33 1.89 ;
      RECT 1.475 0.085 1.805 0.58 ;
      RECT 1.555 1.79 1.77 2.635 ;
      RECT 1.66 0.995 1.89 1.425 ;
      RECT 2.4 0.085 2.675 0.745 ;
      RECT 2.415 1.625 2.675 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__and3_2
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 2.675 2.465 ;
        RECT 1.465 1.025 2.675 1.545 ;
      LAYER mcon ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 2.69 2.34 ;
        RECT 0.085 2.08 2.675 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.085 2.675 0.855 ;
      RECT 0.085 0.855 1.295 1.375 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_6
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 1.755 2.465 ;
        RECT 1.005 1.025 1.755 1.545 ;
      LAYER mcon ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.085 2.08 1.755 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.085 0.085 1.755 0.855 ;
      RECT 0.085 0.855 0.835 1.375 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_4
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 5.43 2.465 ;
        RECT 2.835 1.025 5.43 1.545 ;
      LAYER mcon ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 2.905 2.125 3.075 2.295 ;
        RECT 3.365 2.125 3.535 2.295 ;
        RECT 3.825 2.125 3.995 2.295 ;
        RECT 4.285 2.125 4.455 2.295 ;
        RECT 4.745 2.125 4.915 2.295 ;
        RECT 5.205 2.125 5.375 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 5.45 2.34 ;
        RECT 0.085 2.08 5.435 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.085 0.085 5.43 0.855 ;
      RECT 0.085 0.855 2.665 1.375 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_12
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 3.595 2.465 ;
        RECT 1.905 1.025 3.595 1.545 ;
      LAYER mcon ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 2.905 2.125 3.075 2.295 ;
        RECT 3.365 2.125 3.535 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 3.61 2.34 ;
        RECT 0.085 2.08 3.595 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.085 3.595 0.855 ;
      RECT 0.085 0.855 1.735 1.375 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_8
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 1.295 2.465 ;
        RECT 0.775 1.005 1.295 1.545 ;
      LAYER mcon ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.085 2.08 1.295 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.085 0.085 1.295 0.835 ;
      RECT 0.085 0.835 0.605 1.375 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_3
MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.74 1.02 4.975 1.275 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.637500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.635 4.975 0.85 ;
        RECT 3.19 0.85 3.57 1.445 ;
        RECT 3.19 1.445 4.36 1.615 ;
        RECT 3.19 1.615 3.52 2.125 ;
        RECT 4.03 1.615 4.36 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.695 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.695 0.995 ;
      RECT 0.5 0.995 3.02 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 2.125 0.875 2.635 ;
      RECT 1.035 0.255 1.205 0.655 ;
      RECT 1.035 0.655 3.02 0.825 ;
      RECT 1.075 1.555 2.995 1.725 ;
      RECT 1.075 1.725 1.285 2.465 ;
      RECT 1.375 0.085 1.705 0.485 ;
      RECT 1.455 1.895 1.785 2.635 ;
      RECT 1.875 0.255 2.045 0.655 ;
      RECT 1.955 1.725 2.125 2.465 ;
      RECT 2.215 0.085 2.555 0.485 ;
      RECT 2.295 1.895 2.655 2.635 ;
      RECT 2.735 0.255 4.975 0.465 ;
      RECT 2.735 0.465 3.02 0.655 ;
      RECT 2.825 1.725 2.995 2.295 ;
      RECT 2.825 2.295 4.975 2.465 ;
      RECT 3.69 1.785 3.86 2.295 ;
      RECT 4.53 1.445 4.975 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__einvp_4
MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.42 1.02 8.195 1.275 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.027500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.87 0.635 8.195 0.85 ;
        RECT 4.87 0.85 5.25 1.445 ;
        RECT 4.87 1.445 7.72 1.615 ;
        RECT 4.87 1.615 5.2 2.125 ;
        RECT 5.71 1.615 6.04 2.125 ;
        RECT 6.55 1.615 6.88 2.125 ;
        RECT 7.39 1.615 7.72 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.695 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.695 0.995 ;
      RECT 0.5 0.995 4.7 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 2.125 0.875 2.635 ;
      RECT 1.035 0.255 1.205 0.655 ;
      RECT 1.035 0.655 4.7 0.825 ;
      RECT 1.075 1.555 4.7 1.725 ;
      RECT 1.075 1.725 1.285 2.465 ;
      RECT 1.375 0.085 1.705 0.485 ;
      RECT 1.455 1.895 1.785 2.635 ;
      RECT 1.875 0.255 2.045 0.655 ;
      RECT 1.955 1.725 2.125 2.465 ;
      RECT 2.215 0.085 2.545 0.485 ;
      RECT 2.295 1.895 2.625 2.635 ;
      RECT 2.715 0.255 2.885 0.655 ;
      RECT 2.795 1.725 2.965 2.465 ;
      RECT 3.055 0.085 3.385 0.485 ;
      RECT 3.135 1.895 3.465 2.635 ;
      RECT 3.555 0.255 3.725 0.655 ;
      RECT 3.635 1.725 3.805 2.465 ;
      RECT 3.895 0.085 4.235 0.485 ;
      RECT 3.975 1.895 4.305 2.635 ;
      RECT 4.405 0.255 8.195 0.465 ;
      RECT 4.405 0.465 4.7 0.655 ;
      RECT 4.475 1.725 4.7 2.295 ;
      RECT 4.475 2.295 8.195 2.465 ;
      RECT 5.37 1.785 5.54 2.295 ;
      RECT 6.21 1.785 6.38 2.295 ;
      RECT 7.05 1.785 7.22 2.295 ;
      RECT 7.89 1.445 8.195 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
  END
END sky130_fd_sc_hd__einvp_8
MACRO sky130_fd_sc_hd__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.975 2.215 1.955 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.223500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.545 1.725 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.62 0.255 2.215 0.805 ;
        RECT 1.62 0.805 1.795 2.125 ;
        RECT 1.62 2.125 2.215 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 1.45 0.825 ;
      RECT 0.085 1.895 1.45 2.065 ;
      RECT 0.085 2.065 0.345 2.465 ;
      RECT 0.515 0.085 1.45 0.485 ;
      RECT 0.515 2.235 1.45 2.635 ;
      RECT 0.715 0.825 1.45 1.895 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__einvp_1
MACRO sky130_fd_sc_hd__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.85 0.765 3.135 1.615 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.354000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 0.595 2.68 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.875 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.875 0.995 ;
      RECT 0.5 0.995 2.18 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 0.515 0.085 0.875 0.485 ;
      RECT 0.515 2.125 0.875 2.635 ;
      RECT 1.045 0.255 1.24 0.655 ;
      RECT 1.045 0.655 2.18 0.825 ;
      RECT 1.045 1.555 2.155 1.725 ;
      RECT 1.045 1.725 1.285 2.465 ;
      RECT 1.41 0.085 1.77 0.485 ;
      RECT 1.455 1.895 1.785 2.635 ;
      RECT 1.94 0.255 3.135 0.425 ;
      RECT 1.94 0.425 2.18 0.655 ;
      RECT 1.985 1.725 2.155 2.295 ;
      RECT 1.985 2.295 3.135 2.465 ;
      RECT 2.85 0.425 3.135 0.595 ;
      RECT 2.85 1.785 3.135 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__einvp_2
MACRO sky130_fd_sc_hd__clkinvlp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.6 1.665 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.436750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.81 0.315 1.445 0.75 ;
        RECT 0.81 0.75 1.235 2.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.225 1.835 0.555 2.625 ;
      RECT 0.225 2.625 1.74 2.635 ;
      RECT 0.295 0.085 0.625 0.745 ;
      RECT 1.44 1.455 1.74 2.625 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__clkinvlp_2
MACRO sky130_fd_sc_hd__clkinvlp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.425 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.714000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.255 1.215 0.68 ;
        RECT 0.595 0.68 0.955 1.015 ;
        RECT 0.595 1.015 2.015 1.295 ;
        RECT 0.595 1.295 0.955 2.465 ;
        RECT 1.685 1.295 2.015 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 0.085 0.425 0.575 ;
      RECT 0.095 1.495 0.425 2.635 ;
      RECT 1.155 1.465 1.485 2.635 ;
      RECT 1.675 0.085 2.005 0.775 ;
      RECT 2.215 1.465 2.545 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__clkinvlp_4
MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 1.415 1.275 ;
        RECT 1.15 1.275 1.415 1.445 ;
        RECT 1.15 1.445 3.575 1.615 ;
        RECT 3.275 1.075 3.605 1.245 ;
        RECT 3.275 1.245 3.575 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.685 1.075 3.095 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 0.995 4.94 1.445 ;
        RECT 4.295 1.445 6.935 1.615 ;
        RECT 6.715 0.995 6.935 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.11 1.075 6.46 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.785 3.915 1.955 ;
        RECT 1.845 1.955 2.095 2.125 ;
        RECT 2.685 1.955 2.935 2.125 ;
        RECT 3.745 1.445 4.125 1.615 ;
        RECT 3.745 1.615 3.915 1.785 ;
        RECT 3.955 0.645 7.275 0.82 ;
        RECT 3.955 0.82 4.125 1.445 ;
        RECT 5.255 1.785 7.275 1.955 ;
        RECT 5.255 1.955 5.505 2.125 ;
        RECT 6.095 1.955 6.345 2.125 ;
        RECT 7.105 0.82 7.275 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.125 0.255 0.455 0.725 ;
      RECT 0.125 0.725 1.295 0.735 ;
      RECT 0.125 0.735 3.785 0.905 ;
      RECT 0.165 1.445 0.415 2.635 ;
      RECT 0.585 1.445 0.835 1.785 ;
      RECT 0.585 1.785 1.675 1.955 ;
      RECT 0.585 1.955 0.835 2.465 ;
      RECT 0.625 0.085 0.795 0.555 ;
      RECT 0.965 0.255 1.295 0.725 ;
      RECT 1.005 2.125 1.255 2.635 ;
      RECT 1.425 1.955 1.675 2.295 ;
      RECT 1.425 2.295 3.395 2.465 ;
      RECT 1.465 0.085 1.635 0.555 ;
      RECT 1.805 0.255 2.135 0.725 ;
      RECT 1.805 0.725 2.975 0.735 ;
      RECT 2.265 2.125 2.515 2.295 ;
      RECT 2.305 0.085 2.475 0.555 ;
      RECT 2.645 0.255 2.975 0.725 ;
      RECT 3.105 2.125 3.395 2.295 ;
      RECT 3.145 0.085 3.315 0.555 ;
      RECT 3.485 0.255 7.245 0.475 ;
      RECT 3.485 0.475 3.785 0.735 ;
      RECT 3.565 2.125 3.785 2.635 ;
      RECT 3.955 2.125 4.255 2.465 ;
      RECT 4.085 1.785 5.085 1.955 ;
      RECT 4.085 1.955 4.255 2.125 ;
      RECT 4.425 2.125 4.665 2.635 ;
      RECT 4.835 1.955 5.085 2.295 ;
      RECT 4.835 2.295 6.765 2.465 ;
      RECT 5.675 2.125 5.925 2.295 ;
      RECT 6.515 2.135 6.765 2.295 ;
      RECT 6.935 2.125 7.215 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__o22ai_4
MACRO sky130_fd_sc_hd__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.215 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.22 1.075 1.585 1.245 ;
        RECT 1.405 1.245 1.585 1.445 ;
        RECT 1.405 1.445 1.725 1.615 ;
        RECT 1.525 1.615 1.725 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.665 0.325 1.99 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 0.995 1.005 1.415 ;
        RECT 0.835 1.415 1.235 1.665 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.650250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495 0.645 0.845 0.825 ;
        RECT 0.495 0.825 0.665 1.835 ;
        RECT 0.495 1.835 1.335 2.045 ;
        RECT 0.835 2.045 1.335 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.295 1.345 0.475 ;
      RECT 0.135 2.175 0.345 2.635 ;
      RECT 1.015 0.475 1.345 0.695 ;
      RECT 1.015 0.695 2.215 0.825 ;
      RECT 1.185 0.825 2.215 0.865 ;
      RECT 1.535 0.085 1.705 0.525 ;
      RECT 1.875 0.28 2.215 0.695 ;
      RECT 1.895 1.455 2.215 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__o22ai_1
MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.165 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.075 3.225 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.2 1.075 0.985 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.075 1.925 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.645 0.865 0.725 ;
        RECT 0.535 0.725 2.34 0.905 ;
        RECT 1.375 0.645 1.705 0.725 ;
        RECT 1.415 1.445 3.065 1.625 ;
        RECT 1.415 1.625 1.665 2.125 ;
        RECT 2.095 0.905 2.34 1.445 ;
        RECT 2.815 1.625 3.065 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.09 0.305 2.68 0.475 ;
      RECT 0.09 0.475 0.365 0.905 ;
      RECT 0.15 1.455 1.245 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.295 ;
      RECT 0.995 2.295 2.085 2.465 ;
      RECT 1.835 1.795 2.085 2.295 ;
      RECT 2.395 1.795 2.645 2.295 ;
      RECT 2.395 2.295 3.485 2.465 ;
      RECT 2.51 0.475 2.68 0.725 ;
      RECT 2.51 0.725 4.365 0.905 ;
      RECT 2.855 0.085 3.025 0.555 ;
      RECT 3.195 0.255 3.525 0.725 ;
      RECT 3.235 1.455 4.33 1.625 ;
      RECT 3.235 1.625 3.485 2.295 ;
      RECT 3.655 1.795 3.905 2.635 ;
      RECT 3.695 0.085 3.865 0.555 ;
      RECT 4.035 0.255 4.365 0.725 ;
      RECT 4.075 1.625 4.33 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__o22ai_2
MACRO sky130_fd_sc_hd__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 0.995 2.175 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.37 0.995 2.63 1.615 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.325 0.335 1.665 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.3 0.265 3.58 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.105 1.845 0.855 2.045 ;
      RECT 0.105 2.045 0.345 2.435 ;
      RECT 0.515 0.265 0.745 1.165 ;
      RECT 0.515 1.165 0.855 1.845 ;
      RECT 0.515 2.225 0.865 2.635 ;
      RECT 0.945 0.085 1.19 0.865 ;
      RECT 1.035 1.045 1.58 1.345 ;
      RECT 1.035 1.345 1.365 2.455 ;
      RECT 1.36 0.265 1.79 0.625 ;
      RECT 1.36 0.625 3.1 0.815 ;
      RECT 1.36 0.815 1.58 1.045 ;
      RECT 1.535 1.785 2.56 1.985 ;
      RECT 1.535 1.985 1.715 2.455 ;
      RECT 1.885 2.155 2.215 2.635 ;
      RECT 2.37 0.085 3.1 0.455 ;
      RECT 2.39 1.985 2.56 2.455 ;
      RECT 2.825 1.495 3.11 2.635 ;
      RECT 2.84 0.815 3.1 1.325 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a21bo_1
MACRO sky130_fd_sc_hd__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.995 3.1 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.27 0.995 3.56 1.615 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.035 1.525 1.325 ;
        RECT 1.33 0.995 1.525 1.035 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.715 0.85 0.885 ;
        RECT 0.15 0.885 0.38 1.835 ;
        RECT 0.15 1.835 0.85 2.005 ;
        RECT 0.52 0.315 0.85 0.715 ;
        RECT 0.595 2.005 0.85 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 0.085 0.345 0.545 ;
      RECT 0.09 2.255 0.425 2.635 ;
      RECT 0.57 1.075 0.9 1.495 ;
      RECT 0.57 1.495 1.285 1.665 ;
      RECT 1.02 0.085 1.22 0.865 ;
      RECT 1.04 2.275 1.37 2.635 ;
      RECT 1.115 1.665 1.285 1.895 ;
      RECT 1.115 1.895 2.225 2.105 ;
      RECT 1.455 0.655 1.865 0.825 ;
      RECT 1.455 1.555 1.865 1.725 ;
      RECT 1.695 0.825 1.865 0.995 ;
      RECT 1.695 0.995 2.175 1.325 ;
      RECT 1.695 1.325 1.865 1.555 ;
      RECT 1.975 0.085 2.305 0.465 ;
      RECT 1.975 2.105 2.225 2.465 ;
      RECT 2.055 1.505 2.515 1.675 ;
      RECT 2.055 1.675 2.225 1.895 ;
      RECT 2.345 0.635 2.74 0.825 ;
      RECT 2.345 0.825 2.515 1.505 ;
      RECT 2.395 1.845 3.565 2.015 ;
      RECT 2.395 2.015 2.725 2.465 ;
      RECT 2.895 2.185 3.065 2.635 ;
      RECT 3.235 0.085 3.565 0.825 ;
      RECT 3.235 2.015 3.565 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a21bo_2
MACRO sky130_fd_sc_hd__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.59 1.01 4.955 1.36 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025 1.01 4.42 1.275 ;
        RECT 4.245 1.275 4.42 1.595 ;
        RECT 4.245 1.595 5.39 1.765 ;
        RECT 5.22 1.055 5.7 1.29 ;
        RECT 5.22 1.29 5.39 1.595 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.5 1.01 0.83 1.625 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 0.615 2.34 0.785 ;
        RECT 1 0.785 1.235 1.595 ;
        RECT 1 1.595 2.41 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.105 0.255 0.54 0.84 ;
      RECT 0.105 0.84 0.33 1.795 ;
      RECT 0.105 1.795 0.565 1.935 ;
      RECT 0.105 1.935 2.87 2.105 ;
      RECT 0.105 2.105 0.55 2.465 ;
      RECT 0.71 0.085 1.05 0.445 ;
      RECT 0.72 2.275 1.05 2.635 ;
      RECT 1.405 0.995 2.81 1.185 ;
      RECT 1.405 1.185 2.53 1.325 ;
      RECT 1.58 0.085 1.91 0.445 ;
      RECT 1.58 2.275 1.91 2.635 ;
      RECT 2.435 2.275 2.77 2.635 ;
      RECT 2.515 0.085 3.285 0.445 ;
      RECT 2.64 0.615 3.645 0.67 ;
      RECT 2.64 0.67 4.965 0.785 ;
      RECT 2.64 0.785 3.01 0.8 ;
      RECT 2.64 0.8 2.81 0.995 ;
      RECT 2.7 1.355 3.305 1.525 ;
      RECT 2.7 1.525 2.87 1.935 ;
      RECT 2.995 0.995 3.305 1.355 ;
      RECT 3.055 1.695 3.225 2.21 ;
      RECT 3.055 2.21 4.065 2.38 ;
      RECT 3.475 0.255 3.645 0.615 ;
      RECT 3.475 0.785 4.965 0.84 ;
      RECT 3.475 0.84 3.645 1.805 ;
      RECT 3.855 0.085 4.185 0.445 ;
      RECT 3.885 1.445 4.065 1.935 ;
      RECT 3.885 1.935 5.825 2.105 ;
      RECT 3.885 2.105 4.065 2.21 ;
      RECT 4.235 2.275 4.565 2.635 ;
      RECT 4.685 0.405 4.965 0.67 ;
      RECT 5.075 2.275 5.405 2.635 ;
      RECT 5.545 0.085 5.825 0.885 ;
      RECT 5.57 1.46 5.825 1.935 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__a21bo_4
MACRO sky130_fd_sc_hd__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 12.15 2.91 ;
        RECT 4.405 1.305 12.15 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.72 0.085 10.89 0.545 ;
      RECT 10.72 1.495 10.97 2.635 ;
      RECT 11.57 0.085 11.74 0.545 ;
      RECT 11.57 1.495 11.82 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_2
MACRO sky130_fd_sc_hd__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 0.995 ;
        RECT 11.19 0.995 12.24 1.325 ;
        RECT 11.19 1.325 11.4 1.445 ;
        RECT 11.99 0.265 12.24 0.995 ;
        RECT 11.99 1.325 12.24 2.325 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 13.07 2.91 ;
        RECT 4.405 1.305 13.07 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 12.88 0.085 ;
      RECT 0 2.635 12.88 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.72 0.085 10.89 0.545 ;
      RECT 10.72 1.495 10.97 2.635 ;
      RECT 11.57 0.085 11.74 0.545 ;
      RECT 11.57 1.495 11.82 2.635 ;
      RECT 12.41 0.085 12.58 0.545 ;
      RECT 12.41 1.495 12.66 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_4
MACRO sky130_fd_sc_hd__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.18 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.5 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 11.69 2.91 ;
        RECT 4.405 1.305 11.69 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.5 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.5 0.085 ;
      RECT 0 2.635 11.5 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.72 0.085 10.89 0.545 ;
      RECT 10.72 1.495 10.97 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_1
MACRO sky130_fd_sc_hd__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.82 1.075 9.575 1.34 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.11 1.075 7.325 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 5.455 1.345 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.075 3.55 1.345 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.755 1.345 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.984350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.645 1.685 0.815 ;
        RECT 0.085 0.815 0.375 1.515 ;
        RECT 0.085 1.515 7.39 1.685 ;
        RECT 0.085 1.685 0.36 2.465 ;
        RECT 1.015 1.685 1.195 2.465 ;
        RECT 1.845 1.685 2.035 2.465 ;
        RECT 2.685 1.685 2.875 2.465 ;
        RECT 3.525 1.685 3.715 2.465 ;
        RECT 4.57 1.685 4.76 2.465 ;
        RECT 5.41 1.685 5.6 2.465 ;
        RECT 6.285 1.685 6.48 2.1 ;
        RECT 7.045 1.685 7.39 1.72 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.095 0.285 2.025 0.475 ;
      RECT 0.53 1.855 0.845 2.635 ;
      RECT 1.39 1.855 1.675 2.635 ;
      RECT 1.855 0.475 2.025 0.615 ;
      RECT 1.855 0.615 3.785 0.825 ;
      RECT 2.195 0.255 5.565 0.445 ;
      RECT 2.205 1.855 2.515 2.635 ;
      RECT 3.045 1.855 3.355 2.635 ;
      RECT 3.975 0.655 9.44 0.905 ;
      RECT 4.075 1.855 4.4 2.635 ;
      RECT 4.93 1.855 5.22 2.635 ;
      RECT 5.785 1.855 6.115 2.27 ;
      RECT 5.785 2.27 7.005 2.465 ;
      RECT 6.1 0.085 6.43 0.485 ;
      RECT 6.705 1.89 8.235 2.06 ;
      RECT 6.705 2.06 7.005 2.27 ;
      RECT 6.96 0.085 7.29 0.485 ;
      RECT 7.555 2.23 7.885 2.635 ;
      RECT 7.825 0.085 8.155 0.485 ;
      RECT 8.045 1.515 9.08 1.685 ;
      RECT 8.045 1.685 8.235 1.89 ;
      RECT 8.055 2.06 8.235 2.465 ;
      RECT 8.41 1.855 8.72 2.635 ;
      RECT 8.665 0.085 8.995 0.485 ;
      RECT 8.89 1.685 9.08 2.465 ;
      RECT 9.265 1.535 9.575 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__o2111ai_4
MACRO sky130_fd_sc_hd__o2111ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.005 3.115 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.615 1.615 ;
        RECT 2.27 1.615 2.615 2.37 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.815 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.255 1.355 1.615 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485 1.075 0.815 1.615 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.857250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.69 0.885 ;
        RECT 0.085 0.885 0.315 1.785 ;
        RECT 0.085 1.785 2.095 2.025 ;
        RECT 0.79 2.025 1.025 2.465 ;
        RECT 1.75 2.025 2.095 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.29 2.195 0.62 2.635 ;
      RECT 1.21 2.255 1.54 2.635 ;
      RECT 1.75 0.255 2.095 0.625 ;
      RECT 1.75 0.625 3.115 0.825 ;
      RECT 2.285 0.085 2.615 0.455 ;
      RECT 2.785 0.255 3.115 0.625 ;
      RECT 2.785 1.795 3.115 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o2111ai_1
MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635 1.075 5.435 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.075 4.455 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.2 1.075 3.185 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.79 1.325 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.355 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.302000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.615 0.935 0.905 ;
        RECT 0.605 0.905 0.865 1.495 ;
        RECT 0.605 1.495 4.005 1.665 ;
        RECT 0.605 1.665 0.865 2.465 ;
        RECT 1.535 1.665 1.725 2.465 ;
        RECT 2.395 1.665 2.575 2.465 ;
        RECT 3.815 1.665 4.005 2.105 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.175 0.26 1.3 0.445 ;
      RECT 0.175 0.445 0.435 0.865 ;
      RECT 0.175 1.525 0.425 2.635 ;
      RECT 1.035 1.835 1.365 2.635 ;
      RECT 1.115 0.445 1.3 0.735 ;
      RECT 1.115 0.735 2.275 0.905 ;
      RECT 1.47 0.255 3.21 0.445 ;
      RECT 1.47 0.445 1.775 0.53 ;
      RECT 1.47 0.53 1.76 0.565 ;
      RECT 1.895 1.84 2.225 2.635 ;
      RECT 1.925 0.62 2.275 0.735 ;
      RECT 2.45 0.655 5.435 0.84 ;
      RECT 2.755 1.835 3.085 2.635 ;
      RECT 2.88 0.445 3.21 0.485 ;
      RECT 3.31 1.835 3.57 2.275 ;
      RECT 3.31 2.275 4.5 2.465 ;
      RECT 3.38 0.365 3.57 0.655 ;
      RECT 3.74 0.085 4.07 0.485 ;
      RECT 4.24 0.365 4.43 0.65 ;
      RECT 4.24 0.65 5.435 0.655 ;
      RECT 4.24 1.515 5.36 1.685 ;
      RECT 4.24 1.685 4.5 2.275 ;
      RECT 4.6 0.085 4.93 0.48 ;
      RECT 4.67 1.855 4.93 2.635 ;
      RECT 5.1 0.365 5.435 0.65 ;
      RECT 5.1 1.685 5.36 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__o2111ai_2
MACRO sky130_fd_sc_hd__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 5.525 1.315 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.58 0.255 0.91 0.715 ;
        RECT 0.58 0.715 6.79 0.905 ;
        RECT 0.58 1.495 6.79 1.665 ;
        RECT 0.58 1.665 0.91 2.465 ;
        RECT 1.42 0.255 1.75 0.715 ;
        RECT 1.42 1.665 1.75 2.465 ;
        RECT 2.26 0.255 2.59 0.715 ;
        RECT 2.26 1.665 2.59 2.465 ;
        RECT 3.1 0.255 3.43 0.715 ;
        RECT 3.1 1.665 3.43 2.465 ;
        RECT 3.94 0.255 4.27 0.715 ;
        RECT 3.94 1.665 4.27 2.465 ;
        RECT 4.78 0.255 5.11 0.715 ;
        RECT 4.78 1.665 5.11 2.465 ;
        RECT 5.62 0.255 5.95 0.715 ;
        RECT 5.62 1.665 5.95 2.465 ;
        RECT 6.46 0.255 6.79 0.715 ;
        RECT 6.46 0.905 6.79 1.495 ;
        RECT 6.46 1.665 6.79 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.18 0.085 0.41 0.885 ;
      RECT 0.2 1.485 0.41 2.635 ;
      RECT 1.08 0.085 1.25 0.545 ;
      RECT 1.08 1.835 1.25 2.635 ;
      RECT 1.92 0.085 2.09 0.545 ;
      RECT 1.92 1.835 2.09 2.635 ;
      RECT 2.76 0.085 2.93 0.545 ;
      RECT 2.76 1.835 2.93 2.635 ;
      RECT 3.6 0.085 3.77 0.545 ;
      RECT 3.6 1.835 3.77 2.635 ;
      RECT 4.44 0.085 4.61 0.545 ;
      RECT 4.44 1.835 4.61 2.635 ;
      RECT 5.28 0.085 5.45 0.545 ;
      RECT 5.28 1.835 5.45 2.635 ;
      RECT 6.12 0.085 6.29 0.545 ;
      RECT 6.12 1.835 6.29 2.635 ;
      RECT 6.96 0.085 7.17 0.885 ;
      RECT 6.96 1.835 7.17 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__inv_16
MACRO sky130_fd_sc_hd__inv_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 2.615 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.685 1.495 3.135 1.665 ;
        RECT 0.685 1.665 1.015 2.465 ;
        RECT 0.765 0.255 0.935 0.725 ;
        RECT 0.765 0.725 3.135 0.905 ;
        RECT 1.525 1.665 1.855 2.465 ;
        RECT 1.605 0.255 1.775 0.725 ;
        RECT 2.365 1.665 3.135 1.685 ;
        RECT 2.365 1.685 2.695 2.465 ;
        RECT 2.445 0.255 2.615 0.725 ;
        RECT 2.785 0.905 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.13 0.085 0.395 0.545 ;
      RECT 0.13 1.495 0.425 2.635 ;
      RECT 1.185 0.085 1.355 0.545 ;
      RECT 1.185 1.835 1.355 2.635 ;
      RECT 2.025 0.085 2.195 0.545 ;
      RECT 2.025 1.835 2.195 2.635 ;
      RECT 2.785 0.085 3.035 0.55 ;
      RECT 2.865 2.175 3.035 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__inv_6
MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.970000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.68 1.075 5.27 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 5.895 0.905 ;
        RECT 0.085 0.905 0.51 1.495 ;
        RECT 0.085 1.495 5.895 1.665 ;
        RECT 0.68 0.255 1.01 0.715 ;
        RECT 0.68 1.665 1.01 2.465 ;
        RECT 1.52 0.255 1.85 0.715 ;
        RECT 1.52 1.665 1.85 2.465 ;
        RECT 2.36 0.255 2.69 0.715 ;
        RECT 2.36 1.665 2.69 2.465 ;
        RECT 3.2 0.255 3.53 0.715 ;
        RECT 3.2 1.665 3.53 2.465 ;
        RECT 4.04 0.255 4.37 0.715 ;
        RECT 4.04 1.665 4.37 2.465 ;
        RECT 4.88 0.255 5.21 0.715 ;
        RECT 4.88 1.665 5.21 2.465 ;
        RECT 5.545 0.905 5.895 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.255 0.085 0.51 0.545 ;
      RECT 0.255 1.835 0.51 2.635 ;
      RECT 1.18 0.085 1.35 0.545 ;
      RECT 1.18 1.835 1.35 2.635 ;
      RECT 2.02 0.085 2.19 0.545 ;
      RECT 2.02 1.835 2.19 2.635 ;
      RECT 2.86 0.085 3.03 0.545 ;
      RECT 2.86 1.835 3.03 2.635 ;
      RECT 3.7 0.085 3.87 0.545 ;
      RECT 3.7 1.835 3.87 2.635 ;
      RECT 4.54 0.085 4.71 0.545 ;
      RECT 4.54 1.835 4.71 2.635 ;
      RECT 5.555 0.085 5.895 0.545 ;
      RECT 5.555 1.835 5.895 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__inv_12
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.32 1.075 0.65 1.315 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.72 0.255 1.05 0.885 ;
        RECT 0.72 1.485 1.05 2.465 ;
        RECT 0.82 0.885 1.05 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.32 0.085 0.55 0.905 ;
      RECT 0.34 1.495 0.55 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__inv_1
MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.255 0.855 0.885 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 0.605 0.885 0.855 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.125 0.085 0.355 0.905 ;
      RECT 0.125 1.495 0.355 2.635 ;
      RECT 1.025 0.085 1.235 0.905 ;
      RECT 1.025 1.495 1.235 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__inv_2
MACRO sky130_fd_sc_hd__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.68 1.075 3.535 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 4.055 0.905 ;
        RECT 0.085 0.905 0.43 1.495 ;
        RECT 0.085 1.495 4.055 1.665 ;
        RECT 0.68 0.255 1.01 0.715 ;
        RECT 0.68 1.665 1.01 2.465 ;
        RECT 1.52 0.255 1.85 0.715 ;
        RECT 1.52 1.665 1.85 2.465 ;
        RECT 2.36 0.255 2.69 0.715 ;
        RECT 2.36 1.665 2.69 2.465 ;
        RECT 3.2 0.255 3.53 0.715 ;
        RECT 3.2 1.665 3.53 2.465 ;
        RECT 3.735 0.905 4.055 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.255 0.085 0.51 0.545 ;
      RECT 0.255 1.835 0.51 2.635 ;
      RECT 1.18 0.085 1.35 0.545 ;
      RECT 1.18 1.835 1.35 2.635 ;
      RECT 2.02 0.085 2.19 0.545 ;
      RECT 2.02 1.835 2.19 2.635 ;
      RECT 2.86 0.085 3.03 0.545 ;
      RECT 2.86 1.835 3.03 2.635 ;
      RECT 3.7 0.085 4.005 0.545 ;
      RECT 3.7 1.835 4 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__inv_8
MACRO sky130_fd_sc_hd__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.735 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 0.255 0.895 0.725 ;
        RECT 0.565 0.725 2.17 0.905 ;
        RECT 0.565 1.495 2.17 1.665 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.405 0.255 1.735 0.725 ;
        RECT 1.405 1.665 2.17 1.685 ;
        RECT 1.405 1.685 1.735 2.465 ;
        RECT 1.905 0.905 2.17 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.13 0.085 0.395 0.545 ;
      RECT 0.13 1.495 0.395 2.635 ;
      RECT 1.065 0.085 1.235 0.545 ;
      RECT 1.065 1.835 1.235 2.635 ;
      RECT 1.905 0.085 2.155 0.55 ;
      RECT 1.905 2.175 2.115 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__inv_4
MACRO sky130_fd_sc_hd__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.775 1.325 ;
        RECT 0.085 1.325 0.4 1.765 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.643500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.665 0.255 2.215 0.545 ;
        RECT 1.765 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.285 1.965 0.565 2.635 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.245 0.085 1.495 0.545 ;
      RECT 1.245 1.915 1.575 2.635 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
      RECT 2.385 0.085 2.675 0.885 ;
      RECT 2.385 1.495 2.675 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__and2_2
MACRO sky130_fd_sc_hd__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 0.775 1.325 ;
        RECT 0.1 1.325 0.365 1.685 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 0.255 2.215 0.545 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.285 1.965 0.565 2.635 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.235 0.085 1.485 0.545 ;
      RECT 1.235 1.915 1.565 2.635 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__and2_1
MACRO sky130_fd_sc_hd__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.995 0.435 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 0.98 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.515 1.72 0.615 ;
        RECT 1.53 0.615 3.135 0.845 ;
        RECT 1.53 1.535 3.135 1.76 ;
        RECT 1.53 1.76 1.72 2.465 ;
        RECT 2.39 0.255 2.58 0.615 ;
        RECT 2.39 1.76 3.135 1.765 ;
        RECT 2.39 1.765 2.58 2.465 ;
        RECT 2.855 0.845 3.135 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.095 0.255 0.425 0.615 ;
      RECT 0.095 0.615 1.36 0.805 ;
      RECT 0.095 1.88 0.425 2.635 ;
      RECT 0.605 1.58 1.36 1.75 ;
      RECT 0.605 1.75 0.785 2.465 ;
      RECT 0.955 0.085 1.285 0.445 ;
      RECT 0.99 1.935 1.32 2.635 ;
      RECT 1.15 0.805 1.36 1.02 ;
      RECT 1.15 1.02 2.685 1.355 ;
      RECT 1.15 1.355 1.36 1.58 ;
      RECT 1.89 0.085 2.22 0.445 ;
      RECT 1.89 1.935 2.22 2.635 ;
      RECT 2.75 0.085 3.08 0.445 ;
      RECT 2.75 1.935 3.08 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__and2_4
MACRO sky130_fd_sc_hd__and2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.185 0.43 1.955 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.08 1.27 1.615 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.56 0.255 2.215 0.525 ;
        RECT 1.79 1.835 2.215 2.465 ;
        RECT 1.95 0.525 2.215 1.835 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.16 2.175 0.43 2.635 ;
      RECT 0.185 0.28 0.49 0.695 ;
      RECT 0.185 0.695 1.78 0.91 ;
      RECT 0.185 0.91 0.77 0.95 ;
      RECT 0.6 0.95 0.77 2.135 ;
      RECT 0.6 2.135 0.865 2.465 ;
      RECT 0.95 0.085 1.39 0.525 ;
      RECT 1.11 1.835 1.62 2.635 ;
      RECT 1.45 0.91 1.78 1.435 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__and2_0
MACRO sky130_fd_sc_hd__decap_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
      RECT 0.085000  1.545000 5.430000 2.635000 ;
      RECT 2.835000  1.025000 5.430000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_12
MACRO sky130_fd_sc_hd__decap_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
      RECT 0.085000  1.545000 2.675000 2.635000 ;
      RECT 1.465000  1.025000 2.675000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_6
MACRO sky130_fd_sc_hd__decap_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
      RECT 0.085000  1.545000 1.295000 2.635000 ;
      RECT 0.775000  1.005000 1.295000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_3
MACRO sky130_fd_sc_hd__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
      RECT 0.085000  1.545000 1.755000 2.635000 ;
      RECT 1.005000  1.025000 1.755000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_4
MACRO sky130_fd_sc_hd__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
      RECT 0.085000  1.545000 3.595000 2.635000 ;
      RECT 1.905000  1.025000 3.595000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_8
MACRO sky130_fd_sc_hd__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 3.1 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.39 1.075 4.5 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.78 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.485 2.16 1.655 ;
        RECT 0.095 1.655 0.345 2.465 ;
        RECT 0.935 1.655 1.265 2.125 ;
        RECT 1.355 0.675 3.045 0.845 ;
        RECT 1.775 1.655 2.16 2.125 ;
        RECT 1.87 0.845 2.16 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.095 0.255 0.345 0.68 ;
      RECT 0.095 0.68 1.185 0.85 ;
      RECT 0.515 0.085 0.845 0.51 ;
      RECT 0.515 1.825 0.765 2.295 ;
      RECT 0.515 2.295 2.625 2.465 ;
      RECT 1.015 0.255 2.105 0.505 ;
      RECT 1.015 0.505 1.185 0.68 ;
      RECT 1.435 1.825 1.605 2.295 ;
      RECT 2.295 0.255 3.385 0.505 ;
      RECT 2.375 1.485 4.305 1.655 ;
      RECT 2.375 1.655 2.625 2.295 ;
      RECT 2.795 1.825 2.965 2.635 ;
      RECT 3.135 1.655 3.465 2.465 ;
      RECT 3.215 0.505 3.385 0.68 ;
      RECT 3.215 0.68 4.375 0.85 ;
      RECT 3.555 0.085 3.885 0.51 ;
      RECT 3.635 1.825 3.805 2.635 ;
      RECT 3.975 1.655 4.305 2.465 ;
      RECT 4.055 0.255 4.375 0.68 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__a22oi_2
MACRO sky130_fd_sc_hd__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.675 1.7 1.075 ;
        RECT 1.49 1.075 1.84 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 0.995 2.335 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.275 ;
        RECT 0.99 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.575 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.445 1.84 1.495 ;
        RECT 0.095 1.495 2.675 1.625 ;
        RECT 0.095 1.625 0.425 2.295 ;
        RECT 0.095 2.295 1.265 2.465 ;
        RECT 0.82 0.255 2.125 0.505 ;
        RECT 0.935 2.255 1.265 2.295 ;
        RECT 1.615 1.625 2.675 1.665 ;
        RECT 1.945 0.505 2.125 0.655 ;
        RECT 1.945 0.655 2.675 0.825 ;
        RECT 2.505 0.825 2.675 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 0.085 0.545 0.595 ;
      RECT 0.595 1.795 1.475 1.835 ;
      RECT 0.595 1.835 2.125 2.035 ;
      RECT 0.595 2.035 1.21 2.085 ;
      RECT 0.595 2.085 0.825 2.125 ;
      RECT 1.435 2.255 1.81 2.635 ;
      RECT 1.955 2.035 2.125 2.165 ;
      RECT 2.305 0.085 2.635 0.485 ;
      RECT 2.36 1.855 2.625 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__a22oi_1
MACRO sky130_fd_sc_hd__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 5.685 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.91 1.075 7.735 1.285 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.04 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.895 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.445 3.325 1.625 ;
        RECT 0.595 1.625 0.805 2.125 ;
        RECT 1.395 1.625 1.645 2.125 ;
        RECT 2.195 0.645 5.565 0.885 ;
        RECT 2.195 0.885 2.445 1.445 ;
        RECT 2.235 1.625 2.485 2.125 ;
        RECT 3.075 1.625 3.325 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.09 1.455 0.425 2.295 ;
      RECT 0.09 2.295 4.265 2.465 ;
      RECT 0.095 0.255 0.425 0.725 ;
      RECT 0.095 0.725 2.025 0.905 ;
      RECT 0.595 0.085 0.765 0.555 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 0.975 1.795 1.225 2.295 ;
      RECT 1.435 0.085 1.605 0.555 ;
      RECT 1.775 0.255 3.785 0.475 ;
      RECT 1.775 0.475 2.025 0.725 ;
      RECT 1.815 1.795 2.065 2.295 ;
      RECT 2.655 1.795 2.905 2.295 ;
      RECT 3.495 1.455 7.625 1.625 ;
      RECT 3.495 1.625 4.265 2.295 ;
      RECT 3.975 0.255 5.985 0.475 ;
      RECT 4.435 1.795 4.685 2.635 ;
      RECT 4.855 1.625 5.105 2.465 ;
      RECT 5.275 1.795 5.525 2.635 ;
      RECT 5.695 1.625 5.945 2.465 ;
      RECT 5.735 0.475 5.985 0.725 ;
      RECT 5.735 0.725 7.665 0.905 ;
      RECT 6.115 1.795 6.365 2.635 ;
      RECT 6.155 0.085 6.325 0.555 ;
      RECT 6.495 0.255 6.825 0.725 ;
      RECT 6.535 1.625 6.785 2.465 ;
      RECT 6.955 1.795 7.205 2.635 ;
      RECT 6.995 0.085 7.165 0.555 ;
      RECT 7.335 0.255 7.665 0.725 ;
      RECT 7.375 1.625 7.625 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__a22oi_4
MACRO sky130_fd_sc_hd__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 0.955 1.77 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595 0.255 5.925 0.485 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 1.425 6.355 1.5 ;
        RECT 5.755 1.5 5.925 1.875 ;
        RECT 5.76 1.415 6.355 1.425 ;
        RECT 5.765 1.41 6.355 1.415 ;
        RECT 5.77 0.865 6.355 0.89 ;
        RECT 5.775 1.385 6.355 1.41 ;
        RECT 5.785 0.89 6.355 1.385 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.48 0.995 4.815 1.035 ;
        RECT 4.48 1.035 5.24 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.435 1.495 2.12 1.665 ;
      RECT 1.435 1.665 1.785 2.415 ;
      RECT 1.515 0.345 1.705 0.615 ;
      RECT 1.515 0.615 2.12 0.765 ;
      RECT 1.515 0.765 2.335 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.95 0.785 2.335 1.095 ;
      RECT 1.95 1.095 2.12 1.495 ;
      RECT 1.955 1.835 2.25 2.635 ;
      RECT 2.45 1.355 2.755 1.685 ;
      RECT 2.585 0.735 3.1 1.04 ;
      RECT 2.77 0.365 3.445 0.535 ;
      RECT 2.77 2.255 3.58 2.425 ;
      RECT 2.905 1.78 3.265 1.91 ;
      RECT 2.905 1.91 3.175 1.995 ;
      RECT 2.93 1.04 3.1 1.57 ;
      RECT 2.93 1.57 3.265 1.78 ;
      RECT 3.27 0.535 3.445 0.995 ;
      RECT 3.27 0.995 4.22 1.325 ;
      RECT 3.41 2 3.605 2.085 ;
      RECT 3.41 2.085 3.58 2.255 ;
      RECT 3.415 1.995 3.605 2 ;
      RECT 3.42 1.985 3.605 1.995 ;
      RECT 3.435 1.325 3.605 1.985 ;
      RECT 3.72 0.085 4.06 0.53 ;
      RECT 3.75 2.175 4.09 2.635 ;
      RECT 3.775 1.535 5.585 1.705 ;
      RECT 3.775 1.705 4.97 1.865 ;
      RECT 4.24 0.255 4.58 0.655 ;
      RECT 4.24 0.655 5.095 0.695 ;
      RECT 4.24 0.695 5.585 0.825 ;
      RECT 4.28 2.135 4.56 2.635 ;
      RECT 4.8 1.865 4.97 2.465 ;
      RECT 4.955 0.825 5.585 0.865 ;
      RECT 5.14 1.875 5.485 2.635 ;
      RECT 5.255 0.085 5.425 0.525 ;
      RECT 5.415 0.865 5.585 0.995 ;
      RECT 5.415 0.995 5.615 1.325 ;
      RECT 5.415 1.325 5.585 1.535 ;
      RECT 6.095 0.085 6.355 0.595 ;
      RECT 6.095 1.67 6.355 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.925 1.785 3.095 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.68 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.155 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_2
MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.345 5.895 0.745 ;
        RECT 5.635 1.67 5.895 2.455 ;
        RECT 5.725 0.745 5.895 1.67 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.345 4.975 0.995 ;
        RECT 4.745 0.995 5.075 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 1.795 0.775 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.775 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.775 1.07 ;
      RECT 0.605 1.07 0.835 1.4 ;
      RECT 0.605 1.4 0.775 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.235 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.785 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.115 0.765 ;
      RECT 1.51 0.765 2.335 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.945 0.785 2.335 1.095 ;
      RECT 1.945 1.095 2.115 1.495 ;
      RECT 1.955 1.835 2.245 2.635 ;
      RECT 2.445 1.355 2.835 1.625 ;
      RECT 2.445 1.625 2.76 1.685 ;
      RECT 2.69 0.765 3.245 1.095 ;
      RECT 2.81 2.255 3.625 2.425 ;
      RECT 2.815 0.365 3.585 0.535 ;
      RECT 2.9 1.785 3.265 1.995 ;
      RECT 3.005 1.095 3.245 1.635 ;
      RECT 3.005 1.635 3.265 1.785 ;
      RECT 3.415 0.535 3.585 0.995 ;
      RECT 3.415 0.995 4.175 1.165 ;
      RECT 3.455 1.165 4.175 1.325 ;
      RECT 3.455 1.325 3.625 2.255 ;
      RECT 3.755 0.085 4.025 0.61 ;
      RECT 3.815 1.535 5.465 1.735 ;
      RECT 3.815 1.735 4.965 1.865 ;
      RECT 3.93 2.135 4.445 2.635 ;
      RECT 4.195 0.295 4.575 0.805 ;
      RECT 4.345 0.805 4.575 1.505 ;
      RECT 4.345 1.505 5.465 1.535 ;
      RECT 4.625 1.865 4.965 2.435 ;
      RECT 5.135 1.915 5.465 2.635 ;
      RECT 5.155 0.085 5.44 0.715 ;
      RECT 5.245 0.995 5.555 1.325 ;
      RECT 5.245 1.325 5.465 1.505 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 1.445 0.775 1.615 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.445 2.615 1.615 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.925 1.785 3.095 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 0.545 1.415 0.835 1.46 ;
      RECT 0.545 1.46 2.675 1.6 ;
      RECT 0.545 1.6 0.835 1.645 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 3.155 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.385 1.415 2.675 1.46 ;
      RECT 2.385 1.6 2.675 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_1
MACRO sky130_fd_sc_hd__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.255 5.965 0.485 ;
        RECT 5.68 1.875 5.965 2.465 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 0.255 6.775 0.765 ;
        RECT 6.575 1.325 6.775 2.465 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.96 1.835 2.275 2.635 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.46 1.495 2.145 1.665 ;
      RECT 1.46 1.665 1.79 2.415 ;
      RECT 1.54 0.345 1.71 0.615 ;
      RECT 1.54 0.615 2.145 0.765 ;
      RECT 1.54 0.765 2.345 0.785 ;
      RECT 1.88 0.085 2.21 0.445 ;
      RECT 1.975 0.785 2.345 1.095 ;
      RECT 1.975 1.095 2.145 1.495 ;
      RECT 2.475 1.355 2.76 1.685 ;
      RECT 2.72 0.705 3.1 1.035 ;
      RECT 2.845 0.365 3.505 0.535 ;
      RECT 2.905 2.255 3.655 2.425 ;
      RECT 2.93 1.035 3.1 1.575 ;
      RECT 2.93 1.575 3.27 1.995 ;
      RECT 3.335 0.535 3.505 0.995 ;
      RECT 3.335 0.995 4.235 1.165 ;
      RECT 3.485 1.165 4.235 1.325 ;
      RECT 3.485 1.325 3.655 2.255 ;
      RECT 3.745 0.085 4.075 0.53 ;
      RECT 3.825 1.535 5.625 1.705 ;
      RECT 3.825 1.705 4.945 1.865 ;
      RECT 4.265 0.255 4.595 0.655 ;
      RECT 4.265 0.655 5.625 0.825 ;
      RECT 4.755 1.865 4.945 2.465 ;
      RECT 5.1 0.085 5.44 0.485 ;
      RECT 5.455 0.825 5.625 1.535 ;
      RECT 6.135 0.085 6.405 0.595 ;
      RECT 6.945 0.085 7.275 0.595 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.475 1.445 2.645 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.935 1.785 3.105 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.705 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.165 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.415 1.415 2.705 1.46 ;
      RECT 2.415 1.6 2.705 1.645 ;
      RECT 2.875 1.755 3.165 1.8 ;
      RECT 2.875 1.94 3.165 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_4
MACRO sky130_fd_sc_hd__lpflow_inputiso0n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 0.775 1.325 ;
        RECT 0.1 1.325 0.365 1.685 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 0.255 2.215 0.545 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.285 1.965 0.565 2.635 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.235 0.085 1.485 0.545 ;
      RECT 1.235 1.915 1.565 2.635 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0n_1
MACRO sky130_fd_sc_hd__maj3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.125 1.325 ;
        RECT 0.61 1.325 0.78 2.46 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.995 1.905 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.765 2.755 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.602250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255 0.255 3.595 0.825 ;
        RECT 3.255 2.16 3.595 2.465 ;
        RECT 3.265 1.495 3.595 2.16 ;
        RECT 3.37 0.825 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.135 0.255 0.395 0.655 ;
      RECT 0.135 0.655 2.245 0.825 ;
      RECT 0.135 0.825 0.395 2.125 ;
      RECT 0.875 0.085 1.205 0.485 ;
      RECT 0.955 1.715 1.205 2.635 ;
      RECT 1.655 0.255 1.985 0.64 ;
      RECT 1.655 0.64 2.245 0.655 ;
      RECT 1.655 1.815 2.245 2.08 ;
      RECT 2.075 0.825 2.245 1.495 ;
      RECT 2.075 1.495 3.095 1.665 ;
      RECT 2.075 1.665 2.245 1.815 ;
      RECT 2.545 0.085 2.88 0.47 ;
      RECT 2.555 1.845 2.885 2.635 ;
      RECT 2.925 0.995 3.2 1.325 ;
      RECT 2.925 1.325 3.095 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__maj3_1
MACRO sky130_fd_sc_hd__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.45 1.635 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 1.075 2.29 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.89 1.285 ;
        RECT 0.72 1.285 0.89 1.915 ;
        RECT 0.72 1.915 1.79 2.085 ;
        RECT 1.62 2.085 1.79 2.225 ;
        RECT 1.62 2.225 2.63 2.395 ;
        RECT 2.46 1.075 2.945 1.245 ;
        RECT 2.46 1.245 2.63 2.225 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375 0.255 3.705 0.49 ;
        RECT 3.375 1.455 4.975 1.625 ;
        RECT 3.375 1.625 3.705 2.465 ;
        RECT 3.455 0.49 3.705 0.715 ;
        RECT 3.455 0.715 4.975 0.905 ;
        RECT 4.215 0.255 4.545 0.715 ;
        RECT 4.215 1.625 4.545 2.465 ;
        RECT 4.715 0.905 4.975 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.255 0.635 0.66 ;
      RECT 0.085 0.66 2.29 0.715 ;
      RECT 0.085 0.715 3.285 0.885 ;
      RECT 0.085 0.885 0.255 1.455 ;
      RECT 0.085 1.455 0.465 2.465 ;
      RECT 1.12 0.085 1.45 0.49 ;
      RECT 1.12 2.255 1.45 2.635 ;
      RECT 1.62 0.885 1.79 1.545 ;
      RECT 1.62 1.545 2.29 1.745 ;
      RECT 1.96 0.255 2.29 0.66 ;
      RECT 1.96 1.745 2.29 2.055 ;
      RECT 2.845 1.455 3.175 2.635 ;
      RECT 2.86 0.085 3.205 0.545 ;
      RECT 3.115 0.885 3.285 1.075 ;
      RECT 3.115 1.075 4.545 1.285 ;
      RECT 3.875 0.085 4.045 0.545 ;
      RECT 3.875 1.795 4.045 2.635 ;
      RECT 4.715 0.085 4.885 0.545 ;
      RECT 4.715 1.795 4.925 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__maj3_4
MACRO sky130_fd_sc_hd__maj3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 0.995 1.695 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865 0.995 2.155 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.495 ;
        RECT 0.425 1.495 3.07 1.665 ;
        RECT 2.415 1.415 3.07 1.495 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285 0.255 3.615 0.905 ;
        RECT 3.285 1.495 3.615 2.465 ;
        RECT 3.445 0.905 3.615 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.28 0.525 0.655 ;
      RECT 0.085 0.655 3.105 0.825 ;
      RECT 0.085 0.825 0.255 1.835 ;
      RECT 0.085 1.835 2.085 2.005 ;
      RECT 0.085 2.005 0.615 2.465 ;
      RECT 0.975 0.085 1.305 0.485 ;
      RECT 0.975 2.175 1.305 2.635 ;
      RECT 1.755 0.255 2.085 0.655 ;
      RECT 1.755 2.005 2.085 2.465 ;
      RECT 2.535 1.835 2.86 2.635 ;
      RECT 2.635 0.085 2.965 0.485 ;
      RECT 2.925 0.825 3.105 1.075 ;
      RECT 2.925 1.075 3.275 1.245 ;
      RECT 3.785 0.085 4.055 0.905 ;
      RECT 3.785 1.495 4.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__maj3_2
MACRO sky130_fd_sc_hd__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 3.56 1.275 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.31 0.995 4.635 1.615 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.325 ;
        RECT 0.58 0.725 0.78 0.995 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.691250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.295 4.975 0.465 ;
        RECT 2.715 2.255 4.975 2.425 ;
        RECT 4.75 1.785 4.975 2.255 ;
        RECT 4.805 0.465 4.975 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.345 0.345 0.675 ;
      RECT 0.085 0.675 0.26 1.495 ;
      RECT 0.085 1.495 1.395 1.665 ;
      RECT 0.085 1.665 0.26 2.135 ;
      RECT 0.085 2.135 0.345 2.465 ;
      RECT 0.515 0.085 0.835 0.545 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 0.935 1.835 1.735 2.005 ;
      RECT 1.015 0.575 1.255 0.935 ;
      RECT 1.225 1.155 1.985 1.325 ;
      RECT 1.225 1.325 1.395 1.495 ;
      RECT 1.355 2.255 1.685 2.635 ;
      RECT 1.435 0.085 1.685 0.885 ;
      RECT 1.565 1.495 3.465 1.665 ;
      RECT 1.565 1.665 1.735 1.835 ;
      RECT 1.655 1.075 1.985 1.155 ;
      RECT 1.855 0.295 2.025 0.735 ;
      RECT 1.855 0.735 3.465 0.905 ;
      RECT 1.855 2.135 2.08 2.465 ;
      RECT 1.91 1.835 2.885 1.915 ;
      RECT 1.91 1.915 4.35 2.005 ;
      RECT 1.91 2.005 2.08 2.135 ;
      RECT 2.275 0.085 2.445 0.545 ;
      RECT 2.275 2.175 2.525 2.635 ;
      RECT 2.715 2.005 4.35 2.085 ;
      RECT 3.135 0.655 3.465 0.735 ;
      RECT 3.135 1.665 3.465 1.715 ;
      RECT 3.85 0.655 4.345 0.825 ;
      RECT 3.85 0.825 4.105 0.935 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.85 0.765 4.02 0.935 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
    LAYER met1 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 4.08 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 3.79 0.735 4.08 0.78 ;
      RECT 3.79 0.92 4.08 0.965 ;
  END
END sky130_fd_sc_hd__mux2i_2
MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.995 1.07 1.105 ;
        RECT 0.56 1.105 1.24 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 3.55 1.325 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.237500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845 1.075 5.93 1.29 ;
        RECT 5.76 1.29 5.93 1.425 ;
        RECT 5.76 1.425 7.85 1.595 ;
        RECT 7.68 0.995 7.85 1.425 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.194500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.315 3.785 0.485 ;
        RECT 0.095 0.485 0.32 2.255 ;
        RECT 0.095 2.255 3.785 2.425 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.515 0.655 1.7 0.825 ;
      RECT 0.515 1.575 5.58 1.745 ;
      RECT 1.355 0.825 1.7 0.935 ;
      RECT 2.195 0.655 5.485 0.825 ;
      RECT 2.195 1.915 7.165 2.085 ;
      RECT 3.975 0.085 4.305 0.465 ;
      RECT 3.975 2.255 4.305 2.635 ;
      RECT 4.475 0.255 4.645 0.655 ;
      RECT 4.815 0.085 5.145 0.465 ;
      RECT 4.815 2.255 5.145 2.635 ;
      RECT 5.315 0.255 5.485 0.655 ;
      RECT 5.655 0.085 5.98 0.59 ;
      RECT 5.655 2.255 5.985 2.635 ;
      RECT 6.15 0.255 6.325 0.715 ;
      RECT 6.15 0.715 7.165 0.905 ;
      RECT 6.15 0.905 6.45 0.935 ;
      RECT 6.155 1.795 6.325 1.915 ;
      RECT 6.155 2.085 6.325 2.465 ;
      RECT 6.495 2.255 6.825 2.635 ;
      RECT 6.545 0.085 6.795 0.545 ;
      RECT 6.73 1.075 7.51 1.245 ;
      RECT 6.995 0.51 7.165 0.715 ;
      RECT 6.995 1.795 7.165 1.915 ;
      RECT 6.995 2.085 7.165 2.465 ;
      RECT 7.34 0.655 8.195 0.825 ;
      RECT 7.34 0.825 7.51 1.075 ;
      RECT 7.435 0.085 7.765 0.465 ;
      RECT 7.435 2.255 7.765 2.635 ;
      RECT 7.935 0.255 8.195 0.655 ;
      RECT 7.935 1.795 8.195 2.465 ;
      RECT 8.02 0.825 8.195 1.795 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.15 0.765 6.32 0.935 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 6.38 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 6.09 0.735 6.38 0.78 ;
      RECT 6.09 0.92 6.38 0.965 ;
  END
END sky130_fd_sc_hd__mux2i_4
MACRO sky130_fd_sc_hd__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.06 0.42 1.285 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.995 1.125 1.155 ;
        RECT 0.955 1.155 1.205 1.325 ;
        RECT 1.035 1.325 1.205 1.445 ;
        RECT 1.035 1.445 1.235 2.11 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 0.76 3.595 1.62 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.595 0.78 1.455 ;
        RECT 0.59 1.455 0.84 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.255 1.805 0.425 ;
      RECT 0.085 0.425 0.44 0.465 ;
      RECT 0.085 0.465 0.345 0.885 ;
      RECT 0.12 1.455 0.42 2.295 ;
      RECT 0.12 2.295 1.575 2.465 ;
      RECT 0.955 0.655 1.52 0.715 ;
      RECT 0.955 0.715 2.62 0.825 ;
      RECT 0.965 0.425 1.805 0.465 ;
      RECT 1.295 0.825 2.62 0.885 ;
      RECT 1.385 1.075 3.085 1.31 ;
      RECT 1.405 1.48 2.615 1.65 ;
      RECT 1.405 1.65 1.575 2.295 ;
      RECT 1.745 1.835 1.975 2.635 ;
      RECT 1.975 0.085 2.145 0.545 ;
      RECT 2.285 1.65 2.615 2.465 ;
      RECT 2.385 0.255 2.62 0.715 ;
      RECT 2.8 0.255 3.165 0.485 ;
      RECT 2.8 0.485 3.085 1.075 ;
      RECT 2.86 1.31 3.085 2.465 ;
      RECT 3.295 1.835 3.59 2.635 ;
      RECT 3.335 0.085 3.555 0.545 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__mux2i_1
MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.95 1.055 7.735 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.02 1.055 6.77 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655 1.055 5.85 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 1.055 4.475 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.115 1.055 3.08 1.315 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.765 1.315 ;
        RECT 0.595 0.255 0.765 0.715 ;
        RECT 0.595 0.715 1.605 0.885 ;
        RECT 0.595 0.885 0.765 1.055 ;
        RECT 0.595 1.315 0.765 1.485 ;
        RECT 0.595 1.485 1.605 1.725 ;
        RECT 0.595 1.725 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.715 ;
        RECT 1.435 1.725 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.085 0.085 0.425 0.885 ;
      RECT 0.085 1.485 0.425 2.635 ;
      RECT 0.935 0.085 1.265 0.545 ;
      RECT 0.935 1.055 1.945 1.315 ;
      RECT 0.935 1.895 1.265 2.635 ;
      RECT 1.775 0.085 2.025 0.545 ;
      RECT 1.775 0.715 3.045 0.885 ;
      RECT 1.775 0.885 1.945 1.055 ;
      RECT 1.775 1.315 1.945 1.485 ;
      RECT 1.775 1.485 5.005 1.725 ;
      RECT 1.775 1.895 2.445 2.635 ;
      RECT 2.195 0.255 4.305 0.505 ;
      RECT 2.195 0.675 3.045 0.715 ;
      RECT 2.615 1.725 2.785 2.465 ;
      RECT 2.955 1.895 3.285 2.635 ;
      RECT 3.215 0.505 3.385 0.885 ;
      RECT 3.455 1.725 3.625 2.465 ;
      RECT 3.555 0.675 7.735 0.885 ;
      RECT 3.855 1.895 4.045 2.635 ;
      RECT 4.335 1.895 4.665 2.295 ;
      RECT 4.335 2.295 6.445 2.465 ;
      RECT 4.485 0.255 4.755 0.675 ;
      RECT 4.835 1.725 5.005 2.125 ;
      RECT 4.925 0.085 5.605 0.505 ;
      RECT 5.255 1.485 5.525 2.295 ;
      RECT 5.695 1.485 7.735 1.725 ;
      RECT 5.695 1.725 5.945 2.125 ;
      RECT 5.775 0.255 5.945 0.675 ;
      RECT 6.115 0.085 6.445 0.505 ;
      RECT 6.115 1.895 6.445 2.295 ;
      RECT 6.615 0.255 6.785 0.675 ;
      RECT 6.615 1.725 6.785 2.125 ;
      RECT 6.955 0.085 7.285 0.505 ;
      RECT 6.955 1.895 7.285 2.635 ;
      RECT 7.455 0.255 7.735 0.675 ;
      RECT 7.455 1.725 7.735 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__o311a_4
MACRO sky130_fd_sc_hd__o311a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.28 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.45 0.995 1.79 1.325 ;
        RECT 1.52 1.325 1.79 2.07 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 0.995 2.27 1.325 ;
        RECT 1.98 1.325 2.215 2.07 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.84 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.995 3.595 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.355 1.07 ;
        RECT 0.085 1.07 0.435 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.525 0.085 1.195 0.825 ;
      RECT 0.605 0.995 0.775 1.495 ;
      RECT 0.605 1.495 1.35 1.665 ;
      RECT 0.605 1.835 1.01 2.635 ;
      RECT 1.18 1.665 1.35 2.295 ;
      RECT 1.18 2.295 2.715 2.465 ;
      RECT 1.365 0.31 1.66 0.655 ;
      RECT 1.365 0.655 2.76 0.825 ;
      RECT 1.84 0.085 2.215 0.485 ;
      RECT 2.385 1.495 3.595 1.665 ;
      RECT 2.385 1.665 2.715 2.295 ;
      RECT 2.43 0.31 2.76 0.655 ;
      RECT 2.9 1.835 3.135 2.635 ;
      RECT 3.01 0.255 3.595 0.825 ;
      RECT 3.01 0.825 3.18 1.495 ;
      RECT 3.305 1.665 3.595 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o311a_1
MACRO sky130_fd_sc_hd__o311a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.75 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.92 0.995 2.25 1.325 ;
        RECT 1.98 1.325 2.25 2.07 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.73 1.325 ;
        RECT 2.44 1.325 2.675 2.07 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.995 3.3 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.81 0.995 4.055 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.905 1.315 ;
        RECT 0.55 0.255 0.825 0.995 ;
        RECT 0.55 0.995 0.905 1.055 ;
        RECT 0.55 1.315 0.905 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.085 0.38 0.885 ;
      RECT 0.085 1.485 0.38 2.635 ;
      RECT 0.995 0.085 1.665 0.825 ;
      RECT 1.075 0.995 1.245 1.495 ;
      RECT 1.075 1.495 1.81 1.665 ;
      RECT 1.075 1.835 1.47 2.635 ;
      RECT 1.64 1.665 1.81 2.295 ;
      RECT 1.64 2.295 3.175 2.465 ;
      RECT 1.835 0.31 2.12 0.655 ;
      RECT 1.835 0.655 3.22 0.825 ;
      RECT 2.3 0.085 2.675 0.485 ;
      RECT 2.845 1.495 4.055 1.665 ;
      RECT 2.845 1.665 3.175 2.295 ;
      RECT 2.89 0.31 3.22 0.655 ;
      RECT 3.36 1.835 3.595 2.635 ;
      RECT 3.47 0.255 4.055 0.825 ;
      RECT 3.47 0.825 3.64 1.495 ;
      RECT 3.765 1.665 4.055 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o311a_2
MACRO sky130_fd_sc_hd__macro_sparecell
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__macro_sparecell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN LO
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215 1.075 4.965 1.325 ;
      LAYER mcon ;
        RECT 4.775 1.105 4.945 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.135 1.075 5.895 1.325 ;
      LAYER mcon ;
        RECT 5.705 1.105 5.875 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.755 0.915 7.275 2.465 ;
      LAYER mcon ;
        RECT 6.765 1.105 6.935 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.445 1.075 8.205 1.325 ;
      LAYER mcon ;
        RECT 7.625 1.105 7.795 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.375 1.075 9.125 1.325 ;
      LAYER mcon ;
        RECT 8.485 1.105 8.655 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.715 1.075 5.005 1.12 ;
        RECT 4.715 1.12 8.715 1.26 ;
        RECT 4.715 1.26 5.005 1.305 ;
        RECT 5.645 1.075 5.935 1.12 ;
        RECT 5.645 1.26 5.935 1.305 ;
        RECT 6.705 1.075 6.995 1.12 ;
        RECT 6.705 1.26 6.995 1.305 ;
        RECT 7.565 1.075 7.855 1.12 ;
        RECT 7.565 1.26 7.855 1.305 ;
        RECT 8.425 1.075 8.715 1.12 ;
        RECT 8.425 1.26 8.715 1.305 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.34 0.085 ;
        RECT 0.145 0.085 0.355 0.905 ;
        RECT 1.025 0.085 1.255 0.905 ;
        RECT 1.515 0.085 1.805 0.555 ;
        RECT 2.475 0.085 2.645 0.555 ;
        RECT 3.315 0.085 3.59 0.905 ;
        RECT 5.215 0.085 5.385 0.545 ;
        RECT 6.755 0.085 7.095 0.745 ;
        RECT 7.955 0.085 8.125 0.545 ;
        RECT 9.75 0.085 10.025 0.905 ;
        RECT 10.695 0.085 10.865 0.555 ;
        RECT 11.535 0.085 11.825 0.555 ;
        RECT 12.085 0.085 12.315 0.905 ;
        RECT 12.985 0.085 13.195 0.905 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 13.53 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.34 2.805 ;
        RECT 0.145 1.495 0.355 2.635 ;
        RECT 1.025 1.495 1.255 2.635 ;
        RECT 2.815 1.835 3.145 2.635 ;
        RECT 3.87 1.835 4.125 2.635 ;
        RECT 4.795 1.835 4.965 2.635 ;
        RECT 5.635 1.495 5.895 2.635 ;
        RECT 6.255 1.91 6.585 2.635 ;
        RECT 7.445 1.495 7.705 2.635 ;
        RECT 8.375 1.835 8.545 2.635 ;
        RECT 9.215 1.835 9.47 2.635 ;
        RECT 10.195 1.835 10.525 2.635 ;
        RECT 12.085 1.495 12.315 2.635 ;
        RECT 12.985 1.495 13.195 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 0.255 0.855 0.885 ;
      RECT 0.525 0.885 0.775 1.485 ;
      RECT 0.525 1.485 0.855 2.465 ;
      RECT 0.945 1.075 1.275 1.325 ;
      RECT 1.505 1.835 1.805 2.295 ;
      RECT 1.505 2.295 2.645 2.465 ;
      RECT 1.545 0.735 3.145 0.905 ;
      RECT 1.545 0.905 1.76 1.445 ;
      RECT 1.545 1.445 2.305 1.665 ;
      RECT 1.93 1.075 2.7 1.275 ;
      RECT 1.975 0.255 2.305 0.725 ;
      RECT 1.975 0.725 3.145 0.735 ;
      RECT 1.975 1.665 2.305 2.125 ;
      RECT 2.475 1.455 3.59 1.665 ;
      RECT 2.475 1.665 2.645 2.295 ;
      RECT 2.815 0.255 3.145 0.725 ;
      RECT 2.87 1.075 3.59 1.275 ;
      RECT 3.315 1.665 3.59 2.465 ;
      RECT 3.765 0.655 4.625 0.905 ;
      RECT 3.765 0.905 4.045 1.495 ;
      RECT 3.765 1.495 5.465 1.665 ;
      RECT 3.875 0.255 5.045 0.465 ;
      RECT 3.875 0.465 4.205 0.485 ;
      RECT 4.295 1.665 4.625 2.465 ;
      RECT 4.795 0.465 5.045 0.715 ;
      RECT 4.795 0.715 5.895 0.885 ;
      RECT 5.135 1.665 5.465 2.465 ;
      RECT 5.555 0.255 5.895 0.715 ;
      RECT 6.065 0.255 6.585 1.74 ;
      RECT 7.445 0.255 7.785 0.715 ;
      RECT 7.445 0.715 8.545 0.885 ;
      RECT 7.875 1.495 9.575 1.665 ;
      RECT 7.875 1.665 8.205 2.465 ;
      RECT 8.295 0.255 9.465 0.465 ;
      RECT 8.295 0.465 8.545 0.715 ;
      RECT 8.715 0.655 9.575 0.905 ;
      RECT 8.715 1.665 9.045 2.465 ;
      RECT 9.135 0.465 9.465 0.485 ;
      RECT 9.295 0.905 9.575 1.495 ;
      RECT 9.75 1.075 10.47 1.275 ;
      RECT 9.75 1.455 10.865 1.665 ;
      RECT 9.75 1.665 10.025 2.465 ;
      RECT 10.195 0.255 10.525 0.725 ;
      RECT 10.195 0.725 11.365 0.735 ;
      RECT 10.195 0.735 11.795 0.905 ;
      RECT 10.64 1.075 11.41 1.275 ;
      RECT 10.695 1.665 10.865 2.295 ;
      RECT 10.695 2.295 11.835 2.465 ;
      RECT 11.035 0.255 11.365 0.725 ;
      RECT 11.035 1.445 11.795 1.665 ;
      RECT 11.035 1.665 11.365 2.125 ;
      RECT 11.535 1.835 11.835 2.295 ;
      RECT 11.58 0.905 11.795 1.445 ;
      RECT 12.065 1.075 12.395 1.325 ;
      RECT 12.485 0.255 12.815 0.885 ;
      RECT 12.485 1.485 12.815 2.465 ;
      RECT 12.565 0.885 12.815 1.485 ;
    LAYER mcon ;
      RECT 0.565 1.105 0.735 1.275 ;
      RECT 1.085 1.105 1.255 1.275 ;
      RECT 1.57 1.105 1.74 1.275 ;
      RECT 2.1 1.105 2.27 1.275 ;
      RECT 2.96 1.105 3.13 1.275 ;
      RECT 3.82 1.105 3.99 1.275 ;
      RECT 9.345 1.105 9.515 1.275 ;
      RECT 10.205 1.105 10.375 1.275 ;
      RECT 11.065 1.105 11.235 1.275 ;
      RECT 11.605 1.105 11.775 1.275 ;
      RECT 12.09 1.105 12.26 1.275 ;
      RECT 12.605 1.105 12.775 1.275 ;
    LAYER met1 ;
      RECT 0.505 1.075 0.875 1.305 ;
      RECT 1.025 1.075 1.315 1.12 ;
      RECT 1.025 1.12 1.8 1.26 ;
      RECT 1.025 1.26 1.315 1.305 ;
      RECT 1.51 1.075 1.8 1.12 ;
      RECT 1.51 1.26 1.8 1.305 ;
      RECT 2.04 1.075 2.33 1.12 ;
      RECT 2.04 1.12 4.05 1.26 ;
      RECT 2.04 1.26 2.33 1.305 ;
      RECT 2.9 1.075 3.19 1.12 ;
      RECT 2.9 1.26 3.19 1.305 ;
      RECT 3.76 1.075 4.05 1.12 ;
      RECT 3.76 1.26 4.05 1.305 ;
      RECT 9.285 1.075 9.575 1.12 ;
      RECT 9.285 1.12 11.295 1.26 ;
      RECT 9.285 1.26 9.575 1.305 ;
      RECT 10.145 1.075 10.435 1.12 ;
      RECT 10.145 1.26 10.435 1.305 ;
      RECT 11.005 1.075 11.295 1.12 ;
      RECT 11.005 1.26 11.295 1.305 ;
      RECT 11.545 1.075 11.835 1.12 ;
      RECT 11.545 1.12 12.32 1.26 ;
      RECT 11.545 1.26 11.835 1.305 ;
      RECT 12.03 1.075 12.32 1.12 ;
      RECT 12.03 1.26 12.32 1.305 ;
      RECT 12.47 1.075 12.835 1.305 ;
    LAYER pwell ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 3.36 -0.085 3.53 0.085 ;
      RECT 5.66 -0.085 5.83 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 7.51 -0.085 7.68 0.085 ;
      RECT 9.81 -0.085 9.98 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
  END
END sky130_fd_sc_hd__macro_sparecell
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.725 0.325 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 1.065 1.325 1.325 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235 0.255 1.565 0.725 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.655 1.85 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.85 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.33 0.37 0.675 0.545 ;
      RECT 0.415 1.51 1.705 1.68 ;
      RECT 0.415 1.68 0.675 1.905 ;
      RECT 0.495 0.545 0.675 1.51 ;
      RECT 0.855 0.085 1.065 0.895 ;
      RECT 0.875 1.855 1.205 2.635 ;
      RECT 1.535 1.075 1.865 1.245 ;
      RECT 1.535 1.245 1.705 1.51 ;
      RECT 1.735 0.085 2.12 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 20.24 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.315 0.995 ;
        RECT 0.085 0.995 0.665 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.45 1.075 15.65 1.285 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.255 3.255 0.725 ;
        RECT 2.925 0.725 16.475 0.905 ;
        RECT 3.765 0.255 4.095 0.725 ;
        RECT 4.605 0.255 4.935 0.725 ;
        RECT 5.445 0.255 5.775 0.725 ;
        RECT 6.285 0.255 6.615 0.725 ;
        RECT 7.125 0.255 7.455 0.725 ;
        RECT 7.965 0.255 8.295 0.725 ;
        RECT 8.805 0.255 9.135 0.725 ;
        RECT 9.645 0.255 9.975 0.725 ;
        RECT 9.685 1.455 16.475 1.625 ;
        RECT 9.685 1.625 9.935 2.125 ;
        RECT 10.485 0.255 10.815 0.725 ;
        RECT 10.525 1.625 10.775 2.125 ;
        RECT 11.325 0.255 11.655 0.725 ;
        RECT 11.365 1.625 11.615 2.125 ;
        RECT 12.165 0.255 12.495 0.725 ;
        RECT 12.205 1.625 12.455 2.125 ;
        RECT 13.005 0.255 13.335 0.725 ;
        RECT 13.045 1.625 13.295 2.125 ;
        RECT 13.845 0.255 14.175 0.725 ;
        RECT 13.885 1.625 14.135 2.125 ;
        RECT 14.685 0.255 15.015 0.725 ;
        RECT 14.725 1.625 14.975 2.125 ;
        RECT 15.525 0.255 15.855 0.725 ;
        RECT 15.565 1.625 15.815 2.125 ;
        RECT 15.82 0.905 16.475 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 16.56 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 16.75 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 16.56 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 16.56 0.085 ;
      RECT 0 2.635 16.56 2.805 ;
      RECT 0.3 1.495 0.515 2.635 ;
      RECT 0.485 0.085 0.815 0.825 ;
      RECT 0.685 1.495 1.015 2.465 ;
      RECT 0.835 1.065 2.035 1.075 ;
      RECT 0.835 1.075 9.28 1.285 ;
      RECT 0.835 1.285 1.015 1.495 ;
      RECT 0.985 0.255 1.195 1.065 ;
      RECT 1.185 1.455 1.355 2.635 ;
      RECT 1.365 0.085 1.615 0.895 ;
      RECT 1.525 1.285 1.855 2.465 ;
      RECT 1.785 0.255 2.035 1.065 ;
      RECT 2.025 1.455 2.27 2.635 ;
      RECT 2.205 0.085 2.755 0.905 ;
      RECT 2.475 1.455 9.515 1.665 ;
      RECT 2.475 1.665 2.795 2.465 ;
      RECT 2.965 1.835 3.215 2.635 ;
      RECT 3.385 1.665 3.635 2.465 ;
      RECT 3.425 0.085 3.595 0.555 ;
      RECT 3.805 1.835 4.055 2.635 ;
      RECT 4.225 1.665 4.475 2.465 ;
      RECT 4.265 0.085 4.435 0.555 ;
      RECT 4.645 1.835 4.895 2.635 ;
      RECT 5.065 1.665 5.315 2.465 ;
      RECT 5.105 0.085 5.275 0.555 ;
      RECT 5.485 1.835 5.735 2.635 ;
      RECT 5.905 1.665 6.155 2.465 ;
      RECT 5.945 0.085 6.115 0.555 ;
      RECT 6.325 1.835 6.575 2.635 ;
      RECT 6.745 1.665 6.995 2.465 ;
      RECT 6.785 0.085 6.955 0.555 ;
      RECT 7.165 1.835 7.415 2.635 ;
      RECT 7.585 1.665 7.835 2.465 ;
      RECT 7.625 0.085 7.795 0.555 ;
      RECT 8.005 1.835 8.255 2.635 ;
      RECT 8.425 1.665 8.675 2.465 ;
      RECT 8.465 0.085 8.635 0.555 ;
      RECT 8.845 1.835 9.095 2.635 ;
      RECT 9.265 1.665 9.515 2.295 ;
      RECT 9.265 2.295 16.235 2.465 ;
      RECT 9.305 0.085 9.475 0.555 ;
      RECT 10.105 1.795 10.355 2.295 ;
      RECT 10.145 0.085 10.315 0.555 ;
      RECT 10.945 1.795 11.195 2.295 ;
      RECT 10.985 0.085 11.155 0.555 ;
      RECT 11.785 1.795 12.035 2.295 ;
      RECT 11.825 0.085 11.995 0.555 ;
      RECT 12.625 1.795 12.875 2.295 ;
      RECT 12.665 0.085 12.835 0.555 ;
      RECT 13.465 1.795 13.715 2.295 ;
      RECT 13.505 0.085 13.675 0.555 ;
      RECT 14.305 1.795 14.555 2.295 ;
      RECT 14.345 0.085 14.515 0.555 ;
      RECT 15.145 1.795 15.395 2.295 ;
      RECT 15.185 0.085 15.355 0.555 ;
      RECT 15.985 1.795 16.235 2.295 ;
      RECT 16.025 0.085 16.295 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 14.405 2.635 14.575 2.805 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.865 2.635 15.035 2.805 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 15.325 2.635 15.495 2.805 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.785 2.635 15.955 2.805 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 16.245 2.635 16.415 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.065 3.125 1.275 ;
        RECT 2.91 1.275 3.125 1.965 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.48 1.065 0.92 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 0.895 1.665 2.125 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.365 0.895 ;
      RECT 0.085 1.445 1.245 1.655 ;
      RECT 0.085 1.655 0.405 2.465 ;
      RECT 0.575 1.825 0.825 2.635 ;
      RECT 0.995 1.655 1.245 2.295 ;
      RECT 0.995 2.295 2.125 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.835 1.445 2.09 1.89 ;
      RECT 1.835 1.89 2.125 2.295 ;
      RECT 1.875 0.085 2.045 0.895 ;
      RECT 1.875 1.075 2.43 1.245 ;
      RECT 2.215 0.725 2.565 0.895 ;
      RECT 2.215 0.895 2.43 1.075 ;
      RECT 2.26 1.245 2.43 1.445 ;
      RECT 2.26 1.445 2.565 1.615 ;
      RECT 2.395 0.445 2.565 0.725 ;
      RECT 2.395 1.615 2.565 2.46 ;
      RECT 2.775 0.085 3.03 0.845 ;
      RECT 2.775 2.145 3.025 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_2
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.265 1.065 ;
        RECT 0.085 1.065 0.575 1.285 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.27 1.075 8.01 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.255 2.335 0.725 ;
        RECT 2.005 0.725 8.655 0.905 ;
        RECT 2.845 0.255 3.175 0.725 ;
        RECT 3.685 0.255 4.015 0.725 ;
        RECT 4.525 0.255 4.855 0.725 ;
        RECT 5.365 0.255 5.695 0.725 ;
        RECT 5.405 1.445 8.655 1.615 ;
        RECT 5.405 1.615 5.655 2.125 ;
        RECT 6.205 0.255 6.535 0.725 ;
        RECT 6.245 1.615 6.495 2.125 ;
        RECT 7.045 0.255 7.375 0.725 ;
        RECT 7.085 1.615 7.335 2.125 ;
        RECT 7.885 0.255 8.215 0.725 ;
        RECT 7.925 1.615 8.175 2.125 ;
        RECT 8.18 0.905 8.655 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.195 1.455 0.415 2.635 ;
      RECT 0.435 0.085 0.655 0.895 ;
      RECT 0.585 1.455 0.915 2.465 ;
      RECT 0.745 1.065 1.155 1.075 ;
      RECT 0.745 1.075 5 1.285 ;
      RECT 0.745 1.285 0.915 1.455 ;
      RECT 0.825 0.255 1.155 1.065 ;
      RECT 1.085 1.455 1.33 2.635 ;
      RECT 1.325 0.085 1.835 0.905 ;
      RECT 1.555 1.455 5.235 1.665 ;
      RECT 1.555 1.665 1.875 2.465 ;
      RECT 2.045 1.835 2.295 2.635 ;
      RECT 2.465 1.665 2.715 2.465 ;
      RECT 2.505 0.085 2.675 0.555 ;
      RECT 2.885 1.835 3.135 2.635 ;
      RECT 3.305 1.665 3.555 2.465 ;
      RECT 3.345 0.085 3.515 0.555 ;
      RECT 3.725 1.835 3.975 2.635 ;
      RECT 4.145 1.665 4.395 2.465 ;
      RECT 4.185 0.085 4.355 0.555 ;
      RECT 4.565 1.835 4.815 2.635 ;
      RECT 4.985 1.665 5.235 2.295 ;
      RECT 4.985 2.295 8.595 2.465 ;
      RECT 5.025 0.085 5.195 0.555 ;
      RECT 5.825 1.785 6.075 2.295 ;
      RECT 5.865 0.085 6.035 0.555 ;
      RECT 6.665 1.785 6.915 2.295 ;
      RECT 6.705 0.085 6.875 0.555 ;
      RECT 7.505 1.785 7.755 2.295 ;
      RECT 7.545 0.085 7.715 0.555 ;
      RECT 8.345 1.785 8.595 2.295 ;
      RECT 8.385 0.085 8.655 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.32 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 1.8 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.085 0.365 0.905 ;
      RECT 0.085 1.455 2.125 1.665 ;
      RECT 0.085 1.665 0.365 2.465 ;
      RECT 0.535 1.835 0.865 2.635 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.375 1.835 1.625 2.635 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.855 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 2.795 1.075 4.275 1.275 ;
      RECT 3.475 1.575 3.855 2.295 ;
      RECT 3.555 0.085 3.845 0.905 ;
      RECT 4.025 0.255 4.355 0.815 ;
      RECT 4.025 0.815 4.275 1.075 ;
      RECT 4.025 1.275 4.275 1.575 ;
      RECT 4.025 1.575 4.355 2.465 ;
      RECT 4.525 0.085 4.815 0.905 ;
      RECT 4.525 1.495 4.93 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4
MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915 0.275 13.255 0.825 ;
        RECT 12.915 1.495 13.255 2.45 ;
        RECT 13.07 0.825 13.255 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.5 0.255 11.83 2.465 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.345 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.765 0.825 1.675 ;
      LAYER mcon ;
        RECT 0.61 1.105 0.78 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
      LAYER mcon ;
        RECT 2.445 1.105 2.615 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.55 1.075 0.84 1.12 ;
        RECT 0.55 1.12 2.675 1.26 ;
        RECT 0.55 1.26 0.84 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.015 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.885 1.415 9.11 1.525 ;
        RECT 8.885 1.525 10.075 1.725 ;
      LAYER mcon ;
        RECT 8.885 1.445 9.055 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.115 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.825 1.415 9.115 1.46 ;
        RECT 8.825 1.6 9.115 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.59 ;
        RECT 2.905 1.59 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 13.53 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 13.34 0.085 ;
      RECT 0 2.635 13.34 2.805 ;
      RECT 0.085 0.085 0.48 0.595 ;
      RECT 0.085 1.845 1.105 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.515 2.195 0.765 2.635 ;
      RECT 0.875 0.28 1.655 0.56 ;
      RECT 0.935 2.025 1.105 2.255 ;
      RECT 0.935 2.255 2.045 2.465 ;
      RECT 1.295 1.87 1.695 2.075 ;
      RECT 1.38 0.56 1.655 0.59 ;
      RECT 1.38 0.59 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.67 0.62 ;
      RECT 1.44 0.62 1.67 0.63 ;
      RECT 1.445 0.63 1.67 0.635 ;
      RECT 1.46 0.635 1.67 0.645 ;
      RECT 1.475 0.645 1.67 0.655 ;
      RECT 1.475 0.655 1.695 0.665 ;
      RECT 1.495 0.665 1.695 0.705 ;
      RECT 1.505 0.705 1.695 1.87 ;
      RECT 1.825 0.085 2.005 0.545 ;
      RECT 1.865 0.715 2.515 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.515 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 2.69 0.085 3.03 0.555 ;
      RECT 2.69 2.14 3.03 2.635 ;
      RECT 3.255 1.775 3.995 1.955 ;
      RECT 3.255 1.955 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.595 2.275 3.925 2.635 ;
      RECT 3.63 0.085 3.94 0.545 ;
      RECT 3.735 0.885 3.995 1.775 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.11 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.61 1.59 4.915 1.615 ;
      RECT 4.61 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.66 1.275 ;
      RECT 5.03 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.435 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.61 0.085 6.095 0.465 ;
      RECT 5.61 0.635 6.535 0.805 ;
      RECT 5.61 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.765 2.105 ;
      RECT 5.945 2.275 6.275 2.635 ;
      RECT 6.25 0.975 7.66 1.225 ;
      RECT 6.275 0.255 6.535 0.635 ;
      RECT 6.55 2.105 6.765 2.45 ;
      RECT 6.735 0.085 7.63 0.805 ;
      RECT 7.005 2.125 7.96 2.635 ;
      RECT 7.19 1.495 8.005 1.955 ;
      RECT 7.3 1.275 7.66 1.325 ;
      RECT 7.835 0.695 9.04 0.895 ;
      RECT 7.835 0.895 8.005 1.495 ;
      RECT 8.13 2.125 8.935 2.46 ;
      RECT 8.365 1.075 8.595 1.905 ;
      RECT 8.41 0.275 9.825 0.445 ;
      RECT 8.765 1.895 10.465 2.065 ;
      RECT 8.765 2.065 8.935 2.125 ;
      RECT 8.81 0.895 9.04 1.245 ;
      RECT 9.195 2.235 9.525 2.635 ;
      RECT 9.29 0.855 9.465 1.185 ;
      RECT 9.29 1.185 10.895 1.355 ;
      RECT 9.655 0.445 9.825 0.845 ;
      RECT 9.655 0.845 10.545 1.015 ;
      RECT 9.695 2.065 9.91 2.45 ;
      RECT 10.135 2.235 10.465 2.635 ;
      RECT 10.22 0.085 10.39 0.545 ;
      RECT 10.245 1.525 10.465 1.895 ;
      RECT 10.56 0.255 10.895 0.54 ;
      RECT 10.635 1.355 10.895 2.465 ;
      RECT 10.715 0.54 10.895 1.185 ;
      RECT 11.12 0.085 11.33 0.885 ;
      RECT 11.12 1.485 11.33 2.635 ;
      RECT 12.06 0.255 12.27 0.995 ;
      RECT 12.06 0.995 12.9 1.325 ;
      RECT 12.06 1.325 12.27 2.465 ;
      RECT 12.54 0.085 12.745 0.825 ;
      RECT 12.575 1.575 12.745 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 1.785 7.675 1.955 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.735 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.655 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.445 1.755 7.735 1.8 ;
      RECT 7.445 1.94 7.735 1.985 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
  END
END sky130_fd_sc_hd__sdfsbp_1
MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.41 0.275 13.74 0.825 ;
        RECT 13.41 1.495 13.74 2.45 ;
        RECT 13.515 0.825 13.74 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.46 0.255 11.855 2.465 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
      LAYER mcon ;
        RECT 0.605 1.105 0.775 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 2.735 1.59 ;
      LAYER mcon ;
        RECT 2.445 1.105 2.615 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.435 9.115 1.525 ;
        RECT 8.88 1.525 9.935 1.725 ;
      LAYER mcon ;
        RECT 8.94 1.445 9.11 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.1 1.97 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 14.45 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.26 0.085 ;
      RECT 0 2.635 14.26 2.805 ;
      RECT 0.085 0.085 0.7 0.595 ;
      RECT 0.085 1.845 1.185 2.075 ;
      RECT 0.085 2.075 0.345 2.465 ;
      RECT 0.515 2.275 0.845 2.635 ;
      RECT 0.87 0.255 1.67 0.595 ;
      RECT 1.015 2.075 1.185 2.255 ;
      RECT 1.015 2.255 2.105 2.465 ;
      RECT 1.355 1.845 1.695 2.085 ;
      RECT 1.495 0.595 1.67 0.645 ;
      RECT 1.495 0.645 1.695 0.705 ;
      RECT 1.5 0.705 1.695 0.72 ;
      RECT 1.505 0.72 1.695 1.845 ;
      RECT 1.84 0.085 2.09 0.545 ;
      RECT 1.98 0.715 2.53 0.905 ;
      RECT 1.98 0.905 2.235 1.76 ;
      RECT 1.98 1.76 2.535 2.085 ;
      RECT 2.26 0.255 2.53 0.715 ;
      RECT 2.275 2.085 2.535 2.465 ;
      RECT 2.7 0.085 3.1 0.555 ;
      RECT 2.705 2.14 3.1 2.635 ;
      RECT 3.27 0.255 3.47 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.27 1.83 3.995 2 ;
      RECT 3.27 2 3.475 2.325 ;
      RECT 3.64 0.085 3.94 0.545 ;
      RECT 3.645 2.275 3.975 2.635 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.11 0.255 4.335 0.585 ;
      RECT 4.145 2.135 4.44 2.465 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.885 0.92 ;
      RECT 4.665 1.59 4.97 1.615 ;
      RECT 4.665 1.615 4.89 2.465 ;
      RECT 4.715 0.92 4.885 1.445 ;
      RECT 4.715 1.445 4.97 1.59 ;
      RECT 5.055 0.255 5.45 1.225 ;
      RECT 5.055 1.225 7.705 1.275 ;
      RECT 5.06 2.135 5.805 2.465 ;
      RECT 5.14 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.465 1.955 ;
      RECT 5.62 0.635 6.55 0.805 ;
      RECT 5.62 0.805 6.015 1.015 ;
      RECT 5.635 1.395 5.805 2.135 ;
      RECT 5.665 0.085 6.165 0.465 ;
      RECT 5.975 1.575 6.145 1.935 ;
      RECT 5.975 1.935 6.82 2.105 ;
      RECT 6 2.275 6.33 2.635 ;
      RECT 6.305 0.975 7.705 1.225 ;
      RECT 6.335 0.255 6.55 0.635 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 6.72 0.085 7.705 0.805 ;
      RECT 7.06 2.125 8.015 2.635 ;
      RECT 7.355 1.275 7.705 1.325 ;
      RECT 7.385 1.705 8.055 1.955 ;
      RECT 7.885 0.695 9.085 0.895 ;
      RECT 7.885 0.895 8.055 1.705 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.42 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.855 0.515 ;
      RECT 8.82 1.895 10.43 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 8.83 0.895 9.085 1.265 ;
      RECT 9.16 2.235 9.49 2.635 ;
      RECT 9.285 0.855 9.515 1.185 ;
      RECT 9.285 1.185 10.91 1.355 ;
      RECT 9.66 2.065 9.93 2.45 ;
      RECT 9.685 0.515 9.855 0.845 ;
      RECT 9.685 0.845 10.56 1.015 ;
      RECT 10.035 0.085 10.285 0.545 ;
      RECT 10.1 2.235 10.43 2.635 ;
      RECT 10.105 1.525 10.43 1.895 ;
      RECT 10.465 0.255 10.91 0.585 ;
      RECT 10.6 1.355 10.845 2.465 ;
      RECT 10.73 0.585 10.91 1.185 ;
      RECT 11.08 1.485 11.29 2.635 ;
      RECT 11.12 0.085 11.29 0.885 ;
      RECT 12.025 0.085 12.315 0.885 ;
      RECT 12.025 1.485 12.315 2.635 ;
      RECT 12.53 0.255 12.715 0.995 ;
      RECT 12.53 0.995 13.345 1.325 ;
      RECT 12.53 1.325 12.715 2.465 ;
      RECT 12.885 0.085 13.24 0.825 ;
      RECT 12.885 1.635 13.24 2.635 ;
      RECT 13.91 0.085 14.175 0.885 ;
      RECT 13.91 1.485 14.175 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.26 1.785 5.43 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.48 1.105 8.65 1.275 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 5.03 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.2 1.755 5.49 1.8 ;
      RECT 5.2 1.94 5.49 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfsbp_2
MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.265 1.275 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 0.255 4.545 0.26 ;
        RECT 4.295 0.26 4.625 0.735 ;
        RECT 4.295 0.735 10.955 0.905 ;
        RECT 4.295 1.445 10.955 1.615 ;
        RECT 4.295 1.615 4.625 2.465 ;
        RECT 5.135 0.26 5.465 0.735 ;
        RECT 5.135 1.615 5.465 2.465 ;
        RECT 5.215 0.255 5.385 0.26 ;
        RECT 5.975 0.26 6.305 0.735 ;
        RECT 5.975 1.615 6.305 2.465 ;
        RECT 6.055 0.255 6.225 0.26 ;
        RECT 6.815 0.26 7.145 0.735 ;
        RECT 6.815 1.615 7.145 2.465 ;
        RECT 7.655 0.26 7.985 0.735 ;
        RECT 7.655 1.615 7.985 2.465 ;
        RECT 8.495 0.26 8.825 0.735 ;
        RECT 8.495 1.615 8.825 2.465 ;
        RECT 9.335 0.26 9.665 0.735 ;
        RECT 9.335 1.615 9.665 2.465 ;
        RECT 10.175 0.26 10.505 0.735 ;
        RECT 10.175 1.615 10.505 2.465 ;
        RECT 10.68 0.905 10.955 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.095 0.26 0.425 0.735 ;
      RECT 0.095 0.735 1.605 0.905 ;
      RECT 0.095 1.445 1.605 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.595 0.085 0.765 0.565 ;
      RECT 0.595 1.785 0.765 2.635 ;
      RECT 0.935 0.26 1.265 0.735 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.435 0.085 1.605 0.565 ;
      RECT 1.435 0.905 1.605 1.075 ;
      RECT 1.435 1.075 3.745 1.275 ;
      RECT 1.435 1.275 1.605 1.445 ;
      RECT 1.435 1.785 1.605 2.635 ;
      RECT 1.775 0.26 2.105 0.735 ;
      RECT 1.775 0.735 4.125 0.905 ;
      RECT 1.775 1.445 4.125 1.615 ;
      RECT 1.775 1.615 2.105 2.465 ;
      RECT 2.275 0.085 2.445 0.565 ;
      RECT 2.275 1.835 2.445 2.635 ;
      RECT 2.615 0.26 2.945 0.735 ;
      RECT 2.615 1.615 2.945 2.465 ;
      RECT 3.115 0.085 3.285 0.565 ;
      RECT 3.115 1.835 3.285 2.635 ;
      RECT 3.455 0.26 3.785 0.735 ;
      RECT 3.455 1.615 3.785 2.465 ;
      RECT 3.95 0.905 4.125 1.075 ;
      RECT 3.95 1.075 10.51 1.275 ;
      RECT 3.95 1.275 4.125 1.445 ;
      RECT 3.955 0.085 4.125 0.565 ;
      RECT 3.955 1.835 4.125 2.635 ;
      RECT 4.795 0.085 4.965 0.565 ;
      RECT 4.795 1.835 4.965 2.635 ;
      RECT 5.635 0.085 5.805 0.565 ;
      RECT 5.635 1.835 5.805 2.635 ;
      RECT 6.475 0.085 6.645 0.565 ;
      RECT 6.475 1.835 6.645 2.635 ;
      RECT 7.315 0.085 7.485 0.565 ;
      RECT 7.315 1.835 7.485 2.635 ;
      RECT 8.155 0.085 8.325 0.565 ;
      RECT 8.155 1.835 8.325 2.635 ;
      RECT 8.995 0.085 9.165 0.565 ;
      RECT 8.995 1.835 9.165 2.635 ;
      RECT 9.835 0.085 10.005 0.565 ;
      RECT 9.835 1.835 10.005 2.635 ;
      RECT 10.675 0.085 10.845 0.565 ;
      RECT 10.675 1.835 10.845 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
  END
END sky130_fd_sc_hd__bufinv_16
MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.505 1.275 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.26 3.045 0.735 ;
        RECT 2.715 0.735 6.355 0.905 ;
        RECT 2.715 1.445 6.355 1.615 ;
        RECT 2.715 1.615 3.045 2.465 ;
        RECT 3.555 0.26 3.885 0.735 ;
        RECT 3.555 1.615 3.885 2.465 ;
        RECT 4.395 0.26 4.725 0.735 ;
        RECT 4.395 1.615 4.725 2.465 ;
        RECT 5.235 0.26 5.565 0.735 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 5.97 0.905 6.355 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.175 0.085 0.345 0.905 ;
      RECT 0.175 1.445 0.345 2.635 ;
      RECT 0.515 0.26 0.845 0.905 ;
      RECT 0.515 1.545 0.845 2.465 ;
      RECT 0.675 0.905 0.845 1.075 ;
      RECT 0.675 1.075 2.205 1.275 ;
      RECT 0.675 1.275 0.845 1.545 ;
      RECT 1.035 0.26 1.365 0.735 ;
      RECT 1.035 0.735 2.545 0.905 ;
      RECT 1.035 1.445 2.545 1.615 ;
      RECT 1.035 1.615 1.365 2.465 ;
      RECT 1.535 0.085 1.705 0.565 ;
      RECT 1.535 1.785 1.705 2.635 ;
      RECT 1.875 0.26 2.205 0.735 ;
      RECT 1.875 1.615 2.205 2.465 ;
      RECT 2.375 0.085 2.545 0.565 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 5.76 1.275 ;
      RECT 2.375 1.275 2.545 1.445 ;
      RECT 2.375 1.785 2.545 2.635 ;
      RECT 3.215 0.085 3.385 0.565 ;
      RECT 3.215 1.835 3.385 2.635 ;
      RECT 4.055 0.085 4.225 0.565 ;
      RECT 4.055 1.835 4.225 2.635 ;
      RECT 4.895 0.085 5.065 0.565 ;
      RECT 4.895 1.835 5.065 2.635 ;
      RECT 5.735 0.085 5.905 0.565 ;
      RECT 5.735 1.835 5.905 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__bufinv_8
MACRO sky130_fd_sc_hd__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.415 2.175 0.7 ;
        RECT 1.965 0.7 2.355 0.87 ;
        RECT 2.185 0.87 2.355 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.4 1.7 0.695 ;
        RECT 1.53 0.695 1.795 0.865 ;
        RECT 1.625 0.865 1.795 1.075 ;
        RECT 1.625 1.075 1.955 1.245 ;
        RECT 1.625 1.245 1.795 1.26 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.76 1.27 0.995 ;
        RECT 1.065 0.995 1.395 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.755 3.09 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.715 0.765 0.885 ;
        RECT 0.09 0.885 0.345 1.835 ;
        RECT 0.09 1.835 0.765 2.005 ;
        RECT 0.595 0.255 0.765 0.715 ;
        RECT 0.595 2.005 0.765 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.09 0.085 0.345 0.545 ;
      RECT 0.135 2.175 0.385 2.635 ;
      RECT 0.555 1.075 0.885 1.245 ;
      RECT 0.555 1.245 0.725 1.495 ;
      RECT 0.555 1.495 3.045 1.665 ;
      RECT 0.935 1.835 1.185 2.635 ;
      RECT 0.955 0.085 1.285 0.465 ;
      RECT 1.015 0.465 1.185 0.545 ;
      RECT 1.355 1.835 2.645 2.005 ;
      RECT 1.355 2.005 1.605 2.425 ;
      RECT 1.815 2.175 2.145 2.635 ;
      RECT 2.335 2.005 2.585 2.425 ;
      RECT 2.375 0.335 2.705 0.505 ;
      RECT 2.46 0.255 2.705 0.335 ;
      RECT 2.535 0.505 2.705 1.495 ;
      RECT 2.875 0.085 3.135 0.565 ;
      RECT 2.875 1.665 3.045 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a31o_2
MACRO sky130_fd_sc_hd__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.16 1.655 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.7 1.655 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.995 1.24 1.325 ;
        RECT 1.025 1.325 1.24 1.655 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 0.995 2.62 1.655 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.3 0.425 0.81 ;
        RECT 0.095 0.81 0.285 1.575 ;
        RECT 0.095 1.575 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.455 0.995 0.765 1.325 ;
      RECT 0.595 0.085 0.925 0.485 ;
      RECT 0.595 0.655 2.96 0.825 ;
      RECT 0.595 0.825 0.765 0.995 ;
      RECT 0.595 1.495 0.845 2.635 ;
      RECT 1.035 1.825 2.325 1.995 ;
      RECT 1.035 1.995 1.285 2.415 ;
      RECT 1.515 2.165 1.845 2.635 ;
      RECT 1.975 0.315 2.305 0.655 ;
      RECT 2.075 1.995 2.325 2.415 ;
      RECT 2.475 0.085 2.805 0.485 ;
      RECT 2.505 1.825 2.96 1.995 ;
      RECT 2.505 1.995 2.835 2.425 ;
      RECT 2.79 0.825 2.96 1.825 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a31o_1
MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 1.705 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.075 1.055 1.245 ;
        RECT 0.805 0.735 2.17 0.905 ;
        RECT 0.805 0.905 0.975 1.075 ;
        RECT 1.985 0.905 2.17 1.075 ;
        RECT 1.985 1.075 2.315 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.525 1.445 ;
        RECT 0.15 1.445 2.855 1.615 ;
        RECT 2.525 1.075 2.855 1.445 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.575 1.075 4.03 1.285 ;
        RECT 3.815 0.745 4.03 1.075 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.655 6.295 0.825 ;
        RECT 4.535 1.785 6.295 1.955 ;
        RECT 4.595 1.955 4.765 2.465 ;
        RECT 5.435 1.955 5.605 2.465 ;
        RECT 6.125 0.825 6.295 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.175 0.085 0.345 0.905 ;
      RECT 0.175 1.785 2.985 1.955 ;
      RECT 0.175 1.955 0.345 2.465 ;
      RECT 0.515 2.125 0.845 2.635 ;
      RECT 1.015 1.955 1.185 2.465 ;
      RECT 1.355 0.395 2.52 0.565 ;
      RECT 1.355 2.125 1.685 2.635 ;
      RECT 1.855 1.955 2.025 2.465 ;
      RECT 2.195 2.125 2.525 2.635 ;
      RECT 2.35 0.565 2.52 0.7 ;
      RECT 2.35 0.7 3.485 0.805 ;
      RECT 2.35 0.805 3.345 0.87 ;
      RECT 2.7 0.085 2.985 0.53 ;
      RECT 2.815 1.955 2.985 2.295 ;
      RECT 2.815 2.295 3.825 2.465 ;
      RECT 3.155 0.295 3.485 0.7 ;
      RECT 3.155 0.87 3.345 1.455 ;
      RECT 3.155 1.455 4.395 1.625 ;
      RECT 3.155 1.625 3.485 2.115 ;
      RECT 3.655 1.795 3.825 2.295 ;
      RECT 3.735 0.085 4.265 0.565 ;
      RECT 4.095 2.125 4.425 2.635 ;
      RECT 4.225 0.995 5.935 1.325 ;
      RECT 4.225 1.325 4.395 1.455 ;
      RECT 4.935 0.085 5.265 0.485 ;
      RECT 4.935 2.125 5.265 2.635 ;
      RECT 5.775 0.085 6.105 0.485 ;
      RECT 5.775 2.125 6.105 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
  END
END sky130_fd_sc_hd__a31o_4
MACRO sky130_fd_sc_hd__lpflow_inputiso0p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.645 2.175 1.955 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.58 2.655 2.365 ;
        RECT 2.415 0.255 2.655 0.775 ;
        RECT 2.48 0.775 2.655 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 0.085 0.425 0.59 ;
      RECT 0.175 1.785 0.85 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.515 2.185 0.845 2.635 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.615 0.655 0.835 0.805 ;
      RECT 0.615 0.805 1.15 1.135 ;
      RECT 0.615 1.135 0.85 1.785 ;
      RECT 1.02 1.305 2.305 1.325 ;
      RECT 1.02 1.325 1.88 1.475 ;
      RECT 1.02 1.475 1.305 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.49 0.61 ;
      RECT 1.32 0.61 1.49 0.945 ;
      RECT 1.32 0.945 2.305 1.305 ;
      RECT 1.485 2.165 2.17 2.635 ;
      RECT 1.85 0.085 2.245 0.58 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0p_1
MACRO sky130_fd_sc_hd__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.89 1.495 7.3 1.575 ;
        RECT 6.89 1.575 7.22 2.42 ;
        RECT 6.9 0.305 7.23 0.74 ;
        RECT 6.9 0.74 7.3 0.825 ;
        RECT 7.055 0.825 7.3 0.865 ;
        RECT 7.065 1.445 7.3 1.495 ;
        RECT 7.11 0.865 7.3 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.315 1.48 8.65 2.465 ;
        RECT 8.395 0.255 8.65 0.91 ;
        RECT 8.415 0.91 8.65 1.48 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.44 2.175 1.705 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.4 0.085 3.77 0.585 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.61 1.835 3.78 2.635 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.02 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.38 1.905 ;
      RECT 5.49 2.135 5.805 2.635 ;
      RECT 5.585 0.085 5.795 0.615 ;
      RECT 6.04 1.905 6.38 2.465 ;
      RECT 6.06 0.3 6.39 0.825 ;
      RECT 6.19 0.825 6.39 0.995 ;
      RECT 6.19 0.995 6.94 1.325 ;
      RECT 6.19 1.325 6.38 1.53 ;
      RECT 6.55 1.625 6.72 2.635 ;
      RECT 6.56 0.085 6.73 0.695 ;
      RECT 7.41 1.715 7.74 2.445 ;
      RECT 7.42 0.345 7.67 0.615 ;
      RECT 7.47 0.615 7.67 0.995 ;
      RECT 7.47 0.995 8.245 1.325 ;
      RECT 7.47 1.325 7.74 1.715 ;
      RECT 7.905 0.085 8.225 0.545 ;
      RECT 7.93 1.495 8.145 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxbp_1
MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.89 1.495 7.3 1.575 ;
        RECT 6.89 1.575 7.22 2.42 ;
        RECT 6.9 0.305 7.23 0.74 ;
        RECT 6.9 0.74 7.3 0.825 ;
        RECT 7.055 0.825 7.3 0.865 ;
        RECT 7.065 1.445 7.3 1.495 ;
        RECT 7.11 0.865 7.3 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.81 1.495 9.145 2.465 ;
        RECT 8.89 0.265 9.145 0.885 ;
        RECT 8.93 0.885 9.145 1.495 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.44 2.175 1.705 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.4 0.085 3.77 0.585 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.61 1.835 3.78 2.635 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.02 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.38 1.905 ;
      RECT 5.49 2.135 5.805 2.635 ;
      RECT 5.585 0.085 5.795 0.615 ;
      RECT 6.04 1.905 6.38 2.465 ;
      RECT 6.06 0.3 6.39 0.825 ;
      RECT 6.19 0.825 6.39 0.995 ;
      RECT 6.19 0.995 6.94 1.325 ;
      RECT 6.19 1.325 6.38 1.53 ;
      RECT 6.55 1.625 6.72 2.635 ;
      RECT 6.56 0.085 6.73 0.695 ;
      RECT 7.39 1.72 7.565 2.635 ;
      RECT 7.4 0.085 7.57 0.6 ;
      RECT 7.905 0.345 8.165 0.615 ;
      RECT 7.905 1.715 8.235 2.445 ;
      RECT 7.965 0.615 8.165 0.995 ;
      RECT 7.965 0.995 8.76 1.325 ;
      RECT 7.965 1.325 8.235 1.715 ;
      RECT 8.39 0.085 8.72 0.825 ;
      RECT 8.425 1.495 8.64 2.635 ;
      RECT 9.315 0.085 9.565 0.905 ;
      RECT 9.315 1.495 9.565 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxbp_2
MACRO sky130_fd_sc_hd__dlxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 0.955 1.685 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 0.255 5.49 0.82 ;
        RECT 5.14 1.67 5.49 2.455 ;
        RECT 5.32 0.82 5.49 1.67 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555 0.255 6.815 0.825 ;
        RECT 6.555 1.445 6.815 2.465 ;
        RECT 6.6 0.825 6.815 1.445 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.795 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.135 0.785 ;
      RECT 1.855 0.785 2.135 0.875 ;
      RECT 1.855 0.875 2.335 1.235 ;
      RECT 1.855 1.235 2.115 1.495 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.965 1.835 2.245 2.635 ;
      RECT 2.465 1.355 2.795 1.685 ;
      RECT 2.58 0.705 3.135 1.065 ;
      RECT 2.75 2.255 3.61 2.425 ;
      RECT 2.8 0.365 3.475 0.535 ;
      RECT 2.965 1.065 3.135 1.575 ;
      RECT 2.965 1.575 3.29 1.91 ;
      RECT 2.965 1.91 3.195 1.995 ;
      RECT 3.305 0.535 3.475 0.995 ;
      RECT 3.305 0.995 4.175 1.165 ;
      RECT 3.425 2.035 3.65 2.065 ;
      RECT 3.425 2.065 3.63 2.09 ;
      RECT 3.425 2.09 3.61 2.255 ;
      RECT 3.43 2.02 3.65 2.035 ;
      RECT 3.435 2.01 3.65 2.02 ;
      RECT 3.44 1.995 3.65 2.01 ;
      RECT 3.46 1.165 4.175 1.325 ;
      RECT 3.46 1.325 3.65 1.995 ;
      RECT 3.7 0.085 4.045 0.53 ;
      RECT 3.78 2.175 3.98 2.635 ;
      RECT 3.82 1.535 4.515 1.865 ;
      RECT 4.285 0.415 4.55 0.745 ;
      RECT 4.285 1.865 4.515 2.435 ;
      RECT 4.345 0.745 4.55 0.995 ;
      RECT 4.345 0.995 5.15 1.325 ;
      RECT 4.345 1.325 4.515 1.535 ;
      RECT 4.685 1.57 4.97 2.635 ;
      RECT 4.72 0.085 4.97 0.715 ;
      RECT 5.66 0.255 5.91 0.995 ;
      RECT 5.66 0.995 6.43 1.325 ;
      RECT 5.66 1.325 5.91 2.465 ;
      RECT 6.09 0.085 6.385 0.545 ;
      RECT 6.09 1.835 6.385 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.555 1.445 2.725 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.965 1.785 3.135 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.785 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.195 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.495 1.415 2.785 1.46 ;
      RECT 2.495 1.6 2.785 1.645 ;
      RECT 2.905 1.755 3.195 1.8 ;
      RECT 2.905 1.94 3.195 1.985 ;
  END
END sky130_fd_sc_hd__dlxbp_1
MACRO sky130_fd_sc_hd__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 1.755000 0.375000 1.985000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  1.785000 0.315000 1.955000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd2_1
MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.86 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.415 0.255 14.665 0.825 ;
        RECT 14.415 1.445 14.665 2.465 ;
        RECT 14.46 0.825 14.665 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.58 0.255 12.83 0.715 ;
        RECT 12.58 1.63 12.83 2.465 ;
        RECT 12.66 0.715 12.83 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.59 1.095 12.07 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.345 2.145 0.765 ;
        RECT 1.935 0.765 2.335 1.095 ;
        RECT 1.935 1.095 2.155 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 5.885 0.965 6.215 1.065 ;
      LAYER mcon ;
        RECT 6.125 0.765 6.295 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
      LAYER mcon ;
        RECT 9.805 0.765 9.975 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 15.18 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 15.37 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 15.18 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 15.18 0.085 ;
      RECT 0 2.635 15.18 2.805 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.835 0.805 ;
      RECT 0.17 1.795 0.835 1.965 ;
      RECT 0.17 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 1.43 0.085 1.705 0.635 ;
      RECT 1.43 1.885 1.785 2.635 ;
      RECT 2.215 1.875 2.575 2.385 ;
      RECT 2.315 0.265 2.73 0.595 ;
      RECT 2.405 1.25 3.075 1.405 ;
      RECT 2.405 1.405 2.575 1.875 ;
      RECT 2.435 1.235 3.075 1.25 ;
      RECT 2.56 0.595 2.73 1.075 ;
      RECT 2.56 1.075 3.075 1.235 ;
      RECT 2.745 1.575 3.645 1.745 ;
      RECT 2.745 1.745 3.065 1.905 ;
      RECT 2.895 1.905 3.065 2.465 ;
      RECT 2.955 0.305 3.125 0.625 ;
      RECT 2.955 0.625 3.645 0.765 ;
      RECT 2.955 0.765 3.77 0.795 ;
      RECT 3.295 2.215 3.64 2.635 ;
      RECT 3.37 0.085 3.7 0.445 ;
      RECT 3.475 0.795 3.77 1.095 ;
      RECT 3.475 1.095 3.645 1.575 ;
      RECT 4.23 0.305 4.455 2.465 ;
      RECT 4.625 0.705 4.845 1.575 ;
      RECT 4.625 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 4.7 0.265 5.715 0.465 ;
      RECT 5.025 0.645 5.375 1.015 ;
      RECT 5.295 1.195 5.715 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.545 0.465 5.715 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 5.705 2.205 6.085 2.635 ;
      RECT 5.885 0.085 6.055 0.525 ;
      RECT 6.225 0.255 7.375 0.425 ;
      RECT 6.225 0.425 6.555 0.505 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.705 0.595 7.035 0.765 ;
      RECT 6.815 0.765 7.035 0.895 ;
      RECT 6.815 0.895 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.175 1.915 7.505 2.635 ;
      RECT 7.205 0.425 7.375 0.715 ;
      RECT 7.645 0.085 7.975 0.465 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.41 2.085 ;
      RECT 9.56 0.085 9.82 0.525 ;
      RECT 9.62 2.255 10 2.635 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.41 0.545 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.58 0.595 10.91 0.78 ;
      RECT 10.73 0.78 10.91 1.915 ;
      RECT 10.94 2.255 12.41 2.635 ;
      RECT 11.08 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.845 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.925 1.745 ;
      RECT 11.62 0.265 11.845 0.755 ;
      RECT 12.08 0.085 12.41 0.805 ;
      RECT 12.24 0.995 12.48 1.325 ;
      RECT 12.24 1.325 12.41 1.915 ;
      RECT 13 0.085 13.235 0.885 ;
      RECT 13 1.495 13.235 2.635 ;
      RECT 13.455 0.255 13.77 0.995 ;
      RECT 13.455 0.995 14.29 1.325 ;
      RECT 13.455 1.325 13.77 2.415 ;
      RECT 13.95 0.085 14.245 0.545 ;
      RECT 13.95 1.765 14.245 2.635 ;
      RECT 14.835 0.085 15.075 0.885 ;
      RECT 14.835 1.495 15.075 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 0.765 0.775 0.935 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 1.445 11.355 1.615 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 14.405 2.635 14.575 2.805 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.865 2.635 15.035 2.805 ;
    LAYER met1 ;
      RECT 0.545 0.735 0.835 0.78 ;
      RECT 0.545 0.78 5.435 0.92 ;
      RECT 0.545 0.92 0.835 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 8.655 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.515 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.22 0.965 5.435 1.12 ;
      RECT 5.22 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbn_2
MACRO sky130_fd_sc_hd__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.405 4.105 1.575 ;
        RECT 3.775 1.575 4.06 1.675 ;
        RECT 3.825 1.675 4.06 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915 0.255 14.175 0.785 ;
        RECT 13.915 1.47 14.175 2.465 ;
        RECT 13.965 0.785 14.175 1.47 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.5 0.255 12.785 0.715 ;
        RECT 12.5 1.63 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.99 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.345 2.155 0.815 ;
        RECT 1.935 0.815 2.315 1.15 ;
        RECT 1.935 1.15 2.155 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.87 0.735 6.295 0.965 ;
        RECT 5.87 0.965 6.215 1.065 ;
      LAYER mcon ;
        RECT 6.125 0.765 6.295 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
      LAYER mcon ;
        RECT 9.805 0.765 9.975 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 14.45 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.26 0.085 ;
      RECT 0 2.635 14.26 2.805 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.095 1.795 0.835 1.965 ;
      RECT 0.095 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 1.43 0.085 1.705 0.635 ;
      RECT 1.43 1.885 1.785 2.635 ;
      RECT 2.215 1.875 2.575 2.385 ;
      RECT 2.325 0.265 2.655 0.595 ;
      RECT 2.405 1.295 3.075 1.405 ;
      RECT 2.405 1.405 2.67 1.43 ;
      RECT 2.405 1.43 2.63 1.465 ;
      RECT 2.405 1.465 2.605 1.505 ;
      RECT 2.405 1.505 2.575 1.875 ;
      RECT 2.46 1.255 3.075 1.295 ;
      RECT 2.485 0.595 2.655 1.075 ;
      RECT 2.485 1.075 3.075 1.255 ;
      RECT 2.76 1.575 3.605 1.745 ;
      RECT 2.76 1.745 3.14 1.905 ;
      RECT 2.87 0.305 3.04 0.625 ;
      RECT 2.87 0.625 3.645 0.765 ;
      RECT 2.87 0.765 3.77 0.795 ;
      RECT 2.97 1.905 3.14 2.465 ;
      RECT 3.225 0.085 3.555 0.445 ;
      RECT 3.31 2.215 3.64 2.635 ;
      RECT 3.43 0.795 3.77 1.095 ;
      RECT 3.43 1.095 3.605 1.575 ;
      RECT 3.95 0.425 4.33 0.595 ;
      RECT 3.95 0.595 4.12 1.065 ;
      RECT 3.95 1.065 4.4 1.105 ;
      RECT 3.95 1.105 4.41 1.175 ;
      RECT 3.95 1.175 4.445 1.235 ;
      RECT 4.16 0.265 4.33 0.425 ;
      RECT 4.225 1.235 4.445 1.275 ;
      RECT 4.23 2.135 4.445 2.465 ;
      RECT 4.245 1.275 4.445 1.305 ;
      RECT 4.275 1.305 4.445 2.135 ;
      RECT 4.555 0.265 5.655 0.465 ;
      RECT 4.57 0.705 4.79 1.035 ;
      RECT 4.615 1.035 4.79 1.575 ;
      RECT 4.615 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 5 0.735 5.33 1.015 ;
      RECT 5.295 1.195 5.67 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.485 0.465 5.655 0.585 ;
      RECT 5.485 0.585 5.67 0.655 ;
      RECT 5.5 0.655 5.67 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 5.705 2.205 6.085 2.635 ;
      RECT 5.835 0.085 6.005 0.525 ;
      RECT 6.26 0.255 7.35 0.425 ;
      RECT 6.26 0.425 6.59 0.465 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.68 0.61 7.01 0.78 ;
      RECT 6.81 0.78 7.01 0.895 ;
      RECT 6.81 0.895 8.125 1.06 ;
      RECT 6.815 1.06 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.175 1.915 7.505 2.635 ;
      RECT 7.18 0.425 7.35 0.715 ;
      RECT 7.62 0.085 7.975 0.465 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.33 2.085 ;
      RECT 9.56 0.085 9.82 0.525 ;
      RECT 9.62 2.255 10 2.635 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.41 0.545 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.575 0.595 10.905 0.78 ;
      RECT 10.73 0.78 10.905 1.915 ;
      RECT 10.94 2.255 12.33 2.635 ;
      RECT 11.075 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.775 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.855 1.745 ;
      RECT 11.565 0.265 11.775 0.755 ;
      RECT 12 0.085 12.33 0.805 ;
      RECT 12.16 0.995 12.425 1.325 ;
      RECT 12.16 1.325 12.33 1.915 ;
      RECT 12.96 0.255 13.275 0.995 ;
      RECT 12.96 0.995 13.795 1.325 ;
      RECT 12.96 1.325 13.275 2.415 ;
      RECT 13.455 0.085 13.745 0.545 ;
      RECT 13.455 1.765 13.74 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 0.765 0.775 0.935 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.23 1.105 4.4 1.275 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.155 0.765 5.325 0.935 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 1.445 11.355 1.615 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
    LAYER met1 ;
      RECT 0.545 0.735 0.835 0.78 ;
      RECT 0.545 0.78 5.385 0.92 ;
      RECT 0.545 0.92 0.835 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 8.655 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.46 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.17 1.075 4.46 1.12 ;
      RECT 4.17 1.26 4.46 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.095 0.735 5.385 0.78 ;
      RECT 5.095 0.92 5.385 0.965 ;
      RECT 5.17 0.965 5.385 1.12 ;
      RECT 5.17 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbn_1
MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.955 1.195 1.445 ;
        RECT 0.855 1.445 1.24 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.5 0.255 6.83 0.445 ;
        RECT 6.58 0.445 6.83 0.715 ;
        RECT 6.58 0.715 7.22 0.885 ;
        RECT 6.58 1.485 7.22 1.655 ;
        RECT 6.58 1.655 6.83 2.465 ;
        RECT 7.05 0.885 7.22 1.055 ;
        RECT 7.05 1.055 8.195 1.315 ;
        RECT 7.05 1.315 7.22 1.485 ;
        RECT 7.42 0.255 7.72 1.055 ;
        RECT 7.42 1.315 7.72 2.465 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.345 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.725 0.995 4.945 1.325 ;
      LAYER mcon ;
        RECT 4.77 1.105 4.94 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.685 0.995 6.065 1.325 ;
      LAYER mcon ;
        RECT 5.71 1.105 5.88 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.71 1.075 5 1.12 ;
        RECT 4.71 1.12 5.94 1.26 ;
        RECT 4.71 1.26 5 1.305 ;
        RECT 5.65 1.075 5.94 1.12 ;
        RECT 5.65 1.26 5.94 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.195 0.785 ;
      RECT 0.085 1.835 0.345 2.635 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.515 0.785 0.685 2.125 ;
      RECT 0.515 2.125 1.26 2.465 ;
      RECT 1.015 0.255 1.195 0.615 ;
      RECT 1.365 0.255 2.5 0.535 ;
      RECT 1.365 0.705 1.705 1.205 ;
      RECT 1.365 1.205 1.865 1.325 ;
      RECT 1.41 1.325 1.865 1.955 ;
      RECT 1.43 2.125 2.205 2.465 ;
      RECT 1.875 0.705 2.16 1.035 ;
      RECT 2.035 1.205 3.015 1.375 ;
      RECT 2.035 1.375 2.205 2.125 ;
      RECT 2.33 0.535 2.5 0.995 ;
      RECT 2.33 0.995 3.015 1.205 ;
      RECT 2.375 1.575 2.545 1.635 ;
      RECT 2.375 1.635 3.405 1.905 ;
      RECT 2.375 2.075 3.015 2.635 ;
      RECT 2.67 0.085 3.015 0.825 ;
      RECT 3.185 0.255 3.405 1.635 ;
      RECT 3.185 1.905 3.405 1.915 ;
      RECT 3.185 1.915 5.515 2.085 ;
      RECT 3.185 2.085 3.405 2.465 ;
      RECT 3.595 0.255 3.925 0.765 ;
      RECT 3.595 0.765 4.02 0.935 ;
      RECT 3.595 0.935 3.765 1.575 ;
      RECT 3.595 1.575 4.005 1.745 ;
      RECT 3.595 2.255 5.515 2.635 ;
      RECT 3.935 1.105 4.48 1.275 ;
      RECT 4.095 0.085 4.425 0.445 ;
      RECT 4.175 1.275 4.48 1.495 ;
      RECT 4.175 1.495 4.975 1.745 ;
      RECT 4.19 0.615 4.845 0.785 ;
      RECT 4.19 0.785 4.48 1.105 ;
      RECT 4.595 0.255 4.845 0.615 ;
      RECT 5.015 0.255 5.435 0.615 ;
      RECT 5.015 0.615 6.41 0.785 ;
      RECT 5.165 0.995 5.515 1.915 ;
      RECT 5.605 0.085 6.33 0.445 ;
      RECT 5.685 1.495 6.41 2.085 ;
      RECT 5.685 2.085 5.855 2.465 ;
      RECT 6.055 2.255 6.385 2.635 ;
      RECT 6.24 0.785 6.41 1.055 ;
      RECT 6.24 1.055 6.88 1.315 ;
      RECT 6.24 1.315 6.41 1.495 ;
      RECT 7 0.085 7.25 0.545 ;
      RECT 7 1.825 7.25 2.635 ;
      RECT 7.89 0.085 8.195 0.885 ;
      RECT 7.89 1.485 8.195 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 1.445 1.7 1.615 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.99 0.765 2.16 0.935 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.85 0.765 4.02 0.935 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.31 1.445 4.48 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 1.47 1.415 1.76 1.46 ;
      RECT 1.47 1.46 4.54 1.6 ;
      RECT 1.47 1.6 1.76 1.645 ;
      RECT 1.93 0.735 2.22 0.78 ;
      RECT 1.93 0.78 4.08 0.92 ;
      RECT 1.93 0.92 2.22 0.965 ;
      RECT 3.79 0.735 4.08 0.78 ;
      RECT 3.79 0.92 4.08 0.965 ;
      RECT 4.25 1.415 4.54 1.46 ;
      RECT 4.25 1.6 4.54 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_4
MACRO sky130_fd_sc_hd__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.955 1.195 1.445 ;
        RECT 0.855 1.445 1.24 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.57 0.255 6.84 0.825 ;
        RECT 6.57 1.495 6.84 2.465 ;
        RECT 6.67 0.825 6.84 1.055 ;
        RECT 6.67 1.055 7.275 1.315 ;
        RECT 6.67 1.315 6.84 1.495 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.34 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.705 0.955 6.05 1.265 ;
        RECT 4.705 1.265 4.925 1.325 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.195 0.785 ;
      RECT 0.085 1.835 0.345 2.635 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.515 0.785 0.685 2.125 ;
      RECT 0.515 2.125 1.26 2.465 ;
      RECT 1.015 0.255 1.195 0.615 ;
      RECT 1.365 0.255 2.5 0.535 ;
      RECT 1.365 0.705 1.705 1.205 ;
      RECT 1.365 1.205 1.865 1.325 ;
      RECT 1.41 1.325 1.865 1.955 ;
      RECT 1.43 2.125 2.205 2.465 ;
      RECT 1.875 0.705 2.16 1.035 ;
      RECT 2.035 1.205 3.015 1.375 ;
      RECT 2.035 1.375 2.205 2.125 ;
      RECT 2.33 0.535 2.5 0.995 ;
      RECT 2.33 0.995 3.015 1.205 ;
      RECT 2.375 1.575 2.545 1.635 ;
      RECT 2.375 1.635 3.405 1.905 ;
      RECT 2.375 2.075 3.015 2.635 ;
      RECT 2.67 0.085 3.015 0.825 ;
      RECT 3.185 0.255 3.405 1.635 ;
      RECT 3.185 1.905 3.405 1.915 ;
      RECT 3.185 1.915 5.49 2.085 ;
      RECT 3.185 2.085 3.405 2.465 ;
      RECT 3.575 0.255 3.925 0.765 ;
      RECT 3.575 0.765 4 0.935 ;
      RECT 3.575 0.935 3.745 1.575 ;
      RECT 3.575 1.575 4.04 1.745 ;
      RECT 3.575 2.255 5.53 2.635 ;
      RECT 3.915 1.105 4.46 1.275 ;
      RECT 4.095 0.085 4.425 0.445 ;
      RECT 4.17 0.615 4.825 0.785 ;
      RECT 4.17 0.785 4.46 1.105 ;
      RECT 4.21 1.275 4.46 1.495 ;
      RECT 4.21 1.495 5.01 1.745 ;
      RECT 4.595 0.255 4.825 0.615 ;
      RECT 5.1 0.255 5.31 0.615 ;
      RECT 5.1 0.615 6.4 0.785 ;
      RECT 5.18 1.435 5.65 1.605 ;
      RECT 5.18 1.605 5.49 1.915 ;
      RECT 5.49 0.085 6.4 0.445 ;
      RECT 5.7 1.775 6.4 2.085 ;
      RECT 5.7 2.085 5.87 2.465 ;
      RECT 5.82 1.435 6.4 1.775 ;
      RECT 6.07 2.255 6.4 2.635 ;
      RECT 6.23 0.785 6.4 0.995 ;
      RECT 6.23 0.995 6.5 1.325 ;
      RECT 6.23 1.325 6.4 1.435 ;
      RECT 7.01 0.085 7.275 0.885 ;
      RECT 7.01 1.485 7.275 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 1.445 1.7 1.615 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.99 0.765 2.16 0.935 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.83 0.765 4 0.935 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.29 1.445 4.46 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
    LAYER met1 ;
      RECT 1.47 1.415 1.76 1.46 ;
      RECT 1.47 1.46 4.52 1.6 ;
      RECT 1.47 1.6 1.76 1.645 ;
      RECT 1.93 0.735 2.22 0.78 ;
      RECT 1.93 0.78 4.06 0.92 ;
      RECT 1.93 0.92 2.22 0.965 ;
      RECT 3.77 0.735 4.06 0.78 ;
      RECT 3.77 0.92 4.06 0.965 ;
      RECT 4.23 1.415 4.52 1.46 ;
      RECT 4.23 1.6 4.52 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_2
MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.85 0.955 1.19 1.325 ;
        RECT 0.88 1.325 1.19 1.445 ;
        RECT 0.88 1.445 1.235 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.53 0.255 6.815 0.825 ;
        RECT 6.53 1.495 6.815 2.465 ;
        RECT 6.645 0.825 6.815 1.495 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.34 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.71 0.955 6.01 1.265 ;
        RECT 4.71 1.265 4.93 1.325 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.19 0.785 ;
      RECT 0.085 1.835 0.345 2.635 ;
      RECT 0.51 0.785 0.68 1.46 ;
      RECT 0.51 1.46 0.71 1.755 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.54 1.755 0.71 2.125 ;
      RECT 0.54 2.125 1.255 2.465 ;
      RECT 1.015 0.255 1.19 0.615 ;
      RECT 1.36 0.255 2.495 0.535 ;
      RECT 1.36 0.705 1.7 1.205 ;
      RECT 1.36 1.205 1.86 1.325 ;
      RECT 1.405 1.325 1.86 1.955 ;
      RECT 1.425 2.125 2.2 2.465 ;
      RECT 1.87 0.705 2.155 1.035 ;
      RECT 2.03 1.205 3.01 1.375 ;
      RECT 2.03 1.375 2.2 2.125 ;
      RECT 2.325 0.535 2.495 0.995 ;
      RECT 2.325 0.995 3.01 1.205 ;
      RECT 2.37 1.575 2.54 1.635 ;
      RECT 2.37 1.635 3.4 1.905 ;
      RECT 2.37 2.075 3.01 2.635 ;
      RECT 2.665 0.085 3.01 0.825 ;
      RECT 3.18 0.255 3.4 1.635 ;
      RECT 3.18 1.905 3.4 1.915 ;
      RECT 3.18 1.915 5.45 2.085 ;
      RECT 3.18 2.085 3.4 2.465 ;
      RECT 3.58 0.255 3.91 0.765 ;
      RECT 3.58 0.765 4.005 0.935 ;
      RECT 3.58 0.935 3.75 1.575 ;
      RECT 3.58 1.575 3.99 1.745 ;
      RECT 3.58 2.255 5.49 2.635 ;
      RECT 3.92 1.105 4.465 1.275 ;
      RECT 4.08 0.085 4.41 0.445 ;
      RECT 4.16 1.275 4.465 1.495 ;
      RECT 4.16 1.495 4.96 1.745 ;
      RECT 4.175 0.615 4.83 0.785 ;
      RECT 4.175 0.785 4.465 1.105 ;
      RECT 4.58 0.255 4.83 0.615 ;
      RECT 5.01 0.255 5.27 0.615 ;
      RECT 5.01 0.615 6.36 0.785 ;
      RECT 5.14 1.435 5.61 1.605 ;
      RECT 5.14 1.605 5.45 1.915 ;
      RECT 5.505 0.085 6.36 0.445 ;
      RECT 5.66 1.775 6.36 2.085 ;
      RECT 5.66 2.085 5.83 2.465 ;
      RECT 5.78 1.435 6.36 1.775 ;
      RECT 6.03 2.255 6.36 2.635 ;
      RECT 6.19 0.785 6.36 0.995 ;
      RECT 6.19 0.995 6.46 1.325 ;
      RECT 6.19 1.325 6.36 1.435 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 0.765 2.155 0.935 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.835 0.765 4.005 0.935 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.295 1.445 4.465 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.525 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 1.925 0.735 2.215 0.78 ;
      RECT 1.925 0.78 4.065 0.92 ;
      RECT 1.925 0.92 2.215 0.965 ;
      RECT 3.775 0.735 4.065 0.78 ;
      RECT 3.775 0.92 4.065 0.965 ;
      RECT 4.235 1.415 4.525 1.46 ;
      RECT 4.235 1.6 4.525 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_1
MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 0.995 2.01 1.445 ;
        RECT 1.84 1.445 2.275 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.28 0.995 1.61 1.45 ;
        RECT 1.4 1.45 1.61 1.785 ;
        RECT 1.4 1.785 1.72 2.375 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.88 0.995 1.05 1.62 ;
        RECT 0.88 1.62 1.23 2.375 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.37 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 1.455 4.055 1.625 ;
        RECT 2.48 1.625 2.73 2.465 ;
        RECT 2.52 0.255 2.77 0.725 ;
        RECT 2.52 0.725 4.055 0.905 ;
        RECT 3.28 0.255 3.61 0.725 ;
        RECT 3.32 1.625 3.57 2.465 ;
        RECT 3.81 0.905 4.055 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.115 1.495 0.71 1.665 ;
      RECT 0.115 1.665 0.45 2.45 ;
      RECT 0.12 0.085 0.37 0.585 ;
      RECT 0.54 0.655 2.35 0.825 ;
      RECT 0.54 0.825 0.71 1.495 ;
      RECT 0.7 0.305 0.87 0.655 ;
      RECT 1.07 0.085 1.4 0.485 ;
      RECT 1.57 0.305 1.74 0.655 ;
      RECT 1.96 0.085 2.34 0.485 ;
      RECT 2.005 1.795 2.255 2.635 ;
      RECT 2.18 0.825 2.35 1.075 ;
      RECT 2.18 1.075 3.64 1.245 ;
      RECT 2.9 1.795 3.15 2.635 ;
      RECT 2.94 0.085 3.11 0.555 ;
      RECT 3.74 1.795 3.99 2.635 ;
      RECT 3.78 0.085 3.95 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__or4_4
MACRO sky130_fd_sc_hd__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.32 1.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.44 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.68 0.76 ;
        RECT 2.405 1.495 2.68 2.465 ;
        RECT 2.51 0.76 2.68 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.495 0.41 1.785 ;
      RECT 0.085 1.785 1.68 1.955 ;
      RECT 0.09 0.085 0.425 0.585 ;
      RECT 0.625 0.305 0.795 0.655 ;
      RECT 0.625 0.655 2.235 0.825 ;
      RECT 0.995 0.085 1.325 0.485 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.51 1.495 2.235 1.665 ;
      RECT 1.51 1.665 1.68 1.785 ;
      RECT 1.835 0.085 2.215 0.485 ;
      RECT 1.915 1.835 2.195 2.635 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.34 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
      RECT 2.85 0.085 3.02 1 ;
      RECT 2.85 1.455 3.02 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__or4_2
MACRO sky130_fd_sc_hd__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.32 1.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.755 0.44 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 1.495 0.41 1.785 ;
      RECT 0.09 1.785 1.68 1.955 ;
      RECT 0.095 0.085 0.425 0.585 ;
      RECT 0.625 0.305 0.795 0.655 ;
      RECT 0.625 0.655 2.235 0.825 ;
      RECT 0.995 0.085 1.325 0.485 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.51 1.495 2.235 1.665 ;
      RECT 1.51 1.665 1.68 1.785 ;
      RECT 1.835 0.085 2.215 0.485 ;
      RECT 1.915 1.835 2.195 2.635 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.335 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__or4_1
MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.775 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.255 3.595 0.825 ;
        RECT 3.21 1.495 3.595 2.465 ;
        RECT 3.315 0.825 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.2 0.255 0.485 0.715 ;
      RECT 0.2 0.715 1.155 0.885 ;
      RECT 0.2 1.785 1.155 2.005 ;
      RECT 0.2 2.005 0.485 2.465 ;
      RECT 0.655 0.085 0.925 0.545 ;
      RECT 0.655 2.175 0.925 2.635 ;
      RECT 0.945 0.885 1.155 1.785 ;
      RECT 1.325 0.255 1.725 1.055 ;
      RECT 1.325 1.055 2.42 1.615 ;
      RECT 1.325 1.615 1.725 2.465 ;
      RECT 1.915 0.255 2.195 0.715 ;
      RECT 1.915 0.715 3.04 0.885 ;
      RECT 1.915 1.785 3.04 2.005 ;
      RECT 1.915 2.005 2.195 2.465 ;
      RECT 2.59 0.885 3.04 0.995 ;
      RECT 2.59 0.995 3.145 1.325 ;
      RECT 2.59 1.325 3.04 1.785 ;
      RECT 2.715 0.085 3.04 0.545 ;
      RECT 2.715 2.175 3.04 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345 0.895 2.155 1.275 ;
        RECT 8.93 0.895 10.71 1.275 ;
      LAYER mcon ;
        RECT 1.525 1.105 1.695 1.275 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 9.345 1.105 9.515 1.275 ;
        RECT 9.805 1.105 9.975 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 2.215 1.12 ;
        RECT 1.465 1.12 10.035 1.26 ;
        RECT 1.465 1.26 2.215 1.305 ;
        RECT 9.285 1.075 10.035 1.12 ;
        RECT 9.285 1.26 10.035 1.305 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.455 10.48 1.665 ;
        RECT 0.615 1.665 0.785 2.465 ;
        RECT 1.475 1.665 1.645 2.465 ;
        RECT 2.325 0.28 2.55 1.415 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.335 1.665 2.505 2.465 ;
        RECT 3.155 0.28 3.41 1.415 ;
        RECT 3.195 1.665 3.365 2.465 ;
        RECT 4.015 0.28 4.255 1.415 ;
        RECT 4.055 1.665 4.225 2.465 ;
        RECT 4.905 0.28 5.255 1.415 ;
        RECT 5.08 1.665 5.25 2.465 ;
        RECT 5.925 0.28 6.175 1.415 ;
        RECT 5.965 1.665 6.135 2.465 ;
        RECT 6.785 0.28 7.035 1.415 ;
        RECT 6.825 1.665 6.995 2.465 ;
        RECT 7.645 0.28 7.895 1.415 ;
        RECT 7.685 1.665 7.855 2.465 ;
        RECT 8.505 0.28 8.755 1.415 ;
        RECT 8.545 1.665 8.715 2.465 ;
        RECT 9.405 1.665 9.575 2.465 ;
        RECT 10.265 1.665 10.435 2.465 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.495 0.44 2.465 ;
        RECT 10.61 1.835 10.94 2.465 ;
      LAYER mcon ;
        RECT 0.13 2.125 0.3 2.295 ;
        RECT 10.72 2.125 10.89 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.965 1.835 1.295 2.465 ;
      LAYER mcon ;
        RECT 0.99 2.125 1.16 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.825 1.835 2.155 2.465 ;
      LAYER mcon ;
        RECT 1.89 2.125 2.06 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685 1.835 3.015 2.465 ;
      LAYER mcon ;
        RECT 2.77 2.125 2.94 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.545 1.835 3.875 2.465 ;
      LAYER mcon ;
        RECT 3.69 2.125 3.86 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.425 1.835 4.755 2.465 ;
      LAYER mcon ;
        RECT 4.55 2.125 4.72 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.45 1.835 5.78 2.465 ;
      LAYER mcon ;
        RECT 5.45 2.125 5.62 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.315 1.835 6.645 2.465 ;
      LAYER mcon ;
        RECT 6.37 2.125 6.54 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.175 1.835 7.505 2.465 ;
      LAYER mcon ;
        RECT 7.23 2.125 7.4 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.035 1.835 8.365 2.465 ;
      LAYER mcon ;
        RECT 8.13 2.125 8.3 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.895 1.835 9.225 2.465 ;
      LAYER mcon ;
        RECT 8.96 2.125 9.13 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 1.835 10.085 2.465 ;
      LAYER mcon ;
        RECT 9.82 2.125 9.99 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.08 0.36 2.14 ;
        RECT 0.07 2.14 10.97 2.34 ;
        RECT 0.93 2.08 1.22 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.71 2.08 3 2.14 ;
        RECT 3.63 2.08 3.92 2.14 ;
        RECT 4.49 2.08 4.78 2.14 ;
        RECT 5.39 2.08 5.68 2.14 ;
        RECT 6.31 2.08 6.6 2.14 ;
        RECT 7.17 2.08 7.46 2.14 ;
        RECT 8.07 2.08 8.36 2.14 ;
        RECT 8.9 2.08 9.19 2.14 ;
        RECT 9.76 2.08 10.05 2.14 ;
        RECT 10.66 2.08 10.95 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 1.855 0.085 2.125 0.61 ;
      RECT 2.72 0.085 2.985 0.61 ;
      RECT 3.58 0.085 3.845 0.61 ;
      RECT 4.465 0.085 4.73 0.61 ;
      RECT 5.49 0.085 5.755 0.61 ;
      RECT 6.35 0.085 6.575 0.61 ;
      RECT 7.21 0.085 7.475 0.61 ;
      RECT 8.07 0.085 8.335 0.61 ;
      RECT 8.93 0.085 9.195 0.61 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.46 1.755 1.63 ;
        RECT 0.155 1.63 0.375 2.435 ;
        RECT 1.025 0.28 1.25 0.725 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.045 1.63 1.235 2.435 ;
        RECT 1.475 0.895 1.755 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.8 0.875 2.465 ;
      LAYER mcon ;
        RECT 0.6 2.125 0.77 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.405 1.8 1.735 2.465 ;
      LAYER mcon ;
        RECT 1.5 2.125 1.67 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.54 2.08 0.83 2.14 ;
        RECT 1.44 2.08 1.73 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.56 0.085 0.855 0.61 ;
      RECT 1.42 0.085 1.75 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.66 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 0.105 0.895 0.275 1.46 ;
        RECT 0.105 1.46 3.135 1.63 ;
        RECT 0.645 1.63 0.815 2.435 ;
        RECT 1.03 0.28 1.29 0.725 ;
        RECT 1.505 1.63 1.675 2.435 ;
        RECT 1.89 0.28 2.145 0.725 ;
        RECT 2.365 1.63 2.535 2.435 ;
        RECT 2.835 0.895 3.135 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.8 0.465 2.465 ;
      LAYER mcon ;
        RECT 0.195 2.125 0.365 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.995 1.8 1.325 2.465 ;
      LAYER mcon ;
        RECT 1.055 2.125 1.225 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.855 1.8 2.185 2.465 ;
      LAYER mcon ;
        RECT 1.955 2.125 2.125 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.715 1.8 3.045 2.465 ;
      LAYER mcon ;
        RECT 2.835 2.125 3.005 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 3.15 2.34 ;
        RECT 0.135 2.08 0.425 2.14 ;
        RECT 0.995 2.08 1.285 2.14 ;
        RECT 1.895 2.08 2.185 2.14 ;
        RECT 2.775 2.08 3.065 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.565 0.085 0.86 0.555 ;
      RECT 1.46 0.085 1.72 0.555 ;
      RECT 2.315 0.085 2.615 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.255 0.84 0.76 ;
        RECT 0.59 0.76 1.295 0.945 ;
        RECT 0.595 0.945 1.295 1.29 ;
        RECT 0.595 1.29 0.765 2.465 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.665 0.425 2.465 ;
      LAYER mcon ;
        RECT 0.155 2.125 0.325 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.935 1.665 1.295 2.465 ;
      LAYER mcon ;
        RECT 1.055 2.125 1.225 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.095 2.08 0.385 2.14 ;
        RECT 0.995 2.08 1.285 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 1.01 0.085 1.295 0.59 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.695 5.44 0.865 ;
        RECT 0.115 0.865 0.285 1.46 ;
        RECT 0.115 1.46 5.44 1.63 ;
        RECT 0.595 1.63 0.765 2.435 ;
        RECT 1.44 1.63 1.61 2.435 ;
        RECT 1.535 0.28 1.725 0.695 ;
        RECT 2.28 1.63 2.45 2.435 ;
        RECT 2.395 0.28 2.585 0.695 ;
        RECT 3.12 1.63 3.29 2.435 ;
        RECT 3.255 0.28 3.445 0.695 ;
        RECT 3.96 1.63 4.13 2.435 ;
        RECT 4.115 0.28 4.305 0.695 ;
        RECT 4.8 1.63 4.97 2.435 ;
        RECT 5.17 0.865 5.44 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.8 0.425 2.465 ;
        RECT 5.14 1.8 5.47 2.465 ;
      LAYER mcon ;
        RECT 0.13 2.125 0.3 2.295 ;
        RECT 5.255 2.125 5.425 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.94 1.8 1.27 2.465 ;
      LAYER mcon ;
        RECT 0.99 2.125 1.16 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.78 1.8 2.11 2.465 ;
      LAYER mcon ;
        RECT 1.89 2.125 2.06 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.62 1.8 2.95 2.465 ;
      LAYER mcon ;
        RECT 2.77 2.125 2.94 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.46 1.8 3.79 2.465 ;
      LAYER mcon ;
        RECT 3.495 2.125 3.665 2.295 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.3 1.8 4.63 2.465 ;
      LAYER mcon ;
        RECT 4.355 2.125 4.525 2.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.08 0.36 2.14 ;
        RECT 0.07 2.14 5.91 2.34 ;
        RECT 0.93 2.08 1.22 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.71 2.08 3 2.14 ;
        RECT 3.435 2.08 3.725 2.14 ;
        RECT 4.295 2.08 4.585 2.14 ;
        RECT 5.195 2.08 5.485 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 1.035 0.085 1.365 0.525 ;
      RECT 1.895 0.085 2.225 0.525 ;
      RECT 2.755 0.085 3.085 0.525 ;
      RECT 3.615 0.085 3.945 0.525 ;
      RECT 4.475 0.085 4.805 0.525 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8
MACRO sky130_fd_sc_hd__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.5 1.075 3.08 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.415 2.33 2.355 ;
        RECT 2 1.075 2.33 1.415 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 1.075 1.83 1.245 ;
        RECT 1.5 1.245 1.82 2.355 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.075 1.32 1.245 ;
        RECT 1.015 1.245 1.32 2.355 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.44 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.735 ;
        RECT 0.085 0.735 0.78 0.905 ;
        RECT 0.515 1.485 0.845 2.465 ;
        RECT 0.61 0.905 0.78 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.445 0.345 2.635 ;
      RECT 0.79 0.255 1.12 0.565 ;
      RECT 0.95 0.565 1.12 0.735 ;
      RECT 0.95 0.735 2.96 0.905 ;
      RECT 1.29 0.085 1.54 0.565 ;
      RECT 1.71 0.255 2.04 0.735 ;
      RECT 2.21 0.085 2.46 0.565 ;
      RECT 2.63 0.255 2.96 0.735 ;
      RECT 2.63 1.495 2.96 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o41ai_1
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.17 1.075 7.94 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.31 1.075 5.98 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.075 4.02 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.7 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 2.16 0.905 ;
        RECT 0.515 1.445 3.885 1.615 ;
        RECT 0.515 1.615 0.845 2.465 ;
        RECT 1.355 1.615 1.685 2.465 ;
        RECT 1.87 0.905 2.16 1.445 ;
        RECT 2.715 1.615 3.045 2.125 ;
        RECT 3.555 1.615 3.885 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.085 0.255 2.625 0.465 ;
      RECT 0.085 0.465 0.345 0.905 ;
      RECT 0.085 1.445 0.345 2.635 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.855 1.835 2.105 2.635 ;
      RECT 2.295 1.785 2.545 2.295 ;
      RECT 2.295 2.295 4.225 2.465 ;
      RECT 2.35 0.465 2.625 0.735 ;
      RECT 2.35 0.735 9.865 0.905 ;
      RECT 2.795 0.085 2.965 0.545 ;
      RECT 3.135 0.255 3.465 0.735 ;
      RECT 3.215 1.785 3.385 2.295 ;
      RECT 3.635 0.085 3.805 0.545 ;
      RECT 3.975 0.255 4.305 0.735 ;
      RECT 4.055 1.445 5.985 1.615 ;
      RECT 4.055 1.615 4.225 2.295 ;
      RECT 4.395 1.785 4.645 2.295 ;
      RECT 4.395 2.295 7.685 2.465 ;
      RECT 4.475 0.085 4.645 0.545 ;
      RECT 4.815 0.255 5.145 0.735 ;
      RECT 4.815 1.615 5.145 2.125 ;
      RECT 5.315 0.085 5.485 0.545 ;
      RECT 5.315 1.785 5.485 2.295 ;
      RECT 5.655 0.255 5.985 0.735 ;
      RECT 5.655 1.615 5.985 2.125 ;
      RECT 6.175 0.26 6.505 0.735 ;
      RECT 6.175 1.445 9.865 1.615 ;
      RECT 6.175 1.615 6.505 2.125 ;
      RECT 6.675 0.085 6.845 0.545 ;
      RECT 6.675 1.785 6.845 2.295 ;
      RECT 7.015 0.26 7.345 0.735 ;
      RECT 7.015 1.615 7.345 2.125 ;
      RECT 7.515 0.085 7.685 0.545 ;
      RECT 7.515 1.785 7.685 2.295 ;
      RECT 7.855 0.26 8.185 0.735 ;
      RECT 7.855 1.615 8.185 2.465 ;
      RECT 8.355 0.085 8.525 0.545 ;
      RECT 8.355 1.835 8.525 2.635 ;
      RECT 8.695 0.26 9.025 0.735 ;
      RECT 8.695 1.615 9.025 2.465 ;
      RECT 9.195 0.085 9.365 0.545 ;
      RECT 9.195 1.835 9.365 2.635 ;
      RECT 9.535 0.26 9.865 0.735 ;
      RECT 9.535 1.615 9.865 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__o41ai_4
MACRO sky130_fd_sc_hd__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.72 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 1.075 4.54 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595 1.075 3.58 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 1.075 2.325 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.44 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 0.845 0.885 ;
        RECT 0.515 1.505 2.205 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 0.61 0.885 0.845 1.445 ;
        RECT 0.61 1.445 2.205 1.505 ;
        RECT 1.875 1.665 2.205 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.255 1.265 0.465 ;
      RECT 0.085 0.465 0.345 0.905 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 1.015 0.465 1.265 0.735 ;
      RECT 1.015 0.735 5.705 0.905 ;
      RECT 1.015 1.835 1.265 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.455 1.835 1.705 2.295 ;
      RECT 1.455 2.295 2.545 2.465 ;
      RECT 1.875 0.255 2.205 0.735 ;
      RECT 2.375 0.085 2.545 0.545 ;
      RECT 2.375 1.445 3.465 1.615 ;
      RECT 2.375 1.615 2.545 2.295 ;
      RECT 2.715 0.255 3.045 0.735 ;
      RECT 2.715 1.835 3.045 2.295 ;
      RECT 2.715 2.295 4.445 2.465 ;
      RECT 3.215 0.085 3.45 0.545 ;
      RECT 3.215 1.615 3.465 2.125 ;
      RECT 3.695 0.255 4.025 0.735 ;
      RECT 3.695 1.445 5.705 1.615 ;
      RECT 3.695 1.615 3.945 2.125 ;
      RECT 4.115 1.835 4.445 2.295 ;
      RECT 4.195 0.085 4.365 0.545 ;
      RECT 4.535 0.255 4.865 0.735 ;
      RECT 4.615 1.615 4.785 2.465 ;
      RECT 4.955 1.785 5.285 2.635 ;
      RECT 5.035 0.085 5.205 0.545 ;
      RECT 5.375 0.255 5.705 0.735 ;
      RECT 5.455 1.615 5.705 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__o41ai_2
MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.43 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.97 0.62 1.305 0.995 ;
        RECT 0.97 0.995 1.43 1.325 ;
        RECT 0.97 1.325 1.305 1.695 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.445 9.575 1.725 ;
        RECT 6.275 0.615 9.575 0.855 ;
        RECT 9.325 0.855 9.575 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.085 0.085 0.445 0.825 ;
      RECT 0.085 1.785 0.445 2.635 ;
      RECT 0.6 0.995 0.8 1.615 ;
      RECT 0.615 0.28 0.8 0.995 ;
      RECT 0.615 1.615 0.8 2.465 ;
      RECT 0.97 0.085 1.305 0.445 ;
      RECT 0.97 1.865 1.305 2.635 ;
      RECT 1.475 0.255 1.985 0.825 ;
      RECT 1.475 1.495 1.825 2.465 ;
      RECT 1.6 0.825 1.985 1.025 ;
      RECT 1.6 1.025 5.925 1.275 ;
      RECT 1.6 1.275 1.825 1.495 ;
      RECT 1.995 1.895 9.575 2.065 ;
      RECT 1.995 2.065 2.245 2.465 ;
      RECT 2.155 0.255 2.485 0.655 ;
      RECT 2.155 0.655 6.105 0.855 ;
      RECT 2.415 2.235 2.745 2.635 ;
      RECT 2.655 0.085 2.985 0.485 ;
      RECT 2.915 2.065 3.085 2.465 ;
      RECT 3.155 0.275 3.325 0.655 ;
      RECT 3.255 2.235 3.585 2.635 ;
      RECT 3.495 0.085 3.825 0.485 ;
      RECT 3.755 2.065 3.925 2.465 ;
      RECT 3.995 0.255 4.165 0.655 ;
      RECT 4.095 2.235 4.425 2.635 ;
      RECT 4.335 0.085 4.665 0.485 ;
      RECT 4.595 2.065 4.765 2.465 ;
      RECT 4.835 0.275 5.005 0.655 ;
      RECT 4.935 2.235 5.265 2.635 ;
      RECT 5.175 0.085 5.505 0.485 ;
      RECT 5.435 2.065 9.575 2.465 ;
      RECT 5.675 0.255 9.575 0.445 ;
      RECT 5.675 0.445 6.105 0.655 ;
      RECT 6.175 1.025 9.155 1.275 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 1.105 0.775 1.275 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.58 1.105 6.75 1.275 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.545 1.075 0.835 1.12 ;
      RECT 0.545 1.12 6.81 1.26 ;
      RECT 0.545 1.26 0.835 1.305 ;
      RECT 6.52 1.075 6.81 1.12 ;
      RECT 6.52 1.26 6.81 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_8
MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 0.765 0.78 1.675 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.765 1.28 1.425 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 1.445 5.895 1.725 ;
        RECT 4.145 0.615 5.895 0.855 ;
        RECT 5.675 0.855 5.895 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.28 0.345 0.665 ;
      RECT 0.085 0.665 0.32 1.765 ;
      RECT 0.085 1.765 0.345 2.465 ;
      RECT 0.515 0.085 0.93 0.595 ;
      RECT 0.515 1.845 0.93 2.635 ;
      RECT 1.1 0.255 1.725 0.595 ;
      RECT 1.1 1.595 1.725 1.765 ;
      RECT 1.1 1.765 1.355 2.465 ;
      RECT 1.45 0.595 1.725 1.025 ;
      RECT 1.45 1.025 3.81 1.275 ;
      RECT 1.45 1.275 1.725 1.595 ;
      RECT 1.565 1.935 5.895 2.105 ;
      RECT 1.565 2.105 1.81 2.465 ;
      RECT 1.895 0.255 2.175 0.655 ;
      RECT 1.895 0.655 3.975 0.855 ;
      RECT 1.895 1.895 5.895 1.935 ;
      RECT 1.98 2.275 2.31 2.635 ;
      RECT 2.345 0.085 2.675 0.485 ;
      RECT 2.48 2.105 2.65 2.465 ;
      RECT 2.82 2.275 3.15 2.635 ;
      RECT 2.845 0.275 3.015 0.655 ;
      RECT 3.185 0.085 3.515 0.485 ;
      RECT 3.32 2.105 5.895 2.465 ;
      RECT 3.685 0.255 5.735 0.445 ;
      RECT 3.685 0.445 3.975 0.655 ;
      RECT 3.98 1.025 5.505 1.275 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.15 1.105 0.32 1.275 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.31 1.105 4.48 1.275 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 0.085 1.075 0.38 1.12 ;
      RECT 0.085 1.12 4.54 1.26 ;
      RECT 0.085 1.26 0.38 1.305 ;
      RECT 4.25 1.075 4.54 1.12 ;
      RECT 4.25 1.26 4.54 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_4
MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.355 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 1.075 1.24 1.63 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.601000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.495 3.595 2.465 ;
        RECT 3.125 0.255 3.595 0.825 ;
        RECT 3.255 0.825 3.595 1.495 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.28 0.345 0.615 ;
      RECT 0.085 0.615 1.185 0.825 ;
      RECT 0.085 1.785 0.74 2.005 ;
      RECT 0.085 2.005 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.445 ;
      RECT 0.515 2.175 0.845 2.635 ;
      RECT 0.525 0.825 0.74 1.785 ;
      RECT 1.015 0.255 2.025 0.465 ;
      RECT 1.015 0.465 1.185 0.615 ;
      RECT 1.015 1.8 1.805 2.005 ;
      RECT 1.015 2.005 1.27 2.46 ;
      RECT 1.355 0.635 1.685 0.885 ;
      RECT 1.41 0.885 1.685 1.075 ;
      RECT 1.41 1.075 2.535 1.325 ;
      RECT 1.41 1.325 1.805 1.8 ;
      RECT 1.44 2.175 1.805 2.635 ;
      RECT 1.855 0.465 2.025 0.735 ;
      RECT 1.855 0.735 2.955 0.905 ;
      RECT 2.195 0.085 2.955 0.565 ;
      RECT 2.705 0.905 2.955 0.995 ;
      RECT 2.705 0.995 3.085 1.325 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__ebufn_1
MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 0.765 0.78 1.675 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.765 1.28 1.275 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905 1.445 4.055 1.625 ;
        RECT 1.905 1.625 3.625 1.765 ;
        RECT 3.295 0.635 4.055 0.855 ;
        RECT 3.295 1.765 3.625 2.125 ;
        RECT 3.825 0.855 4.055 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.28 0.345 0.615 ;
      RECT 0.085 0.615 0.32 1.845 ;
      RECT 0.085 1.845 0.345 2.465 ;
      RECT 0.515 0.085 0.85 0.595 ;
      RECT 0.515 1.845 0.95 2.635 ;
      RECT 1.02 0.255 1.73 0.595 ;
      RECT 1.12 1.445 1.735 1.765 ;
      RECT 1.12 1.765 1.41 2.465 ;
      RECT 1.45 0.595 1.73 1.025 ;
      RECT 1.45 1.025 2.965 1.275 ;
      RECT 1.45 1.275 1.735 1.445 ;
      RECT 1.6 1.935 3.125 2.105 ;
      RECT 1.6 2.105 1.81 2.465 ;
      RECT 1.9 0.255 2.17 0.655 ;
      RECT 1.9 0.655 3.125 0.855 ;
      RECT 1.98 2.275 2.31 2.635 ;
      RECT 2.34 0.085 2.67 0.485 ;
      RECT 2.48 2.105 3.125 2.295 ;
      RECT 2.48 2.295 4.055 2.465 ;
      RECT 2.84 0.275 4.05 0.465 ;
      RECT 2.84 0.465 3.125 0.655 ;
      RECT 3.245 1.025 3.655 1.275 ;
      RECT 3.795 1.795 4.055 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.15 1.105 0.32 1.275 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.38 1.105 3.55 1.275 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
    LAYER met1 ;
      RECT 0.085 1.075 0.38 1.12 ;
      RECT 0.085 1.12 3.61 1.26 ;
      RECT 0.085 1.26 0.38 1.305 ;
      RECT 3.32 1.075 3.61 1.12 ;
      RECT 3.32 1.26 3.61 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_2
MACRO sky130_fd_sc_hd__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.635 1.075 3.075 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.075 2.465 1.285 ;
        RECT 1.98 1.285 2.285 1.705 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.075 1.23 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.4 1.075 1.79 1.275 ;
        RECT 1.5 1.275 1.79 1.705 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.345 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295 0.265 3.625 0.735 ;
        RECT 3.295 0.735 4.055 0.905 ;
        RECT 3.295 1.875 4.055 2.045 ;
        RECT 3.295 2.045 3.545 2.465 ;
        RECT 3.745 0.905 4.055 1.875 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.12 -0.085 0.29 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.17 0.255 0.5 0.635 ;
      RECT 0.17 0.635 0.715 0.805 ;
      RECT 0.25 1.495 1.33 1.67 ;
      RECT 0.25 1.67 0.58 2.465 ;
      RECT 0.545 0.805 0.715 1.445 ;
      RECT 0.545 1.445 1.33 1.495 ;
      RECT 0.67 0.295 1.855 0.465 ;
      RECT 0.75 1.85 0.99 2.635 ;
      RECT 1.085 0.645 1.47 0.735 ;
      RECT 1.085 0.735 2.785 0.905 ;
      RECT 1.16 1.67 1.33 1.875 ;
      RECT 1.16 1.875 2.625 2.045 ;
      RECT 1.55 2.045 2.305 2.465 ;
      RECT 2.115 0.085 2.285 0.555 ;
      RECT 2.455 0.27 2.785 0.735 ;
      RECT 2.455 1.455 3.415 1.625 ;
      RECT 2.455 1.625 2.625 1.875 ;
      RECT 2.795 1.795 3.125 2.635 ;
      RECT 2.955 0.085 3.125 0.905 ;
      RECT 3.245 1.075 3.575 1.285 ;
      RECT 3.245 1.285 3.415 1.455 ;
      RECT 3.715 2.215 4.055 2.635 ;
      RECT 3.795 0.085 3.965 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o221a_2
MACRO sky130_fd_sc_hd__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.075 3.605 1.445 ;
        RECT 3.005 1.445 4.775 1.615 ;
        RECT 4.525 1.075 5.035 1.275 ;
        RECT 4.525 1.275 4.775 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 4.355 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.075 1.52 1.445 ;
        RECT 1.025 1.445 2.745 1.615 ;
        RECT 2.415 1.075 2.745 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.69 1.075 2.245 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 5.235 0.725 6.405 0.735 ;
        RECT 5.235 0.735 6.92 0.905 ;
        RECT 5.315 1.785 5.9 1.955 ;
        RECT 5.315 1.955 5.525 2.465 ;
        RECT 5.73 1.445 6.92 1.615 ;
        RECT 5.73 1.615 5.9 1.785 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.115 1.615 6.365 2.465 ;
        RECT 6.575 0.905 6.92 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.085 0.255 2.955 0.475 ;
      RECT 0.085 0.475 0.345 0.895 ;
      RECT 0.145 1.455 0.395 2.635 ;
      RECT 0.515 0.645 0.845 0.865 ;
      RECT 0.565 1.445 0.845 1.785 ;
      RECT 0.565 1.785 5.145 1.955 ;
      RECT 0.565 1.955 0.815 2.465 ;
      RECT 0.61 0.865 0.845 1.445 ;
      RECT 0.985 2.125 1.235 2.635 ;
      RECT 1.015 0.475 1.185 0.905 ;
      RECT 1.355 0.645 2.535 0.715 ;
      RECT 1.355 0.715 3.885 0.725 ;
      RECT 1.355 0.725 4.725 0.905 ;
      RECT 1.405 2.125 1.655 2.295 ;
      RECT 1.405 2.295 2.495 2.465 ;
      RECT 1.825 1.955 2.075 2.125 ;
      RECT 2.245 2.125 2.495 2.295 ;
      RECT 2.665 2.125 3.425 2.635 ;
      RECT 3.145 0.085 3.385 0.545 ;
      RECT 3.555 0.255 3.885 0.715 ;
      RECT 3.595 2.125 3.845 2.295 ;
      RECT 3.595 2.295 4.685 2.465 ;
      RECT 4.015 1.955 4.265 2.125 ;
      RECT 4.055 0.085 4.225 0.555 ;
      RECT 4.395 0.255 4.725 0.725 ;
      RECT 4.435 2.125 4.685 2.295 ;
      RECT 4.855 2.125 5.105 2.635 ;
      RECT 4.895 0.085 5.065 0.905 ;
      RECT 4.975 1.445 5.375 1.615 ;
      RECT 4.975 1.615 5.145 1.785 ;
      RECT 5.205 1.075 6.405 1.275 ;
      RECT 5.205 1.275 5.375 1.445 ;
      RECT 5.695 2.125 5.945 2.635 ;
      RECT 5.735 0.085 5.905 0.555 ;
      RECT 6.535 1.795 6.785 2.635 ;
      RECT 6.575 0.085 6.83 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__o221a_4
MACRO sky130_fd_sc_hd__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 1.075 3.13 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.075 2.49 1.285 ;
        RECT 2.005 1.285 2.38 1.705 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925 1.075 1.255 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.075 1.815 1.325 ;
        RECT 1.495 1.325 1.815 1.705 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.415 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.37 0.265 4.055 0.905 ;
        RECT 3.39 1.875 4.055 2.465 ;
        RECT 3.805 0.905 4.055 1.875 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.24 1.455 1.325 1.625 ;
      RECT 0.24 1.625 0.54 2.465 ;
      RECT 0.245 0.255 0.575 0.645 ;
      RECT 0.245 0.645 0.755 0.825 ;
      RECT 0.585 0.825 0.755 1.455 ;
      RECT 0.735 1.795 0.985 2.635 ;
      RECT 0.745 0.305 1.93 0.475 ;
      RECT 1.155 1.625 1.325 1.875 ;
      RECT 1.155 1.875 2.72 2.045 ;
      RECT 1.16 0.645 1.545 0.735 ;
      RECT 1.16 0.735 2.86 0.905 ;
      RECT 1.575 2.045 2.38 2.465 ;
      RECT 2.19 0.085 2.36 0.555 ;
      RECT 2.53 0.27 2.86 0.735 ;
      RECT 2.55 1.455 3.47 1.625 ;
      RECT 2.55 1.625 2.72 1.875 ;
      RECT 2.89 1.795 3.22 2.635 ;
      RECT 3.03 0.085 3.2 0.905 ;
      RECT 3.3 1.075 3.635 1.285 ;
      RECT 3.3 1.285 3.47 1.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o221a_1
MACRO sky130_fd_sc_hd__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 2.095000 0.375000 2.325000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.125000 0.315000 2.295000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.29 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.17 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 5.925 4.595 6.095 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 6.17 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 5.87 3.455 6.16 3.5 ;
        RECT 5.87 3.64 6.16 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 6.63 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 6.44 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.29 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.29 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 6.44 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.865 0.085 6.155 0.81 ;
      RECT 5.865 2.985 6.155 3.955 ;
      RECT 5.865 4.63 6.155 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 5.93 3.485 6.1 3.655 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 6.44 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
      RECT 5.925 0.32 6.095 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 7.045 4.595 7.215 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 7.29 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 6.93 3.455 7.22 3.5 ;
        RECT 6.93 3.64 7.22 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 7.405 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 7.36 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 7.36 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.825 0.085 6.155 0.845 ;
      RECT 5.905 1.61 6.075 2.635 ;
      RECT 6.755 0.085 7.005 0.925 ;
      RECT 6.755 1.61 6.935 2.635 ;
      RECT 6.985 2.985 7.275 3.955 ;
      RECT 6.985 4.63 7.275 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.585 5.355 6.755 5.525 ;
      RECT 6.99 3.485 7.16 3.655 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.045 5.355 7.215 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 7.36 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
      LAYER mcon ;
        RECT 1.42 2.115 1.59 2.285 ;
        RECT 1.78 2.115 1.95 2.285 ;
        RECT 2.14 2.115 2.31 2.285 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.37 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
      LAYER nwell ;
        RECT 1.92 1.305 2.98 4.135 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
      LAYER pwell ;
        RECT 0.145 4.595 0.315 5.12 ;
        RECT 6.125 4.595 6.295 5.12 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.5 6.3 3.64 ;
        RECT 0.08 3.455 0.37 3.5 ;
        RECT 0.08 3.64 0.37 3.685 ;
        RECT 6.01 3.455 6.3 3.5 ;
        RECT 6.01 3.64 6.3 3.685 ;
      LAYER nwell ;
        RECT -0.19 1.305 0.65 4.135 ;
        RECT 4.25 1.305 6.63 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 1.89 2.805 ;
      RECT 0 5.355 6.44 5.525 ;
      RECT 0.085 0.085 0.375 0.81 ;
      RECT 0.085 2.985 0.375 3.97 ;
      RECT 0.085 4.63 0.375 5.355 ;
      RECT 2.02 0.085 2.35 0.895 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 2.645 4.515 2.905 5.355 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.115 0.085 3.445 0.9 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.575 4.515 3.765 5.355 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 3.975 0.085 4.305 0.56 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.445 4.515 4.955 5.355 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 4.835 0.085 5.165 0.9 ;
      RECT 4.89 1.625 5.12 2.635 ;
      RECT 4.89 2.635 6.44 2.805 ;
      RECT 4.89 2.805 5.12 3.74 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
      RECT 5.825 0.085 6.155 0.9 ;
      RECT 5.905 1.61 6.075 2.635 ;
      RECT 6.065 2.985 6.355 3.955 ;
      RECT 6.065 4.63 6.355 5.355 ;
    LAYER mcon ;
      RECT 0.14 3.485 0.31 3.655 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 6.07 3.485 6.24 3.655 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
    LAYER met1 ;
      RECT 0 -0.24 6.44 0.24 ;
    LAYER pwell ;
      RECT 0.145 0.32 0.315 0.845 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.375 1.075 9.11 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 1.075 7.105 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.445 1.365 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.075 1.295 1.325 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 1.415 3.185 1.705 ;
        RECT 1.935 0.255 2.265 0.725 ;
        RECT 1.935 0.725 8.665 0.905 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.015 0.905 3.185 1.415 ;
        RECT 3.615 0.255 3.945 0.725 ;
        RECT 4.455 0.255 4.785 0.725 ;
        RECT 5.815 0.255 6.145 0.725 ;
        RECT 6.655 0.255 6.985 0.725 ;
        RECT 7.495 0.255 7.825 0.725 ;
        RECT 8.335 0.255 8.665 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.085 0.255 0.445 0.725 ;
      RECT 0.085 0.725 0.785 0.895 ;
      RECT 0.085 1.535 0.785 1.875 ;
      RECT 0.085 1.875 3.525 2.045 ;
      RECT 0.085 2.045 0.365 2.465 ;
      RECT 0.535 2.215 0.865 2.635 ;
      RECT 0.615 0.085 0.785 0.555 ;
      RECT 0.615 0.895 0.785 1.535 ;
      RECT 0.955 0.255 1.285 0.735 ;
      RECT 0.955 0.735 1.635 0.905 ;
      RECT 0.955 1.535 1.635 1.705 ;
      RECT 1.465 0.905 1.635 1.075 ;
      RECT 1.465 1.075 2.845 1.245 ;
      RECT 1.465 1.245 1.635 1.535 ;
      RECT 1.515 2.215 3.525 2.295 ;
      RECT 1.515 2.295 5.195 2.465 ;
      RECT 1.595 0.085 1.765 0.555 ;
      RECT 2.435 0.085 2.605 0.555 ;
      RECT 3.275 0.085 3.445 0.555 ;
      RECT 3.355 1.075 4.905 1.285 ;
      RECT 3.355 1.285 3.525 1.875 ;
      RECT 3.695 1.455 6.945 1.625 ;
      RECT 3.695 1.625 3.905 2.125 ;
      RECT 4.075 1.795 4.325 2.295 ;
      RECT 4.115 0.085 4.285 0.555 ;
      RECT 4.495 1.625 4.745 2.125 ;
      RECT 4.915 1.795 5.195 2.295 ;
      RECT 4.955 0.085 5.645 0.555 ;
      RECT 5.38 1.795 5.685 2.295 ;
      RECT 5.38 2.295 7.365 2.465 ;
      RECT 5.855 1.625 6.105 2.125 ;
      RECT 6.275 1.795 6.525 2.295 ;
      RECT 6.315 0.085 6.485 0.555 ;
      RECT 6.695 1.625 6.945 2.125 ;
      RECT 7.115 1.455 9.11 1.625 ;
      RECT 7.115 1.625 7.365 2.295 ;
      RECT 7.155 0.085 7.325 0.555 ;
      RECT 7.535 1.795 7.785 2.635 ;
      RECT 7.955 1.625 8.205 2.465 ;
      RECT 7.995 0.085 8.165 0.555 ;
      RECT 8.375 1.795 8.625 2.635 ;
      RECT 8.795 1.625 9.11 2.465 ;
      RECT 8.835 0.085 9.11 0.905 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
  END
END sky130_fd_sc_hd__nor4bb_4
MACRO sky130_fd_sc_hd__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.13 1.075 5.895 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.96 1.275 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.235 1.325 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.78 1.695 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.06 0.255 2.39 0.725 ;
        RECT 2.06 0.725 5.45 0.905 ;
        RECT 2.9 0.255 3.23 0.725 ;
        RECT 2.9 1.445 3.995 1.705 ;
        RECT 3.575 0.905 3.995 1.445 ;
        RECT 4.28 0.255 4.61 0.725 ;
        RECT 5.12 0.255 5.45 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.45 0.465 0.825 ;
      RECT 0.085 0.825 0.255 1.885 ;
      RECT 0.085 1.885 1.915 2.055 ;
      RECT 0.085 2.055 0.345 2.455 ;
      RECT 0.515 2.24 0.845 2.635 ;
      RECT 0.635 0.085 0.805 0.825 ;
      RECT 0.995 1.525 1.575 1.715 ;
      RECT 1.055 0.45 1.25 0.655 ;
      RECT 1.055 0.655 1.575 0.825 ;
      RECT 1.405 0.825 1.575 1.075 ;
      RECT 1.405 1.075 2.39 1.245 ;
      RECT 1.405 1.245 1.575 1.525 ;
      RECT 1.56 0.085 1.89 0.48 ;
      RECT 1.64 2.225 1.97 2.295 ;
      RECT 1.64 2.295 3.65 2.465 ;
      RECT 1.745 1.415 2.73 1.585 ;
      RECT 1.745 1.585 1.915 1.885 ;
      RECT 2.14 1.795 2.31 1.875 ;
      RECT 2.14 1.875 4.61 2.045 ;
      RECT 2.14 2.045 2.31 2.125 ;
      RECT 2.48 2.215 3.65 2.295 ;
      RECT 2.56 0.085 2.73 0.555 ;
      RECT 2.56 1.075 3.405 1.275 ;
      RECT 2.56 1.275 2.73 1.415 ;
      RECT 3.4 0.085 4.11 0.555 ;
      RECT 3.86 2.215 4.99 2.465 ;
      RECT 4.32 1.455 4.61 1.875 ;
      RECT 4.78 0.085 4.95 0.555 ;
      RECT 4.78 1.455 5.87 1.625 ;
      RECT 4.78 1.625 4.99 2.215 ;
      RECT 5.16 1.795 5.37 2.635 ;
      RECT 5.54 1.625 5.87 2.465 ;
      RECT 5.62 0.085 5.895 0.905 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__nor4bb_2
MACRO sky130_fd_sc_hd__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.115 0.995 3.595 1.275 ;
        RECT 3.295 1.275 3.595 1.705 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 0.995 2.945 1.445 ;
        RECT 2.615 1.445 3.085 1.63 ;
        RECT 2.825 1.63 3.085 2.41 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.24 1.325 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.606900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.955 2.055 2.125 ;
        RECT 1.855 0.655 3.085 0.825 ;
        RECT 1.855 0.825 2.055 1.955 ;
        RECT 2.015 0.3 2.215 0.655 ;
        RECT 2.885 0.31 3.085 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.45 0.405 0.825 ;
      RECT 0.085 0.825 0.26 1.885 ;
      RECT 0.085 1.885 1.205 2.07 ;
      RECT 0.085 2.07 0.345 2.455 ;
      RECT 0.515 2.24 0.845 2.635 ;
      RECT 0.655 0.085 0.825 0.825 ;
      RECT 0.995 1.525 1.59 1.715 ;
      RECT 1.035 2.07 1.205 2.295 ;
      RECT 1.035 2.295 2.395 2.465 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.59 0.825 ;
      RECT 1.41 0.825 1.59 0.995 ;
      RECT 1.41 0.995 1.685 1.325 ;
      RECT 1.41 1.325 1.59 1.525 ;
      RECT 1.515 0.085 1.845 0.48 ;
      RECT 2.225 0.995 2.395 2.295 ;
      RECT 2.385 0.085 2.715 0.485 ;
      RECT 3.255 0.085 3.585 0.825 ;
      RECT 3.255 1.875 3.585 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__nor4bb_1
MACRO sky130_fd_sc_hd__dfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.11 0.795 ;
        RECT 8.855 1.445 9.11 2.325 ;
        RECT 8.9 0.795 9.11 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.04 2.635 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.38 0.085 8.685 0.545 ;
      RECT 8.38 1.495 8.685 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.655 1.785 0.825 1.955 ;
      RECT 1.015 1.105 1.185 1.275 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
    LAYER met1 ;
      RECT 0.595 1.755 0.885 1.8 ;
      RECT 0.595 1.8 6.255 1.94 ;
      RECT 0.595 1.94 0.885 1.985 ;
      RECT 0.955 1.075 1.245 1.12 ;
      RECT 0.955 1.12 6.255 1.26 ;
      RECT 0.955 1.26 1.245 1.305 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtn_1
MACRO sky130_fd_sc_hd__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.66 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 0.105 0.895 0.275 1.46 ;
        RECT 0.105 1.46 3.135 1.63 ;
        RECT 0.605 1.63 0.86 2.435 ;
        RECT 1.03 0.28 1.29 0.725 ;
        RECT 1.465 1.63 1.72 2.435 ;
        RECT 1.89 0.28 2.145 0.725 ;
        RECT 2.32 1.63 2.58 2.435 ;
        RECT 2.835 0.895 3.135 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 1.8 0.43 2.635 ;
      RECT 0.565 0.085 0.86 0.555 ;
      RECT 1.03 1.8 1.29 2.635 ;
      RECT 1.46 0.085 1.72 0.555 ;
      RECT 1.89 1.8 2.15 2.635 ;
      RECT 2.315 0.085 2.615 0.555 ;
      RECT 2.75 1.8 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__clkinv_4
MACRO sky130_fd_sc_hd__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.695 5.44 0.865 ;
        RECT 0.115 0.865 0.285 1.46 ;
        RECT 0.115 1.46 5.44 1.63 ;
        RECT 0.565 1.63 0.805 2.435 ;
        RECT 1.405 1.63 1.645 2.435 ;
        RECT 1.535 0.28 1.725 0.695 ;
        RECT 2.245 1.63 2.495 2.435 ;
        RECT 2.395 0.28 2.585 0.695 ;
        RECT 3.08 1.63 3.325 2.435 ;
        RECT 3.255 0.28 3.445 0.695 ;
        RECT 3.92 1.63 4.175 2.435 ;
        RECT 4.115 0.28 4.305 0.695 ;
        RECT 4.765 1.63 5.005 2.435 ;
        RECT 5.17 0.865 5.44 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.135 1.8 0.395 2.635 ;
      RECT 0.975 1.8 1.235 2.635 ;
      RECT 1.035 0.085 1.365 0.525 ;
      RECT 1.815 1.8 2.075 2.635 ;
      RECT 1.895 0.085 2.225 0.525 ;
      RECT 2.665 1.8 2.91 2.635 ;
      RECT 2.755 0.085 3.085 0.525 ;
      RECT 3.495 1.8 3.75 2.635 ;
      RECT 3.615 0.085 3.945 0.525 ;
      RECT 4.345 1.8 4.595 2.635 ;
      RECT 4.475 0.085 4.805 0.525 ;
      RECT 5.175 1.8 5.43 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__clkinv_8
MACRO sky130_fd_sc_hd__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345 0.895 2.155 1.275 ;
        RECT 8.93 0.895 10.71 1.275 ;
      LAYER mcon ;
        RECT 1.525 1.105 1.695 1.275 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 9.345 1.105 9.515 1.275 ;
        RECT 9.805 1.105 9.975 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 2.215 1.12 ;
        RECT 1.465 1.12 10.035 1.26 ;
        RECT 1.465 1.26 2.215 1.305 ;
        RECT 9.285 1.075 10.035 1.12 ;
        RECT 9.285 1.26 10.035 1.305 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.455 10.48 1.665 ;
        RECT 0.575 1.665 0.83 2.465 ;
        RECT 1.435 1.665 1.69 2.45 ;
        RECT 2.325 0.28 2.55 1.415 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.325 1.665 2.55 2.465 ;
        RECT 3.155 0.28 3.41 1.415 ;
        RECT 3.155 1.665 3.41 2.45 ;
        RECT 4.015 0.28 4.255 1.415 ;
        RECT 4.015 1.665 4.255 2.45 ;
        RECT 4.905 0.28 5.255 1.415 ;
        RECT 4.905 1.665 5.28 2.45 ;
        RECT 5.925 0.28 6.175 1.415 ;
        RECT 5.925 1.665 6.175 2.45 ;
        RECT 6.785 0.28 7.035 1.415 ;
        RECT 6.785 1.665 7.035 2.45 ;
        RECT 7.645 0.28 7.895 1.415 ;
        RECT 7.645 1.665 7.895 2.45 ;
        RECT 8.505 0.28 8.755 1.415 ;
        RECT 8.505 1.665 8.755 2.45 ;
        RECT 9.365 1.665 9.605 2.45 ;
        RECT 10.225 1.665 10.48 2.45 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.14 1.495 0.405 2.635 ;
      RECT 1 1.835 1.26 2.635 ;
      RECT 1.855 0.085 2.125 0.61 ;
      RECT 1.865 1.835 2.12 2.635 ;
      RECT 2.72 0.085 2.985 0.61 ;
      RECT 2.72 1.835 2.98 2.635 ;
      RECT 3.58 0.085 3.845 0.61 ;
      RECT 3.585 1.835 3.84 2.635 ;
      RECT 4.465 0.085 4.73 0.61 ;
      RECT 4.465 1.835 4.72 2.635 ;
      RECT 5.49 0.085 5.755 0.61 ;
      RECT 5.49 1.835 5.745 2.12 ;
      RECT 5.49 2.12 5.75 2.635 ;
      RECT 6.35 0.085 6.575 0.61 ;
      RECT 6.355 1.835 6.61 2.635 ;
      RECT 7.21 0.085 7.475 0.61 ;
      RECT 7.215 1.835 7.47 2.635 ;
      RECT 8.07 0.085 8.335 0.61 ;
      RECT 8.075 1.835 8.33 2.635 ;
      RECT 8.93 0.085 9.195 0.61 ;
      RECT 8.935 1.835 9.19 2.635 ;
      RECT 9.795 1.835 10.05 2.635 ;
      RECT 10.65 1.835 10.91 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
  END
END sky130_fd_sc_hd__clkinv_16
MACRO sky130_fd_sc_hd__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.46 1.755 1.63 ;
        RECT 0.155 1.63 0.41 2.435 ;
        RECT 1.01 1.63 1.27 2.435 ;
        RECT 1.025 0.28 1.25 0.725 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.475 0.895 1.755 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.56 0.085 0.855 0.61 ;
      RECT 0.58 1.8 0.84 2.635 ;
      RECT 1.42 0.085 1.75 0.555 ;
      RECT 1.44 1.8 1.695 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__clkinv_2
MACRO sky130_fd_sc_hd__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.84 0.76 ;
        RECT 0.515 0.76 1.295 1.29 ;
        RECT 0.515 1.29 0.845 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.085 1.665 0.345 2.635 ;
      RECT 1.01 0.085 1.295 0.59 ;
      RECT 1.015 1.665 1.295 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__clkinv_1
MACRO sky130_fd_sc_hd__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 1.065 1.325 1.325 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.725 0.325 1.325 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235 0.255 1.565 0.725 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.655 1.85 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.85 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.33 0.37 0.675 0.545 ;
      RECT 0.415 1.51 1.705 1.68 ;
      RECT 0.415 1.68 0.675 1.905 ;
      RECT 0.495 0.545 0.675 1.51 ;
      RECT 0.855 0.085 1.065 0.895 ;
      RECT 0.875 1.855 1.205 2.635 ;
      RECT 1.535 1.075 1.865 1.245 ;
      RECT 1.535 1.245 1.705 1.51 ;
      RECT 1.735 0.085 2.12 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nor2b_1
MACRO sky130_fd_sc_hd__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.48 1.065 0.92 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.065 3.125 1.275 ;
        RECT 2.91 1.275 3.125 1.965 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 0.895 1.665 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.365 0.895 ;
      RECT 0.085 1.445 1.245 1.655 ;
      RECT 0.085 1.655 0.405 2.465 ;
      RECT 0.575 1.825 0.825 2.635 ;
      RECT 0.995 1.655 1.245 2.295 ;
      RECT 0.995 2.295 2.125 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.835 1.445 2.09 1.89 ;
      RECT 1.835 1.89 2.125 2.295 ;
      RECT 1.875 0.085 2.045 0.895 ;
      RECT 1.875 1.075 2.43 1.245 ;
      RECT 2.215 0.725 2.565 0.895 ;
      RECT 2.215 0.895 2.43 1.075 ;
      RECT 2.26 1.245 2.43 1.445 ;
      RECT 2.26 1.445 2.565 1.615 ;
      RECT 2.395 0.445 2.565 0.725 ;
      RECT 2.395 1.615 2.565 2.46 ;
      RECT 2.775 0.085 3.03 0.845 ;
      RECT 2.775 2.145 3.025 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__nor2b_2
MACRO sky130_fd_sc_hd__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 1.8 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.32 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.085 0.365 0.905 ;
      RECT 0.085 1.455 2.125 1.665 ;
      RECT 0.085 1.665 0.365 2.465 ;
      RECT 0.535 1.835 0.865 2.635 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.375 1.835 1.625 2.635 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.855 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 2.795 1.075 4.275 1.275 ;
      RECT 3.475 1.575 3.855 2.295 ;
      RECT 3.555 0.085 3.845 0.905 ;
      RECT 4.025 0.255 4.355 0.815 ;
      RECT 4.025 0.815 4.275 1.075 ;
      RECT 4.025 1.275 4.275 1.575 ;
      RECT 4.025 1.575 4.355 2.465 ;
      RECT 4.525 0.085 4.815 0.905 ;
      RECT 4.525 1.495 4.93 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__nor2b_4
MACRO sky130_fd_sc_hd__lpflow_inputiso1p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.5 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.765 1.275 1.325 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.18 0.825 ;
        RECT 1.645 1.845 2.18 2.465 ;
        RECT 1.865 0.825 2.18 1.845 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.25 0.085 0.49 0.595 ;
      RECT 0.27 1.495 1.695 1.665 ;
      RECT 0.27 1.665 0.66 1.84 ;
      RECT 0.67 0.265 0.95 0.595 ;
      RECT 0.67 0.595 0.84 1.495 ;
      RECT 1.145 1.835 1.475 2.635 ;
      RECT 1.18 0.085 1.395 0.595 ;
      RECT 1.525 0.995 1.695 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1p_1
MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.765 0.45 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.645 2.2 1.955 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.58 2.68 2.365 ;
        RECT 2.445 0.255 2.68 0.775 ;
        RECT 2.505 0.775 2.68 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.095 0.085 0.425 0.59 ;
      RECT 0.175 1.785 0.855 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.515 2.185 0.845 2.635 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.62 0.655 0.835 0.805 ;
      RECT 0.62 0.805 1.175 1.135 ;
      RECT 0.62 1.135 0.855 1.785 ;
      RECT 1.045 1.305 2.335 1.325 ;
      RECT 1.045 1.325 1.905 1.475 ;
      RECT 1.045 1.475 1.33 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.515 0.61 ;
      RECT 1.345 0.61 1.515 0.945 ;
      RECT 1.345 0.945 2.335 1.305 ;
      RECT 1.51 2.165 2.195 2.635 ;
      RECT 1.875 0.085 2.275 0.58 ;
      RECT 2.865 0.085 3.135 0.72 ;
      RECT 2.865 1.68 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__and2b_2
MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.625 3.155 0.995 ;
        RECT 2.9 0.995 3.205 1.325 ;
        RECT 2.9 1.325 3.155 1.745 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 0.975 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.535 2.73 1.745 ;
        RECT 1.525 0.495 1.715 0.615 ;
        RECT 1.525 0.615 2.73 0.825 ;
        RECT 2.44 0.825 2.73 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.09 0.255 0.425 0.615 ;
      RECT 0.09 0.615 1.355 0.805 ;
      RECT 0.09 2.255 0.425 2.635 ;
      RECT 0.165 0.995 0.425 1.325 ;
      RECT 0.165 1.325 0.335 1.915 ;
      RECT 0.165 1.915 3.505 2.085 ;
      RECT 0.515 1.5 1.315 1.745 ;
      RECT 0.955 0.085 1.285 0.445 ;
      RECT 0.99 2.275 1.32 2.635 ;
      RECT 1.11 1.435 1.32 1.485 ;
      RECT 1.11 1.485 1.315 1.5 ;
      RECT 1.145 0.805 1.355 0.995 ;
      RECT 1.145 0.995 2.26 1.355 ;
      RECT 1.145 1.355 1.32 1.435 ;
      RECT 1.885 0.085 2.215 0.445 ;
      RECT 1.905 2.275 2.235 2.635 ;
      RECT 2.745 0.085 3.075 0.445 ;
      RECT 2.745 2.275 3.075 2.635 ;
      RECT 3.33 0.495 3.5 0.675 ;
      RECT 3.33 0.675 3.545 0.845 ;
      RECT 3.335 1.53 3.545 1.7 ;
      RECT 3.335 1.7 3.505 1.915 ;
      RECT 3.375 0.845 3.545 1.53 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__and2b_4
MACRO sky130_fd_sc_hd__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.645 2.175 1.955 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.58 2.655 2.365 ;
        RECT 2.415 0.255 2.655 0.775 ;
        RECT 2.48 0.775 2.655 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 0.085 0.425 0.59 ;
      RECT 0.175 1.785 0.85 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.515 2.185 0.845 2.635 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.615 0.655 0.835 0.805 ;
      RECT 0.615 0.805 1.15 1.135 ;
      RECT 0.615 1.135 0.85 1.785 ;
      RECT 1.02 1.305 2.305 1.325 ;
      RECT 1.02 1.325 1.88 1.475 ;
      RECT 1.02 1.475 1.305 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.49 0.61 ;
      RECT 1.32 0.61 1.49 0.945 ;
      RECT 1.32 0.945 2.305 1.305 ;
      RECT 1.485 2.165 2.17 2.635 ;
      RECT 1.85 0.085 2.245 0.58 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__and2b_1
MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.39 0.725 3.64 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.655 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.735 1.72 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.97 1.075 1.32 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.909000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.12 1.495 2.67 1.665 ;
        RECT 1.12 1.665 1.45 2.465 ;
        RECT 2.14 1.665 2.47 2.465 ;
        RECT 2.42 0.255 2.93 0.825 ;
        RECT 2.42 0.825 2.67 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.485 0.425 0.715 ;
      RECT 0.085 0.715 1.27 0.905 ;
      RECT 0.085 0.905 0.26 2.065 ;
      RECT 0.085 2.065 0.425 2.465 ;
      RECT 0.595 0.085 0.9 0.545 ;
      RECT 0.595 1.835 0.925 2.635 ;
      RECT 1.08 0.365 2.25 0.555 ;
      RECT 1.08 0.555 1.27 0.715 ;
      RECT 1.64 1.835 1.97 2.635 ;
      RECT 1.97 0.555 2.25 1.325 ;
      RECT 2.68 2.175 3.45 2.635 ;
      RECT 2.84 0.995 3.09 1.835 ;
      RECT 2.84 1.835 4.055 2.005 ;
      RECT 3.1 0.085 3.45 0.545 ;
      RECT 3.62 0.255 4.055 0.545 ;
      RECT 3.635 2.005 4.055 2.465 ;
      RECT 3.81 0.545 4.055 1.835 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__nand4bb_1
MACRO sky130_fd_sc_hd__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.995 0.33 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.995 0.975 1.615 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.12 1.075 7.91 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.42 1.075 10.015 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.655 3.99 0.905 ;
        RECT 2.54 1.445 9.59 1.665 ;
        RECT 2.54 1.665 2.79 2.465 ;
        RECT 3.38 1.665 3.71 2.465 ;
        RECT 3.7 0.905 3.99 1.445 ;
        RECT 4.22 1.665 4.55 2.465 ;
        RECT 5.06 1.665 5.39 2.465 ;
        RECT 6.74 1.665 7.07 2.465 ;
        RECT 7.58 1.665 7.91 2.465 ;
        RECT 8.42 1.665 8.75 2.465 ;
        RECT 9.26 1.665 9.59 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.085 0.255 0.345 0.635 ;
      RECT 0.085 0.635 1.455 0.805 ;
      RECT 0.085 1.785 1.455 1.98 ;
      RECT 0.085 1.98 0.37 2.44 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.54 2.195 0.765 2.635 ;
      RECT 0.935 2.15 1.795 2.465 ;
      RECT 1.015 0.255 1.795 0.465 ;
      RECT 1.145 0.805 1.455 1.785 ;
      RECT 1.625 0.465 1.795 1.075 ;
      RECT 1.625 1.075 2.21 1.305 ;
      RECT 1.625 1.305 1.795 2.15 ;
      RECT 2.2 0.255 5.81 0.485 ;
      RECT 2.2 0.485 2.37 0.905 ;
      RECT 2.2 1.495 2.37 2.635 ;
      RECT 2.54 1.075 3.285 1.245 ;
      RECT 2.96 1.835 3.21 2.635 ;
      RECT 3.88 1.835 4.05 2.635 ;
      RECT 4.16 1.075 5.39 1.275 ;
      RECT 4.22 0.655 5.39 0.735 ;
      RECT 4.22 0.735 6.15 0.905 ;
      RECT 4.72 1.835 4.89 2.635 ;
      RECT 5.61 1.835 6.54 2.635 ;
      RECT 5.98 0.255 7.91 0.485 ;
      RECT 5.98 0.485 6.15 0.735 ;
      RECT 6.32 0.655 10.035 0.905 ;
      RECT 7.24 1.835 7.41 2.635 ;
      RECT 8.08 1.835 8.25 2.635 ;
      RECT 8.42 0.085 8.75 0.485 ;
      RECT 8.92 1.835 9.09 2.635 ;
      RECT 9.26 0.085 9.59 0.485 ;
      RECT 9.76 1.445 10.035 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.98 1.105 2.15 1.275 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.28 1.105 4.45 1.275 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
    LAYER met1 ;
      RECT 1.92 1.075 2.21 1.12 ;
      RECT 1.92 1.12 4.51 1.26 ;
      RECT 1.92 1.26 2.21 1.305 ;
      RECT 4.22 1.075 4.51 1.12 ;
      RECT 4.22 1.26 4.51 1.305 ;
  END
END sky130_fd_sc_hd__nand4bb_4
MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 1.17 0.89 1.34 ;
        RECT 0.61 1.07 0.89 1.17 ;
        RECT 0.61 1.34 0.89 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.07 0.33 1.615 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.72 1.075 4.615 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945 1.075 5.875 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085 0.655 2.415 1.445 ;
        RECT 2.085 1.445 5.455 1.665 ;
        RECT 2.085 1.665 2.335 2.465 ;
        RECT 2.925 1.665 3.255 2.465 ;
        RECT 3.245 1.075 3.55 1.445 ;
        RECT 4.285 1.665 4.615 2.465 ;
        RECT 5.125 1.665 5.455 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.255 0.345 0.73 ;
      RECT 0.085 0.73 1.23 0.9 ;
      RECT 0.085 1.785 1.23 1.98 ;
      RECT 0.085 1.98 0.37 2.44 ;
      RECT 0.515 0.085 0.765 0.545 ;
      RECT 0.54 2.195 0.765 2.635 ;
      RECT 0.935 0.255 1.575 0.56 ;
      RECT 0.935 2.15 1.575 2.465 ;
      RECT 1.06 0.9 1.23 1.785 ;
      RECT 1.4 0.56 1.575 0.715 ;
      RECT 1.4 0.715 1.58 1.41 ;
      RECT 1.4 1.41 1.575 2.15 ;
      RECT 1.745 0.255 3.675 0.485 ;
      RECT 1.745 0.485 1.915 0.585 ;
      RECT 1.745 1.495 1.915 2.635 ;
      RECT 2.505 1.835 2.755 2.635 ;
      RECT 2.745 1.075 3.075 1.275 ;
      RECT 2.925 0.655 4.615 0.905 ;
      RECT 3.425 1.835 4.115 2.635 ;
      RECT 3.865 0.255 5.035 0.485 ;
      RECT 4.785 0.485 5.035 0.735 ;
      RECT 4.785 0.735 5.895 0.905 ;
      RECT 4.785 1.835 4.955 2.635 ;
      RECT 5.205 0.085 5.375 0.565 ;
      RECT 5.545 0.255 5.895 0.735 ;
      RECT 5.625 1.445 5.895 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.06 1.105 1.23 1.275 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 1 1.075 3.135 1.305 ;
  END
END sky130_fd_sc_hd__nand4bb_2
MACRO sky130_fd_sc_hd__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.065 4 1.31 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.05 1.065 2.395 1.48 ;
        RECT 2.05 1.48 5.47 1.705 ;
        RECT 4.225 1.075 5.47 1.48 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.4 1.035 ;
        RECT 0.09 1.035 1.43 1.415 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.58 1.585 1.88 1.705 ;
        RECT 0.58 1.705 1.745 2.035 ;
        RECT 0.595 0.37 0.785 0.615 ;
        RECT 0.595 0.615 1.645 0.695 ;
        RECT 0.595 0.695 3.905 0.865 ;
        RECT 1.455 0.255 1.645 0.615 ;
        RECT 1.6 0.865 3.905 0.895 ;
        RECT 1.6 0.895 1.88 1.585 ;
        RECT 2.275 0.675 3.905 0.695 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.09 0.085 0.425 0.805 ;
      RECT 0.18 1.795 0.375 2.215 ;
      RECT 0.18 2.215 2.115 2.465 ;
      RECT 0.955 0.085 1.285 0.445 ;
      RECT 0.955 2.205 2.115 2.215 ;
      RECT 1.835 0.085 2.115 0.525 ;
      RECT 1.915 1.875 5.625 2.105 ;
      RECT 1.915 2.105 2.115 2.205 ;
      RECT 2.285 0.255 4.335 0.505 ;
      RECT 2.285 2.275 2.615 2.635 ;
      RECT 2.785 2.105 2.975 2.465 ;
      RECT 3.145 2.275 3.475 2.635 ;
      RECT 3.645 2.105 3.835 2.465 ;
      RECT 4.005 2.275 4.335 2.635 ;
      RECT 4.075 0.505 4.335 0.735 ;
      RECT 4.075 0.735 5.195 0.905 ;
      RECT 4.505 0.085 4.695 0.565 ;
      RECT 4.505 2.105 4.685 2.465 ;
      RECT 4.865 0.255 5.195 0.735 ;
      RECT 4.865 2.275 5.195 2.635 ;
      RECT 5.365 0.085 5.625 0.885 ;
      RECT 5.365 2.105 5.625 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__a21oi_4
MACRO sky130_fd_sc_hd__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815 0.995 1.425 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.035 0.645 1.495 ;
        RECT 0.145 1.495 1.93 1.675 ;
        RECT 1.605 1.075 1.935 1.245 ;
        RECT 1.605 1.245 1.93 1.495 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.8 0.995 3.075 1.625 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.255 1.3 0.615 ;
        RECT 0.955 0.615 2.615 0.785 ;
        RECT 2.295 0.255 2.615 0.615 ;
        RECT 2.315 0.785 2.615 2.115 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.1 0.085 0.395 0.865 ;
      RECT 0.11 1.855 2.145 2.025 ;
      RECT 0.11 2.025 1.22 2.105 ;
      RECT 0.11 2.105 0.37 2.465 ;
      RECT 0.54 2.275 0.87 2.635 ;
      RECT 1.05 2.105 1.22 2.465 ;
      RECT 1.475 2.195 1.645 2.635 ;
      RECT 1.76 0.085 2.09 0.445 ;
      RECT 1.815 2.025 2.145 2.285 ;
      RECT 1.815 2.285 3.09 2.465 ;
      RECT 2.785 1.795 3.09 2.285 ;
      RECT 2.795 0.085 3.125 0.825 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a21oi_2
MACRO sky130_fd_sc_hd__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.85 0.995 1.265 1.325 ;
        RECT 1.035 0.375 1.265 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.74 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.675 0.335 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.447000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.68 1.685 ;
        RECT 0.095 1.685 0.37 2.455 ;
        RECT 0.505 0.645 0.835 0.825 ;
        RECT 0.505 0.825 0.68 1.495 ;
        RECT 0.61 0.265 0.835 0.645 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.11 0.085 0.44 0.475 ;
      RECT 0.54 1.855 1.745 2.025 ;
      RECT 0.54 2.025 0.87 2.455 ;
      RECT 0.85 1.525 1.745 1.855 ;
      RECT 1.04 2.195 1.235 2.635 ;
      RECT 1.415 2.025 1.745 2.455 ;
      RECT 1.445 0.085 1.745 0.815 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__a21oi_1
MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235 0.995 3.405 1.445 ;
        RECT 3.235 1.445 3.67 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675 0.995 3.005 1.45 ;
        RECT 2.795 1.45 3.005 1.785 ;
        RECT 2.795 1.785 3.115 2.375 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875 1.455 5.435 1.625 ;
        RECT 3.875 1.625 4.125 2.465 ;
        RECT 3.915 0.255 4.165 0.725 ;
        RECT 3.915 0.725 5.435 0.905 ;
        RECT 4.675 0.255 5.005 0.725 ;
        RECT 4.715 1.625 4.965 2.465 ;
        RECT 5.205 0.905 5.435 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.085 0.45 0.4 0.825 ;
      RECT 0.085 0.825 0.255 1.865 ;
      RECT 0.085 1.865 1.295 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.515 2.205 0.845 2.635 ;
      RECT 0.655 0.085 0.825 0.825 ;
      RECT 0.99 1.525 1.595 1.695 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.595 0.825 ;
      RECT 1.125 2.035 1.295 2.295 ;
      RECT 1.125 2.295 2.445 2.465 ;
      RECT 1.405 0.825 1.595 0.995 ;
      RECT 1.405 0.995 1.695 1.325 ;
      RECT 1.405 1.325 1.595 1.525 ;
      RECT 1.51 1.955 2.105 2.125 ;
      RECT 1.515 0.085 1.845 0.48 ;
      RECT 1.935 0.655 3.745 0.825 ;
      RECT 1.935 0.825 2.105 1.955 ;
      RECT 2.095 0.305 2.265 0.655 ;
      RECT 2.275 0.995 2.445 2.295 ;
      RECT 2.465 0.085 2.795 0.485 ;
      RECT 2.965 0.305 3.135 0.655 ;
      RECT 3.355 0.085 3.735 0.485 ;
      RECT 3.4 1.795 3.65 2.635 ;
      RECT 3.575 0.825 3.745 1.075 ;
      RECT 3.575 1.075 5.035 1.245 ;
      RECT 4.295 1.795 4.545 2.635 ;
      RECT 4.335 0.085 4.505 0.555 ;
      RECT 5.135 1.795 5.385 2.635 ;
      RECT 5.175 0.085 5.345 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__or4bb_4
MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 0.995 3.27 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 2.125 3.12 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 0.415 4.055 0.76 ;
        RECT 3.78 1.495 4.055 2.465 ;
        RECT 3.885 0.76 4.055 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.45 0.4 0.825 ;
      RECT 0.085 0.825 0.255 1.865 ;
      RECT 0.085 1.865 1.915 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.515 2.205 0.845 2.635 ;
      RECT 0.655 0.085 0.825 0.825 ;
      RECT 0.99 1.525 1.575 1.695 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.575 0.825 ;
      RECT 1.405 0.825 1.575 1.075 ;
      RECT 1.405 1.075 1.83 1.245 ;
      RECT 1.405 1.245 1.575 1.525 ;
      RECT 1.47 0.085 1.845 0.485 ;
      RECT 1.51 2.205 2.255 2.375 ;
      RECT 1.745 1.415 2.395 1.585 ;
      RECT 1.745 1.585 1.915 1.865 ;
      RECT 2.015 0.305 2.185 0.655 ;
      RECT 2.015 0.655 3.61 0.825 ;
      RECT 2.085 1.785 3.12 1.955 ;
      RECT 2.085 1.955 2.255 2.205 ;
      RECT 2.225 0.995 2.395 1.415 ;
      RECT 2.37 0.085 2.7 0.485 ;
      RECT 2.87 0.305 3.04 0.655 ;
      RECT 2.95 1.495 3.61 1.665 ;
      RECT 2.95 1.665 3.12 1.785 ;
      RECT 3.21 0.085 3.59 0.485 ;
      RECT 3.29 1.835 3.57 2.635 ;
      RECT 3.44 0.825 3.61 0.995 ;
      RECT 3.44 0.995 3.715 1.325 ;
      RECT 3.44 1.325 3.61 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__or4bb_1
MACRO sky130_fd_sc_hd__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.64 0.995 3.295 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 2.125 3.145 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.24 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.415 4.08 0.76 ;
        RECT 3.805 1.495 4.08 2.465 ;
        RECT 3.91 0.76 4.08 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.45 0.405 0.825 ;
      RECT 0.085 0.825 0.26 1.865 ;
      RECT 0.085 1.865 1.94 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.515 2.205 0.845 2.635 ;
      RECT 0.66 0.085 0.83 0.825 ;
      RECT 0.995 1.525 1.6 1.695 ;
      RECT 1.08 0.45 1.25 0.655 ;
      RECT 1.08 0.655 1.6 0.825 ;
      RECT 1.41 0.825 1.6 1.075 ;
      RECT 1.41 1.075 1.855 1.245 ;
      RECT 1.41 1.245 1.6 1.525 ;
      RECT 1.495 0.085 1.85 0.485 ;
      RECT 1.535 2.205 2.28 2.375 ;
      RECT 1.77 1.415 2.42 1.585 ;
      RECT 1.77 1.585 1.94 1.865 ;
      RECT 2.025 0.305 2.195 0.655 ;
      RECT 2.025 0.655 3.635 0.825 ;
      RECT 2.11 1.785 3.145 1.955 ;
      RECT 2.11 1.955 2.28 2.205 ;
      RECT 2.25 0.995 2.42 1.415 ;
      RECT 2.395 0.085 2.725 0.485 ;
      RECT 2.895 0.305 3.065 0.655 ;
      RECT 2.975 1.495 3.635 1.665 ;
      RECT 2.975 1.665 3.145 1.785 ;
      RECT 3.235 0.085 3.615 0.485 ;
      RECT 3.315 1.835 3.595 2.635 ;
      RECT 3.465 0.825 3.635 0.995 ;
      RECT 3.465 0.995 3.74 1.325 ;
      RECT 3.465 1.325 3.635 1.495 ;
      RECT 4.25 0.085 4.42 1.025 ;
      RECT 4.25 1.44 4.42 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__or4bb_2
MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.735 2.415 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.59 0.085 1.325 0.565 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.335 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.99 1.495 2.235 1.665 ;
      RECT 0.99 1.665 1.41 1.915 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.495 0.655 2.235 0.825 ;
      RECT 1.835 0.085 2.215 0.485 ;
      RECT 1.915 1.835 2.195 2.635 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.295 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1
MACRO sky130_fd_sc_hd__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.325 ;
        RECT 1.46 1.325 1.7 2.405 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.33 0.995 2.675 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.006000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.26 2.675 0.825 ;
        RECT 1.945 0.825 2.16 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.09 1.495 0.44 2.635 ;
      RECT 0.175 0.085 0.345 0.905 ;
      RECT 0.515 0.255 0.845 0.735 ;
      RECT 0.515 0.735 1.7 0.905 ;
      RECT 1.015 0.085 1.185 0.565 ;
      RECT 1.37 0.255 1.7 0.735 ;
      RECT 2.33 1.495 2.675 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__o31ai_1
MACRO sky130_fd_sc_hd__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.055 1.24 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 1.055 2.22 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 1.055 3.205 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.755 4.515 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.063500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.495 4.515 1.665 ;
        RECT 2.335 1.665 2.665 2.125 ;
        RECT 3.175 1.665 3.505 2.465 ;
        RECT 3.675 0.595 4.005 1.495 ;
        RECT 4.175 1.665 4.515 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.09 0.255 0.445 0.715 ;
      RECT 0.09 0.715 3.505 0.885 ;
      RECT 0.09 1.495 2.125 1.665 ;
      RECT 0.09 1.665 0.445 2.465 ;
      RECT 0.615 0.085 0.785 0.545 ;
      RECT 0.615 1.835 0.785 2.635 ;
      RECT 0.955 0.255 1.285 0.715 ;
      RECT 0.955 1.665 1.285 2.465 ;
      RECT 1.455 0.085 1.965 0.545 ;
      RECT 1.455 1.835 1.625 2.295 ;
      RECT 1.455 2.295 3.005 2.465 ;
      RECT 1.795 1.665 2.125 2.125 ;
      RECT 2.175 0.255 2.505 0.715 ;
      RECT 2.675 0.085 3.005 0.545 ;
      RECT 2.835 1.835 3.005 2.295 ;
      RECT 3.175 0.255 4.515 0.425 ;
      RECT 3.175 0.425 3.505 0.715 ;
      RECT 3.675 1.835 4.005 2.635 ;
      RECT 4.175 0.425 4.515 0.585 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__o31ai_2
MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.055 1.78 1.425 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.055 3.605 1.425 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.055 5.94 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.055 7.735 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.683800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.445 7.735 1.695 ;
        RECT 5.77 1.695 5.94 2.465 ;
        RECT 6.11 0.645 7.28 0.885 ;
        RECT 6.11 0.885 6.295 1.445 ;
        RECT 6.61 1.695 6.78 2.465 ;
        RECT 7.45 1.695 7.735 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.09 0.255 0.445 0.715 ;
      RECT 0.09 0.715 5.94 0.885 ;
      RECT 0.09 1.595 2.125 1.895 ;
      RECT 0.09 1.895 0.445 2.465 ;
      RECT 0.615 0.085 0.785 0.545 ;
      RECT 0.615 2.065 0.785 2.635 ;
      RECT 0.955 0.255 1.285 0.715 ;
      RECT 0.955 1.895 1.285 2.465 ;
      RECT 1.455 0.085 1.625 0.545 ;
      RECT 1.455 2.065 1.625 2.635 ;
      RECT 1.795 0.255 2.125 0.715 ;
      RECT 1.795 1.895 2.125 2.205 ;
      RECT 1.795 2.205 3.885 2.465 ;
      RECT 2.295 0.085 2.465 0.545 ;
      RECT 2.295 1.595 3.605 1.765 ;
      RECT 2.295 1.765 2.465 2.035 ;
      RECT 2.635 0.255 2.965 0.715 ;
      RECT 2.635 1.935 2.965 2.205 ;
      RECT 3.135 0.085 3.305 0.545 ;
      RECT 3.135 1.765 3.605 1.865 ;
      RECT 3.135 1.865 5.6 2.035 ;
      RECT 3.475 0.255 3.805 0.715 ;
      RECT 3.995 0.085 4.64 0.545 ;
      RECT 4.08 2.035 5.6 2.465 ;
      RECT 4.81 0.395 4.98 0.715 ;
      RECT 5.15 0.085 5.6 0.545 ;
      RECT 5.77 0.255 7.735 0.475 ;
      RECT 5.77 0.475 5.94 0.715 ;
      RECT 6.11 1.89 6.44 2.635 ;
      RECT 6.95 1.89 7.28 2.635 ;
      RECT 7.45 0.475 7.735 0.885 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__o31ai_4
MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.955 1.785 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 0.415 5.48 0.745 ;
        RECT 5.14 1.67 5.48 2.465 ;
        RECT 5.31 0.745 5.48 1.67 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555 0.255 6.815 0.825 ;
        RECT 6.555 1.505 6.815 2.465 ;
        RECT 6.625 0.825 6.815 1.505 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.48 1.495 2.165 1.665 ;
      RECT 1.48 1.665 1.81 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.165 0.785 ;
      RECT 1.875 0.085 2.23 0.445 ;
      RECT 1.98 1.835 2.295 2.635 ;
      RECT 1.995 0.785 2.165 0.905 ;
      RECT 1.995 0.905 2.365 1.235 ;
      RECT 1.995 1.235 2.165 1.495 ;
      RECT 2.495 1.355 2.78 2.005 ;
      RECT 2.565 0.705 3.12 1.035 ;
      RECT 2.79 0.365 3.525 0.535 ;
      RECT 2.92 2.105 3.62 2.115 ;
      RECT 2.92 2.115 3.615 2.13 ;
      RECT 2.92 2.13 3.61 2.275 ;
      RECT 2.95 1.035 3.12 1.415 ;
      RECT 2.95 1.415 3.29 1.91 ;
      RECT 3.355 0.535 3.525 0.995 ;
      RECT 3.355 0.995 4.225 1.165 ;
      RECT 3.36 2.075 3.63 2.09 ;
      RECT 3.36 2.09 3.625 2.105 ;
      RECT 3.375 2.06 3.63 2.075 ;
      RECT 3.42 2.03 3.63 2.06 ;
      RECT 3.43 2.015 3.63 2.03 ;
      RECT 3.46 1.165 4.225 1.325 ;
      RECT 3.46 1.325 3.63 2.015 ;
      RECT 3.765 0.085 4.095 0.61 ;
      RECT 3.78 2.175 3.95 2.635 ;
      RECT 3.8 1.535 4.58 1.62 ;
      RECT 3.8 1.62 4.55 1.865 ;
      RECT 4.3 0.415 4.47 0.66 ;
      RECT 4.3 0.66 4.58 0.84 ;
      RECT 4.3 1.865 4.55 2.435 ;
      RECT 4.395 0.84 4.58 0.995 ;
      RECT 4.395 0.995 5.14 1.325 ;
      RECT 4.395 1.325 4.58 1.535 ;
      RECT 4.64 0.085 4.97 0.495 ;
      RECT 4.72 1.83 4.97 2.635 ;
      RECT 5.66 0.255 5.91 0.995 ;
      RECT 5.66 0.995 6.455 1.325 ;
      RECT 5.66 1.325 5.91 2.465 ;
      RECT 6.09 0.085 6.385 0.545 ;
      RECT 6.09 1.835 6.385 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.495 1.785 2.665 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.955 1.445 3.125 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.185 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.725 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.435 1.755 2.725 1.8 ;
      RECT 2.435 1.94 2.725 1.985 ;
      RECT 2.895 1.415 3.185 1.46 ;
      RECT 2.895 1.6 3.185 1.645 ;
  END
END sky130_fd_sc_hd__dlxbn_1
MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.955 1.81 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215 0.415 5.465 0.66 ;
        RECT 5.215 0.66 5.5 0.825 ;
        RECT 5.215 1.495 5.5 1.71 ;
        RECT 5.215 1.71 5.465 2.455 ;
        RECT 5.33 0.825 5.5 0.995 ;
        RECT 5.33 0.995 5.905 1.325 ;
        RECT 5.33 1.325 5.5 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.05 0.255 7.305 0.825 ;
        RECT 7.05 1.445 7.305 2.465 ;
        RECT 7.095 0.825 7.305 1.055 ;
        RECT 7.095 1.055 7.735 1.325 ;
        RECT 7.095 1.325 7.305 1.445 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.475 1.495 2.16 1.665 ;
      RECT 1.475 1.665 1.805 2.415 ;
      RECT 1.555 0.345 1.725 0.615 ;
      RECT 1.555 0.615 2.16 0.765 ;
      RECT 1.555 0.765 2.36 0.785 ;
      RECT 1.895 0.085 2.225 0.445 ;
      RECT 1.975 1.835 2.29 2.635 ;
      RECT 1.99 0.785 2.36 1.095 ;
      RECT 1.99 1.095 2.16 1.495 ;
      RECT 2.49 1.355 2.775 2.005 ;
      RECT 2.735 0.705 3.115 1.035 ;
      RECT 2.86 0.365 3.52 0.535 ;
      RECT 2.92 2.255 3.67 2.425 ;
      RECT 2.945 1.035 3.115 1.415 ;
      RECT 2.945 1.415 3.285 1.995 ;
      RECT 3.35 0.535 3.52 0.995 ;
      RECT 3.35 0.995 4.22 1.165 ;
      RECT 3.5 1.165 4.22 1.325 ;
      RECT 3.5 1.325 3.67 2.255 ;
      RECT 3.76 0.085 4.09 0.825 ;
      RECT 3.84 2.135 4.14 2.635 ;
      RECT 3.86 1.535 4.58 1.865 ;
      RECT 4.36 0.415 4.58 0.825 ;
      RECT 4.36 1.865 4.58 2.435 ;
      RECT 4.41 0.825 4.58 0.995 ;
      RECT 4.41 0.995 5.16 1.325 ;
      RECT 4.41 1.325 4.58 1.535 ;
      RECT 4.76 0.085 5.045 0.825 ;
      RECT 4.76 1.495 5.045 2.635 ;
      RECT 5.635 0.085 5.905 0.545 ;
      RECT 5.635 1.835 5.905 2.635 ;
      RECT 6.075 0.255 6.405 0.995 ;
      RECT 6.075 0.995 6.925 1.325 ;
      RECT 6.075 1.325 6.405 2.465 ;
      RECT 6.585 0.085 6.88 0.545 ;
      RECT 6.585 1.835 6.88 2.635 ;
      RECT 7.475 0.085 7.735 0.885 ;
      RECT 7.475 1.495 7.735 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.49 1.785 2.66 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.95 1.445 3.12 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.72 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.43 1.755 2.72 1.8 ;
      RECT 2.43 1.94 2.72 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxbn_2
MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.075 3.645 1.325 ;
        RECT 3.475 1.325 3.645 1.445 ;
        RECT 3.475 1.445 4.965 1.615 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 0.085 1.445 1.685 1.615 ;
        RECT 1.515 1.075 1.895 1.245 ;
        RECT 1.515 1.245 1.685 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 5.235 0.725 6.92 0.905 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.075 0.275 6.405 0.725 ;
        RECT 6.115 1.415 6.92 1.655 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 6.61 0.905 6.92 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.135 1.785 2.065 1.955 ;
      RECT 0.135 1.955 0.385 2.465 ;
      RECT 0.175 0.085 0.345 0.895 ;
      RECT 0.515 0.255 1.685 0.475 ;
      RECT 0.515 0.475 0.765 0.905 ;
      RECT 0.555 2.125 0.805 2.635 ;
      RECT 0.935 0.645 1.27 0.735 ;
      RECT 0.935 0.735 2.525 0.905 ;
      RECT 0.975 1.955 1.225 2.465 ;
      RECT 1.395 2.125 1.645 2.635 ;
      RECT 1.815 1.955 2.065 2.295 ;
      RECT 1.815 2.295 2.905 2.465 ;
      RECT 1.855 0.085 2.025 0.555 ;
      RECT 1.855 1.455 2.065 1.785 ;
      RECT 2.195 0.255 2.525 0.735 ;
      RECT 2.235 0.905 2.445 1.415 ;
      RECT 2.235 1.415 2.62 1.965 ;
      RECT 2.235 1.965 2.485 2.125 ;
      RECT 2.615 1.075 3.145 1.245 ;
      RECT 2.655 2.135 2.905 2.295 ;
      RECT 2.695 0.085 3.385 0.555 ;
      RECT 2.955 0.725 4.725 0.905 ;
      RECT 2.955 0.905 3.145 1.075 ;
      RECT 2.955 1.245 3.145 1.495 ;
      RECT 2.955 1.495 3.305 1.665 ;
      RECT 3.135 1.665 3.305 1.785 ;
      RECT 3.135 1.785 4.265 1.965 ;
      RECT 3.175 2.135 3.425 2.635 ;
      RECT 3.555 0.255 3.885 0.725 ;
      RECT 3.595 2.135 3.845 2.295 ;
      RECT 3.595 2.295 4.685 2.465 ;
      RECT 4.015 1.965 4.265 2.125 ;
      RECT 4.055 0.085 4.225 0.555 ;
      RECT 4.395 0.255 4.725 0.725 ;
      RECT 4.435 1.785 4.685 2.295 ;
      RECT 4.855 1.795 5.105 2.635 ;
      RECT 4.895 0.085 5.065 0.895 ;
      RECT 5.135 1.075 6.44 1.245 ;
      RECT 5.135 1.245 5.46 1.615 ;
      RECT 5.695 2.165 5.945 2.635 ;
      RECT 5.735 0.085 5.905 0.555 ;
      RECT 6.535 1.825 6.785 2.635 ;
      RECT 6.575 0.085 6.745 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.23 1.445 5.4 1.615 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
    LAYER met1 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.46 5.46 1.6 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 5.17 1.415 5.46 1.46 ;
      RECT 5.17 1.6 5.46 1.645 ;
  END
END sky130_fd_sc_hd__a2bb2o_4
MACRO sky130_fd_sc_hd__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.24 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 0.995 1.7 1.375 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.28 0.765 3.54 1.655 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.355 3.08 1.655 ;
        RECT 2.82 0.765 3.08 1.355 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.81 ;
        RECT 0.085 0.81 0.26 1.525 ;
        RECT 0.085 1.525 0.345 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.085 0.945 0.53 ;
      RECT 0.515 1.325 0.685 1.805 ;
      RECT 0.515 1.805 1.275 1.975 ;
      RECT 0.515 2.235 0.845 2.635 ;
      RECT 1.105 1.975 1.275 2.2 ;
      RECT 1.105 2.2 2.245 2.37 ;
      RECT 1.18 0.255 1.35 0.655 ;
      RECT 1.18 0.655 2.06 0.825 ;
      RECT 1.52 0.085 2.24 0.485 ;
      RECT 1.54 1.545 2.06 1.715 ;
      RECT 1.54 1.715 1.71 1.905 ;
      RECT 1.89 0.825 2.06 1.545 ;
      RECT 1.99 1.895 2.4 2.065 ;
      RECT 1.99 2.065 2.245 2.2 ;
      RECT 1.99 2.37 2.245 2.465 ;
      RECT 2.23 0.7 2.58 0.87 ;
      RECT 2.23 0.87 2.4 1.895 ;
      RECT 2.41 0.255 2.58 0.7 ;
      RECT 2.415 2.255 2.745 2.425 ;
      RECT 2.575 1.835 3.515 2.005 ;
      RECT 2.575 2.005 2.745 2.255 ;
      RECT 2.915 2.175 3.165 2.635 ;
      RECT 3.155 0.085 3.555 0.595 ;
      RECT 3.335 2.005 3.515 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a2bb2o_1
MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345 0.995 1.675 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845 0.995 2.135 1.375 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.73 0.765 3.99 1.655 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.355 3.53 1.655 ;
        RECT 3.27 0.765 3.53 1.355 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.255 0.78 0.81 ;
        RECT 0.525 0.81 0.695 1.525 ;
        RECT 0.525 1.525 0.78 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.185 0.085 0.355 0.93 ;
      RECT 0.185 1.445 0.355 2.635 ;
      RECT 0.865 0.995 1.12 1.325 ;
      RECT 0.95 0.085 1.38 0.53 ;
      RECT 0.95 1.325 1.12 1.805 ;
      RECT 0.95 1.805 1.71 1.975 ;
      RECT 0.95 2.235 1.28 2.635 ;
      RECT 1.54 1.975 1.71 2.2 ;
      RECT 1.54 2.2 2.67 2.37 ;
      RECT 1.615 0.255 1.785 0.655 ;
      RECT 1.615 0.655 2.51 0.825 ;
      RECT 1.955 0.085 2.69 0.485 ;
      RECT 1.975 1.545 2.51 1.715 ;
      RECT 1.975 1.715 2.145 1.905 ;
      RECT 2.34 0.825 2.51 1.545 ;
      RECT 2.44 1.895 2.85 2.065 ;
      RECT 2.44 2.065 2.67 2.2 ;
      RECT 2.5 2.37 2.67 2.465 ;
      RECT 2.68 0.7 3.03 0.87 ;
      RECT 2.68 0.87 2.85 1.895 ;
      RECT 2.86 0.255 3.03 0.7 ;
      RECT 2.875 2.255 3.205 2.425 ;
      RECT 3.035 1.835 3.965 2.005 ;
      RECT 3.035 2.005 3.205 2.255 ;
      RECT 3.375 2.175 3.625 2.635 ;
      RECT 3.605 0.085 4.005 0.595 ;
      RECT 3.795 2.005 3.965 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a2bb2o_2
MACRO sky130_fd_sc_hd__lpflow_bleeder_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_bleeder_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN SHORT
    ANTENNAGATEAREA  0.270000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.275 1.04 1.975 1.73 ;
    END
  END SHORT
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.285 0.085 0.615 0.87 ;
      RECT 2.145 0.54 2.475 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__lpflow_bleeder_1
MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.065 1.295 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 4.975 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.155 1.075 6.185 1.295 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.495 1.075 7.505 1.295 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.075 3.145 1.28 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.635 1.605 0.805 ;
        RECT 0.15 0.805 0.32 1.575 ;
        RECT 0.15 1.575 1.605 1.745 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.435 1.745 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 0.095 1.915 0.425 2.635 ;
      RECT 0.49 1.075 1.945 1.245 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 0.935 1.915 1.265 2.635 ;
      RECT 1.775 0.085 2.125 0.465 ;
      RECT 1.775 0.645 3.905 0.815 ;
      RECT 1.775 0.815 1.945 1.075 ;
      RECT 1.775 1.245 1.945 1.455 ;
      RECT 1.775 1.455 2.965 1.625 ;
      RECT 1.775 1.915 2.125 2.635 ;
      RECT 2.295 0.255 2.465 0.645 ;
      RECT 2.375 1.795 2.545 2.295 ;
      RECT 2.375 2.295 3.405 2.465 ;
      RECT 2.635 0.085 2.965 0.465 ;
      RECT 2.715 1.955 3.045 2.125 ;
      RECT 2.795 1.625 2.965 1.955 ;
      RECT 3.155 0.295 4.245 0.465 ;
      RECT 3.235 1.535 7.37 1.705 ;
      RECT 3.235 1.705 3.405 2.295 ;
      RECT 3.575 1.915 3.905 2.635 ;
      RECT 4.075 0.465 4.245 0.645 ;
      RECT 4.075 0.645 5.165 0.815 ;
      RECT 4.075 1.705 4.245 2.465 ;
      RECT 4.415 0.295 6.105 0.465 ;
      RECT 4.415 1.915 4.745 2.635 ;
      RECT 4.935 1.705 5.105 2.465 ;
      RECT 5.345 1.915 6.035 2.635 ;
      RECT 5.355 0.645 7.285 0.815 ;
      RECT 6.275 1.705 6.445 2.465 ;
      RECT 6.615 0.085 6.945 0.465 ;
      RECT 6.615 1.915 6.945 2.635 ;
      RECT 7.115 0.255 7.285 0.645 ;
      RECT 7.115 1.705 7.285 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__a41o_4
MACRO sky130_fd_sc_hd__a41o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785 0.73 4.005 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085 1.075 3.55 1.245 ;
        RECT 3.335 0.745 3.55 1.075 ;
        RECT 3.335 1.245 3.55 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.995 2.855 1.435 ;
        RECT 2.685 1.435 3.09 1.625 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2 0.995 2.335 1.625 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.4 1.075 1.73 1.295 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.295 0.765 0.755 ;
        RECT 0.595 0.755 0.785 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.095 0.085 0.425 0.805 ;
      RECT 0.095 1.495 0.425 2.635 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 0.98 0.635 2.545 0.805 ;
      RECT 0.98 0.805 1.15 1.495 ;
      RECT 0.98 1.495 1.785 1.665 ;
      RECT 1.015 1.835 1.265 2.635 ;
      RECT 1.455 1.665 1.785 2.425 ;
      RECT 1.495 0.255 1.705 0.635 ;
      RECT 1.875 0.085 2.205 0.465 ;
      RECT 1.955 1.795 3.965 1.965 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.335 2.175 2.585 2.635 ;
      RECT 2.375 0.295 4.045 0.465 ;
      RECT 2.375 0.465 2.545 0.635 ;
      RECT 2.795 1.965 2.965 2.465 ;
      RECT 3.335 2.175 3.585 2.635 ;
      RECT 3.795 1.965 3.965 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a41o_2
MACRO sky130_fd_sc_hd__a41o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 0.995 1.915 1.325 ;
        RECT 1.535 1.325 1.835 1.62 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.7 0.415 2.65 0.6 ;
        RECT 2.225 0.6 2.445 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705 0.995 3.085 1.625 ;
        RECT 2.88 0.395 3.085 0.995 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 0.995 3.57 1.625 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.635 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.3 0.425 0.56 ;
        RECT 0.085 0.56 0.345 2.165 ;
        RECT 0.085 2.165 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.515 0.735 1.53 0.81 ;
      RECT 0.515 0.81 1.335 0.905 ;
      RECT 0.515 0.905 0.685 1.825 ;
      RECT 0.515 1.825 1.365 1.995 ;
      RECT 0.595 0.085 0.925 0.565 ;
      RECT 0.595 2.175 0.845 2.635 ;
      RECT 1.035 1.995 1.365 2.425 ;
      RECT 1.115 0.3 1.53 0.735 ;
      RECT 1.535 1.795 3.505 1.965 ;
      RECT 1.535 1.965 1.705 2.465 ;
      RECT 1.915 2.175 2.165 2.635 ;
      RECT 2.375 1.965 2.545 2.465 ;
      RECT 2.845 2.175 3.095 2.635 ;
      RECT 3.255 0.085 3.595 0.81 ;
      RECT 3.335 1.965 3.505 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a41o_1
MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645 0.995 7.8 1.285 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.87 0.62 8.195 0.825 ;
        RECT 4.87 1.455 8.195 1.625 ;
        RECT 4.87 1.625 5.2 2.125 ;
        RECT 5.71 1.625 6.04 2.125 ;
        RECT 6.55 1.625 6.88 2.125 ;
        RECT 7.39 1.625 7.72 2.125 ;
        RECT 7.97 0.825 8.195 1.455 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.09 0.255 0.345 0.655 ;
      RECT 0.09 0.655 0.845 0.825 ;
      RECT 0.09 1.495 0.845 1.665 ;
      RECT 0.09 1.665 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 0.825 0.845 0.995 ;
      RECT 0.515 0.995 4.475 1.325 ;
      RECT 0.515 1.325 0.845 1.495 ;
      RECT 0.515 1.835 0.845 2.635 ;
      RECT 1.015 0.255 1.285 0.655 ;
      RECT 1.015 0.655 4.7 0.825 ;
      RECT 1.015 1.495 4.7 1.665 ;
      RECT 1.015 1.665 1.24 2.465 ;
      RECT 1.41 1.835 1.74 2.635 ;
      RECT 1.455 0.085 1.785 0.485 ;
      RECT 1.91 1.665 2.08 2.465 ;
      RECT 1.955 0.255 2.125 0.655 ;
      RECT 2.25 1.835 2.58 2.635 ;
      RECT 2.295 0.085 2.625 0.485 ;
      RECT 2.75 1.665 2.92 2.465 ;
      RECT 2.795 0.255 2.965 0.655 ;
      RECT 3.09 1.835 3.42 2.635 ;
      RECT 3.135 0.085 3.465 0.485 ;
      RECT 3.59 1.665 3.76 2.465 ;
      RECT 3.635 0.255 3.805 0.655 ;
      RECT 3.93 1.835 4.28 2.635 ;
      RECT 3.975 0.085 4.315 0.485 ;
      RECT 4.45 1.665 4.7 2.295 ;
      RECT 4.45 2.295 8.195 2.465 ;
      RECT 4.485 0.255 8.195 0.45 ;
      RECT 4.485 0.45 4.7 0.655 ;
      RECT 5.37 1.795 5.54 2.295 ;
      RECT 6.21 1.795 6.38 2.295 ;
      RECT 7.05 1.795 7.22 2.295 ;
      RECT 7.89 1.795 8.195 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
  END
END sky130_fd_sc_hd__einvn_8
MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.765 1.755 1.955 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.65 1.725 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.275600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.16 0.255 1.755 0.595 ;
        RECT 1.16 0.595 1.33 2.125 ;
        RECT 1.16 2.125 1.755 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.085 0.255 0.36 0.655 ;
      RECT 0.085 0.655 0.99 0.825 ;
      RECT 0.085 1.895 0.99 2.065 ;
      RECT 0.085 2.065 0.4 2.465 ;
      RECT 0.53 0.085 0.99 0.485 ;
      RECT 0.57 2.235 0.99 2.635 ;
      RECT 0.82 0.825 0.99 1.895 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__einvn_0
MACRO sky130_fd_sc_hd__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.275 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.325 1.385 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.694800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.445 3.135 1.695 ;
        RECT 2.365 0.595 2.695 0.845 ;
        RECT 2.365 0.845 2.615 1.445 ;
        RECT 2.785 1.695 3.135 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.84 0.825 ;
      RECT 0.085 1.555 0.895 1.725 ;
      RECT 0.085 1.725 0.345 2.465 ;
      RECT 0.495 0.825 0.84 0.995 ;
      RECT 0.495 0.995 2.035 1.275 ;
      RECT 0.495 1.275 0.895 1.555 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 1.895 0.895 2.635 ;
      RECT 1.015 0.255 1.28 0.655 ;
      RECT 1.015 0.655 2.195 0.825 ;
      RECT 1.07 1.445 1.775 1.865 ;
      RECT 1.07 1.865 2.615 2.085 ;
      RECT 1.07 2.085 1.24 2.465 ;
      RECT 1.41 2.255 2.275 2.635 ;
      RECT 1.45 0.085 1.78 0.485 ;
      RECT 1.95 0.255 3.135 0.425 ;
      RECT 1.95 0.425 2.195 0.655 ;
      RECT 2.445 2.085 2.615 2.465 ;
      RECT 2.865 0.425 3.135 0.775 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__einvn_2
MACRO sky130_fd_sc_hd__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.53 0.62 4.975 1.325 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.62 4.36 1.48 ;
        RECT 3.19 1.48 3.52 2.075 ;
        RECT 4.03 1.48 4.36 2.075 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.845 0.825 ;
      RECT 0.085 1.495 0.845 1.665 ;
      RECT 0.085 1.665 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 0.825 0.845 0.995 ;
      RECT 0.515 0.995 3.02 1.325 ;
      RECT 0.515 1.325 0.845 1.495 ;
      RECT 0.515 1.835 0.845 2.635 ;
      RECT 1.015 0.255 1.285 0.655 ;
      RECT 1.015 0.655 2.995 0.825 ;
      RECT 1.015 1.495 3.02 1.665 ;
      RECT 1.015 1.665 1.24 2.465 ;
      RECT 1.41 1.835 1.74 2.635 ;
      RECT 1.455 0.085 1.785 0.485 ;
      RECT 1.91 1.665 2.08 2.465 ;
      RECT 1.955 0.255 2.125 0.655 ;
      RECT 2.25 1.835 2.64 2.635 ;
      RECT 2.295 0.085 2.625 0.485 ;
      RECT 2.81 1.665 3.02 2.295 ;
      RECT 2.81 2.295 4.975 2.465 ;
      RECT 2.825 0.255 4.975 0.45 ;
      RECT 2.825 0.45 2.995 0.655 ;
      RECT 3.69 1.65 3.86 2.295 ;
      RECT 4.53 1.65 4.975 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__einvn_4
MACRO sky130_fd_sc_hd__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.765 2.215 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.51 1.725 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 1.785 2.215 2.465 ;
        RECT 1.62 0.255 2.215 0.595 ;
        RECT 1.62 0.595 1.8 1.785 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.255 0.37 0.615 ;
      RECT 0.085 0.615 1.45 0.785 ;
      RECT 0.085 1.895 0.87 2.065 ;
      RECT 0.085 2.065 0.37 2.465 ;
      RECT 0.54 0.085 1.44 0.445 ;
      RECT 0.54 2.235 0.87 2.635 ;
      RECT 0.685 0.785 1.45 1.615 ;
      RECT 0.685 1.615 0.87 1.895 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__einvn_1
MACRO sky130_fd_sc_hd__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.955 1.81 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215 0.415 5.465 0.685 ;
        RECT 5.215 0.685 5.5 0.825 ;
        RECT 5.215 1.495 5.5 1.64 ;
        RECT 5.215 1.64 5.465 2.455 ;
        RECT 5.33 0.825 5.5 0.995 ;
        RECT 5.33 0.995 5.895 1.325 ;
        RECT 5.33 1.325 5.5 1.495 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.475 1.495 2.16 1.665 ;
      RECT 1.475 1.665 1.805 2.415 ;
      RECT 1.555 0.345 1.725 0.615 ;
      RECT 1.555 0.615 2.16 0.765 ;
      RECT 1.555 0.765 2.36 0.785 ;
      RECT 1.895 0.085 2.225 0.445 ;
      RECT 1.975 1.835 2.29 2.635 ;
      RECT 1.99 0.785 2.36 1.095 ;
      RECT 1.99 1.095 2.16 1.495 ;
      RECT 2.49 1.355 2.775 2.005 ;
      RECT 2.735 0.705 3.115 1.035 ;
      RECT 2.86 0.365 3.52 0.535 ;
      RECT 2.92 2.255 3.67 2.425 ;
      RECT 2.945 1.035 3.115 1.415 ;
      RECT 2.945 1.415 3.285 1.995 ;
      RECT 3.35 0.535 3.52 0.995 ;
      RECT 3.35 0.995 4.22 1.165 ;
      RECT 3.5 1.165 4.22 1.325 ;
      RECT 3.5 1.325 3.67 2.255 ;
      RECT 3.76 0.085 4.09 0.825 ;
      RECT 3.84 2.135 4.14 2.635 ;
      RECT 3.86 1.535 4.58 1.865 ;
      RECT 4.36 0.415 4.58 0.825 ;
      RECT 4.36 1.865 4.58 2.435 ;
      RECT 4.41 0.825 4.58 0.995 ;
      RECT 4.41 0.995 5.16 1.325 ;
      RECT 4.41 1.325 4.58 1.535 ;
      RECT 4.76 0.085 5.045 0.825 ;
      RECT 4.76 1.495 5.045 2.635 ;
      RECT 5.635 0.085 5.895 0.55 ;
      RECT 5.635 1.755 5.895 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.49 1.785 2.66 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.95 1.445 3.12 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.72 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.43 1.755 2.72 1.8 ;
      RECT 2.43 1.94 2.72 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_2
MACRO sky130_fd_sc_hd__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.175 0.415 5.435 0.745 ;
        RECT 5.175 1.67 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.67 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.785 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.115 0.765 ;
      RECT 1.51 0.765 2.32 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.945 0.785 2.32 1.235 ;
      RECT 1.945 1.235 2.115 1.495 ;
      RECT 1.955 1.835 2.245 2.635 ;
      RECT 2.445 1.355 2.78 2.005 ;
      RECT 2.56 0.735 3.265 1.04 ;
      RECT 2.745 2.255 3.605 2.425 ;
      RECT 2.765 0.365 3.605 0.535 ;
      RECT 2.95 1.04 3.265 1.56 ;
      RECT 2.95 1.56 3.285 1.91 ;
      RECT 3.295 2.09 3.62 2.105 ;
      RECT 3.295 2.105 3.605 2.255 ;
      RECT 3.39 2.045 3.645 2.065 ;
      RECT 3.39 2.065 3.63 2.085 ;
      RECT 3.39 2.085 3.62 2.09 ;
      RECT 3.405 2.035 3.645 2.045 ;
      RECT 3.43 2.01 3.645 2.035 ;
      RECT 3.435 0.535 3.605 0.995 ;
      RECT 3.435 0.995 4.2 1.325 ;
      RECT 3.435 1.325 3.645 1.45 ;
      RECT 3.455 1.45 3.645 2.01 ;
      RECT 3.775 0.085 4.045 0.545 ;
      RECT 3.775 2.175 4.095 2.635 ;
      RECT 3.815 1.535 4.54 1.865 ;
      RECT 4.295 0.26 4.54 0.72 ;
      RECT 4.295 1.865 4.54 2.435 ;
      RECT 4.37 0.72 4.54 0.995 ;
      RECT 4.37 0.995 5.095 1.325 ;
      RECT 4.37 1.325 4.54 1.535 ;
      RECT 4.72 1.57 5.005 2.635 ;
      RECT 4.755 0.085 4.98 0.715 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.95 1.445 3.12 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.675 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_1
MACRO sky130_fd_sc_hd__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.24 0.415 5.525 0.745 ;
        RECT 5.24 1.495 5.525 2.455 ;
        RECT 5.355 0.745 5.525 0.995 ;
        RECT 5.355 0.995 6.815 1.325 ;
        RECT 5.355 1.325 5.525 1.495 ;
        RECT 6.115 0.385 6.385 0.995 ;
        RECT 6.115 1.325 6.385 2.455 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.48 1.165 4.2 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.74 0.085 4.07 0.53 ;
      RECT 3.82 2.135 4.12 2.635 ;
      RECT 3.84 1.535 4.605 1.865 ;
      RECT 4.385 0.415 4.605 0.745 ;
      RECT 4.385 1.865 4.605 2.435 ;
      RECT 4.435 0.745 4.605 0.995 ;
      RECT 4.435 0.995 5.185 1.325 ;
      RECT 4.435 1.325 4.605 1.535 ;
      RECT 4.785 0.085 5.07 0.715 ;
      RECT 4.785 1.495 5.07 2.635 ;
      RECT 5.695 0.085 5.945 0.825 ;
      RECT 5.695 1.495 5.945 2.635 ;
      RECT 6.555 0.085 6.815 0.715 ;
      RECT 6.555 1.495 6.815 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_4
MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s6s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.575 1.7 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.08 0.255 4.515 0.825 ;
        RECT 4.08 1.495 4.515 2.465 ;
        RECT 4.155 0.825 4.515 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.255 0.525 0.655 ;
      RECT 0.085 0.655 1.08 0.825 ;
      RECT 0.085 1.87 1.08 2.04 ;
      RECT 0.085 2.04 0.525 2.465 ;
      RECT 0.695 0.085 1.08 0.485 ;
      RECT 0.695 2.21 1.08 2.635 ;
      RECT 0.745 0.825 1.08 0.995 ;
      RECT 0.745 0.995 1.155 1.325 ;
      RECT 0.745 1.325 1.08 1.87 ;
      RECT 1.25 0.255 1.52 0.825 ;
      RECT 1.25 1.495 1.975 1.675 ;
      RECT 1.25 1.675 1.52 2.465 ;
      RECT 1.325 0.825 1.52 0.995 ;
      RECT 1.325 0.995 1.975 1.495 ;
      RECT 1.69 0.255 1.94 0.655 ;
      RECT 1.69 0.655 2.495 0.825 ;
      RECT 1.69 1.845 2.495 2.04 ;
      RECT 1.69 2.04 1.94 2.465 ;
      RECT 2.11 0.085 2.495 0.485 ;
      RECT 2.11 2.21 2.495 2.635 ;
      RECT 2.145 0.825 2.495 0.995 ;
      RECT 2.145 0.995 2.57 1.325 ;
      RECT 2.145 1.325 2.495 1.845 ;
      RECT 2.665 0.255 2.915 0.825 ;
      RECT 2.665 1.495 3.39 1.675 ;
      RECT 2.665 1.675 2.915 2.465 ;
      RECT 2.74 0.825 2.915 0.995 ;
      RECT 2.74 0.995 3.39 1.495 ;
      RECT 3.085 0.255 3.355 0.655 ;
      RECT 3.085 0.655 3.91 0.825 ;
      RECT 3.085 1.845 3.91 2.04 ;
      RECT 3.085 2.04 3.355 2.465 ;
      RECT 3.525 0.085 3.91 0.485 ;
      RECT 3.525 2.21 3.91 2.635 ;
      RECT 3.56 0.825 3.91 0.995 ;
      RECT 3.56 0.995 3.985 1.325 ;
      RECT 3.56 1.325 3.91 1.845 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1
MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 6.885 1.575 7.215 2.42 ;
        RECT 6.895 0.305 7.225 0.74 ;
        RECT 6.895 0.74 7.275 0.825 ;
        RECT 7.05 0.825 7.275 0.865 ;
        RECT 7.06 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.44 2.175 1.705 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.4 0.085 3.77 0.585 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.61 1.835 3.78 2.635 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.015 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.375 1.905 ;
      RECT 5.49 2.135 5.805 2.635 ;
      RECT 5.585 0.085 5.795 0.615 ;
      RECT 6.035 1.905 6.375 2.465 ;
      RECT 6.055 0.3 6.385 0.825 ;
      RECT 6.185 0.825 6.385 0.995 ;
      RECT 6.185 0.995 6.935 1.325 ;
      RECT 6.185 1.325 6.375 1.53 ;
      RECT 6.545 1.625 6.715 2.635 ;
      RECT 6.555 0.085 6.725 0.695 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxtp_1
MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.065 1.72 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985 0.305 7.32 0.73 ;
        RECT 6.985 0.73 8.655 0.9 ;
        RECT 6.985 1.465 8.655 1.635 ;
        RECT 6.985 1.635 7.32 2.395 ;
        RECT 7.84 0.305 8.175 0.73 ;
        RECT 7.84 1.635 8.17 2.395 ;
        RECT 8.41 0.9 8.655 1.465 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.44 2.175 1.705 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.89 0.365 2.22 0.535 ;
      RECT 1.89 0.535 2.06 2.065 ;
      RECT 1.89 2.065 2.125 2.44 ;
      RECT 2.23 0.705 2.81 1.035 ;
      RECT 2.23 1.035 2.47 1.905 ;
      RECT 2.37 2.19 3.44 2.36 ;
      RECT 2.4 0.365 3.15 0.535 ;
      RECT 2.66 1.655 3.1 2.01 ;
      RECT 2.98 0.535 3.15 1.315 ;
      RECT 2.98 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.32 0.765 4.12 1.065 ;
      RECT 3.32 1.065 3.49 1.095 ;
      RECT 3.4 0.085 3.77 0.585 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.61 1.835 3.78 2.635 ;
      RECT 3.95 0.365 4.41 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 0.705 4.84 1.035 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.64 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.84 1.575 ;
      RECT 4.65 1.575 4.97 1.905 ;
      RECT 5.14 0.535 5.31 1.075 ;
      RECT 5.14 1.075 6.23 1.245 ;
      RECT 5.14 1.245 5.31 2.165 ;
      RECT 5.48 1.5 6.59 1.67 ;
      RECT 5.48 1.67 6.34 1.83 ;
      RECT 5.49 2.135 5.705 2.635 ;
      RECT 5.625 0.085 5.795 0.615 ;
      RECT 6.09 0.295 6.45 0.735 ;
      RECT 6.09 0.735 6.59 0.905 ;
      RECT 6.17 1.83 6.34 2.455 ;
      RECT 6.42 0.905 6.59 1.075 ;
      RECT 6.42 1.075 8.24 1.245 ;
      RECT 6.42 1.245 6.59 1.5 ;
      RECT 6.625 0.085 6.795 0.565 ;
      RECT 6.625 1.855 6.805 2.635 ;
      RECT 7.495 0.085 7.665 0.56 ;
      RECT 7.5 1.805 7.67 2.635 ;
      RECT 8.34 1.805 8.51 2.635 ;
      RECT 8.345 0.085 8.515 0.56 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 0.765 2.64 0.935 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.785 3.1 1.955 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.31 0.765 4.48 0.935 ;
      RECT 4.31 1.785 4.48 1.955 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 4.54 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 4.54 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.41 0.735 2.7 0.78 ;
      RECT 2.41 0.92 2.7 0.965 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
      RECT 4.25 0.735 4.54 0.78 ;
      RECT 4.25 0.92 4.54 0.965 ;
      RECT 4.25 1.755 4.54 1.8 ;
      RECT 4.25 1.94 4.54 1.985 ;
  END
END sky130_fd_sc_hd__dfxtp_4
MACRO sky130_fd_sc_hd__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 6.885 1.575 7.215 2.42 ;
        RECT 6.895 0.305 7.225 0.74 ;
        RECT 6.895 0.74 7.275 0.825 ;
        RECT 7.05 0.825 7.275 0.865 ;
        RECT 7.06 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.44 2.175 1.705 2.635 ;
      RECT 1.455 0.085 1.705 0.545 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.4 0.085 3.77 0.585 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.61 1.835 3.78 2.635 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.015 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.375 1.905 ;
      RECT 5.49 2.135 5.805 2.635 ;
      RECT 5.585 0.085 5.795 0.615 ;
      RECT 6.035 1.905 6.375 2.465 ;
      RECT 6.055 0.3 6.385 0.825 ;
      RECT 6.185 0.825 6.385 0.995 ;
      RECT 6.185 0.995 6.935 1.325 ;
      RECT 6.185 1.325 6.375 1.53 ;
      RECT 6.545 1.625 6.715 2.635 ;
      RECT 6.555 0.085 6.725 0.695 ;
      RECT 7.385 1.72 7.555 2.635 ;
      RECT 7.395 0.085 7.565 0.6 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxtp_2
MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.995 5.42 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.55 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.67 0.995 6.855 1.63 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.443500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.635 7.585 0.805 ;
        RECT 6.075 1.915 7.245 2.085 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.045 0.805 7.245 1.915 ;
        RECT 7.415 0.255 7.585 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 3.785 0.805 ;
      RECT 0.175 1.495 5.405 1.665 ;
      RECT 0.175 1.665 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 1.915 0.845 2.635 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.015 1.665 1.185 2.465 ;
      RECT 1.355 0.085 1.685 0.465 ;
      RECT 1.355 1.915 1.685 2.635 ;
      RECT 1.855 0.255 2.025 0.635 ;
      RECT 1.855 1.665 2.025 2.465 ;
      RECT 2.195 0.295 5.565 0.465 ;
      RECT 2.195 1.915 2.525 2.635 ;
      RECT 2.695 1.665 2.865 2.465 ;
      RECT 3.035 1.915 3.365 2.635 ;
      RECT 3.535 1.665 3.705 2.465 ;
      RECT 3.895 1.915 4.225 2.635 ;
      RECT 4.395 1.665 4.565 2.465 ;
      RECT 4.735 2.255 5.065 2.635 ;
      RECT 5.235 1.665 5.405 2.255 ;
      RECT 5.235 2.255 7.665 2.425 ;
      RECT 5.235 2.425 5.405 2.465 ;
      RECT 6.075 0.085 6.405 0.465 ;
      RECT 6.915 0.085 7.245 0.465 ;
      RECT 7.415 1.495 7.665 2.255 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__a31oi_4
MACRO sky130_fd_sc_hd__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.665 1.615 ;
        RECT 2.905 0.995 3.075 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.995 1.755 1.615 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.82 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.82 1.075 4.49 1.275 ;
        RECT 4.265 1.275 4.49 1.625 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.922000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295 0.655 4.505 0.825 ;
        RECT 3.255 0.255 3.425 0.655 ;
        RECT 3.255 0.825 3.57 1.445 ;
        RECT 3.255 1.445 4.085 1.615 ;
        RECT 3.755 1.615 4.085 2.115 ;
        RECT 4.175 0.295 4.505 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.095 0.655 2.105 0.825 ;
      RECT 0.175 1.785 3.505 1.955 ;
      RECT 0.175 1.955 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.125 0.845 2.635 ;
      RECT 1.015 1.955 1.185 2.465 ;
      RECT 1.355 0.295 3.075 0.465 ;
      RECT 1.355 2.125 1.685 2.635 ;
      RECT 1.855 1.955 2.025 2.465 ;
      RECT 2.31 2.125 2.98 2.635 ;
      RECT 3.335 1.955 3.505 2.295 ;
      RECT 3.335 2.295 4.425 2.465 ;
      RECT 3.675 0.085 4.005 0.465 ;
      RECT 4.255 1.795 4.425 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__a31oi_2
MACRO sky130_fd_sc_hd__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.445 1.455 1.665 ;
        RECT 1.27 0.995 1.455 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.335 1.055 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.365 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.215 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.38 0.295 1.785 0.715 ;
        RECT 1.38 0.715 1.795 0.825 ;
        RECT 1.625 0.825 1.795 1.495 ;
        RECT 1.625 1.495 2.21 1.665 ;
        RECT 1.875 1.665 2.21 2.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.09 0.085 0.43 0.815 ;
      RECT 0.09 1.495 0.42 2.635 ;
      RECT 0.59 1.835 1.695 2.005 ;
      RECT 0.59 2.005 0.765 2.415 ;
      RECT 0.935 2.175 1.265 2.635 ;
      RECT 1.47 2.005 1.695 2.415 ;
      RECT 1.955 0.085 2.215 0.565 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__a31oi_1
MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685 0.995 6.855 1.445 ;
        RECT 6.685 1.445 7.265 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.86 0.995 2.495 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.59 0.925 ;
        RECT 0.085 0.925 0.4 1.44 ;
        RECT 0.085 1.44 0.61 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.93 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 0.75 0.995 0.95 1.325 ;
      RECT 0.76 0.085 1.01 0.525 ;
      RECT 0.78 0.695 1.35 0.865 ;
      RECT 0.78 0.865 0.95 0.995 ;
      RECT 0.78 1.325 0.95 1.875 ;
      RECT 0.78 1.875 1.47 2.045 ;
      RECT 0.78 2.215 1.115 2.635 ;
      RECT 1.18 0.255 2.74 0.425 ;
      RECT 1.18 0.425 1.35 0.695 ;
      RECT 1.185 1.535 2.835 1.705 ;
      RECT 1.3 2.045 1.47 2.235 ;
      RECT 1.3 2.235 2.895 2.405 ;
      RECT 1.52 0.595 1.69 1.535 ;
      RECT 1.87 1.895 3.175 2.065 ;
      RECT 1.97 0.655 3.08 0.825 ;
      RECT 2.39 0.425 2.74 0.455 ;
      RECT 2.665 0.995 2.94 1.325 ;
      RECT 2.665 1.325 2.835 1.535 ;
      RECT 2.91 0.255 3.76 0.425 ;
      RECT 2.91 0.425 3.08 0.655 ;
      RECT 3.005 1.525 3.535 1.695 ;
      RECT 3.005 1.695 3.175 1.895 ;
      RECT 3.11 2.235 3.515 2.405 ;
      RECT 3.25 0.595 3.42 1.375 ;
      RECT 3.25 1.375 3.535 1.525 ;
      RECT 3.345 1.895 4.52 2.065 ;
      RECT 3.345 2.065 3.515 2.235 ;
      RECT 3.59 0.425 3.76 1.035 ;
      RECT 3.59 1.035 3.875 1.205 ;
      RECT 3.685 2.235 4.015 2.635 ;
      RECT 3.705 1.205 3.875 1.895 ;
      RECT 3.93 0.085 4.1 0.865 ;
      RECT 4.105 1.445 4.52 1.715 ;
      RECT 4.28 0.415 4.52 1.445 ;
      RECT 4.35 2.065 4.52 2.275 ;
      RECT 4.35 2.275 7.445 2.445 ;
      RECT 4.695 0.265 5.11 0.485 ;
      RECT 4.695 0.485 4.915 0.595 ;
      RECT 4.695 0.595 4.865 2.105 ;
      RECT 5.035 0.72 5.45 0.825 ;
      RECT 5.035 0.825 5.255 0.89 ;
      RECT 5.035 0.89 5.205 2.275 ;
      RECT 5.085 0.655 5.45 0.72 ;
      RECT 5.28 0.32 5.45 0.655 ;
      RECT 5.395 1.445 6.175 1.615 ;
      RECT 5.395 1.615 5.81 2.045 ;
      RECT 5.41 0.995 5.835 1.27 ;
      RECT 5.62 0.63 5.835 0.995 ;
      RECT 6.005 0.255 7.15 0.425 ;
      RECT 6.005 0.425 6.175 1.445 ;
      RECT 6.345 0.595 6.515 1.935 ;
      RECT 6.345 1.935 8.655 2.105 ;
      RECT 6.685 0.425 7.15 0.465 ;
      RECT 7.025 0.73 7.23 0.945 ;
      RECT 7.025 0.945 7.335 1.275 ;
      RECT 7.435 1.495 8.255 1.705 ;
      RECT 7.475 0.295 7.765 0.735 ;
      RECT 7.475 0.735 8.255 0.75 ;
      RECT 7.515 0.75 8.255 0.905 ;
      RECT 7.855 2.275 8.19 2.635 ;
      RECT 7.935 0.085 8.105 0.565 ;
      RECT 8.085 0.905 8.255 0.995 ;
      RECT 8.085 0.995 8.315 1.325 ;
      RECT 8.085 1.325 8.255 1.495 ;
      RECT 8.17 1.875 8.655 1.935 ;
      RECT 8.355 0.255 8.655 0.585 ;
      RECT 8.36 2.105 8.655 2.465 ;
      RECT 8.485 0.585 8.655 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 1.445 3.535 1.615 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 0.765 4.455 0.935 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.425 4.915 0.595 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 0.765 5.835 0.935 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 0.765 7.215 0.935 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 0.425 7.675 0.595 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
    LAYER met1 ;
      RECT 3.305 1.415 3.595 1.46 ;
      RECT 3.305 1.46 5.895 1.6 ;
      RECT 3.305 1.6 3.595 1.645 ;
      RECT 4.225 0.735 4.515 0.78 ;
      RECT 4.225 0.78 7.275 0.92 ;
      RECT 4.225 0.92 4.515 0.965 ;
      RECT 4.685 0.395 4.975 0.44 ;
      RECT 4.685 0.44 7.735 0.58 ;
      RECT 4.685 0.58 4.975 0.625 ;
      RECT 5.605 0.735 5.895 0.78 ;
      RECT 5.605 0.92 5.895 0.965 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.985 0.735 7.275 0.78 ;
      RECT 6.985 0.92 7.275 0.965 ;
      RECT 7.445 0.395 7.735 0.44 ;
      RECT 7.445 0.58 7.735 0.625 ;
  END
END sky130_fd_sc_hd__xor3_1
MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.965 1.075 8.375 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145 0.995 7.315 1.445 ;
        RECT 7.145 1.445 7.725 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.32 0.995 2.955 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.66 1.05 0.925 ;
        RECT 0.545 0.925 0.86 1.44 ;
        RECT 0.545 1.44 1.07 2.045 ;
        RECT 0.8 0.35 1.05 0.66 ;
        RECT 0.82 2.045 1.07 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.3 0.085 0.63 0.465 ;
      RECT 0.3 2.215 0.65 2.635 ;
      RECT 1.21 0.995 1.41 1.325 ;
      RECT 1.22 0.085 1.47 0.525 ;
      RECT 1.24 0.695 1.81 0.865 ;
      RECT 1.24 0.865 1.41 0.995 ;
      RECT 1.24 1.325 1.41 1.875 ;
      RECT 1.24 1.875 1.93 2.045 ;
      RECT 1.24 2.215 1.575 2.635 ;
      RECT 1.64 0.255 3.2 0.425 ;
      RECT 1.64 0.425 1.81 0.695 ;
      RECT 1.645 1.535 3.295 1.705 ;
      RECT 1.76 2.045 1.93 2.235 ;
      RECT 1.76 2.235 3.355 2.405 ;
      RECT 1.98 0.595 2.15 1.535 ;
      RECT 2.33 1.895 3.635 2.065 ;
      RECT 2.43 0.655 3.54 0.825 ;
      RECT 2.85 0.425 3.2 0.455 ;
      RECT 3.125 0.995 3.4 1.325 ;
      RECT 3.125 1.325 3.295 1.535 ;
      RECT 3.37 0.255 4.22 0.425 ;
      RECT 3.37 0.425 3.54 0.655 ;
      RECT 3.465 1.525 3.995 1.695 ;
      RECT 3.465 1.695 3.635 1.895 ;
      RECT 3.57 2.235 3.975 2.405 ;
      RECT 3.71 0.595 3.88 1.375 ;
      RECT 3.71 1.375 3.995 1.525 ;
      RECT 3.805 1.895 4.98 2.065 ;
      RECT 3.805 2.065 3.975 2.235 ;
      RECT 4.05 0.425 4.22 1.035 ;
      RECT 4.05 1.035 4.335 1.205 ;
      RECT 4.145 2.235 4.475 2.635 ;
      RECT 4.165 1.205 4.335 1.895 ;
      RECT 4.39 0.085 4.56 0.865 ;
      RECT 4.565 1.445 4.98 1.715 ;
      RECT 4.74 0.415 4.98 1.445 ;
      RECT 4.81 2.065 4.98 2.275 ;
      RECT 4.81 2.275 7.905 2.445 ;
      RECT 5.155 0.265 5.57 0.485 ;
      RECT 5.155 0.485 5.375 0.595 ;
      RECT 5.155 0.595 5.325 2.105 ;
      RECT 5.495 0.72 5.91 0.825 ;
      RECT 5.495 0.825 5.715 0.89 ;
      RECT 5.495 0.89 5.665 2.275 ;
      RECT 5.545 0.655 5.91 0.72 ;
      RECT 5.74 0.32 5.91 0.655 ;
      RECT 5.855 1.445 6.635 1.615 ;
      RECT 5.855 1.615 6.27 2.045 ;
      RECT 5.87 0.995 6.295 1.27 ;
      RECT 6.08 0.63 6.295 0.995 ;
      RECT 6.465 0.255 7.61 0.425 ;
      RECT 6.465 0.425 6.635 1.445 ;
      RECT 6.805 0.595 6.975 1.935 ;
      RECT 6.805 1.935 9.115 2.105 ;
      RECT 7.145 0.425 7.61 0.465 ;
      RECT 7.485 0.73 7.69 0.945 ;
      RECT 7.485 0.945 7.795 1.275 ;
      RECT 7.895 1.495 8.715 1.705 ;
      RECT 7.935 0.295 8.225 0.735 ;
      RECT 7.935 0.735 8.715 0.75 ;
      RECT 7.975 0.75 8.715 0.905 ;
      RECT 8.315 2.275 8.65 2.635 ;
      RECT 8.395 0.085 8.565 0.565 ;
      RECT 8.545 0.905 8.715 0.995 ;
      RECT 8.545 0.995 8.775 1.325 ;
      RECT 8.545 1.325 8.715 1.495 ;
      RECT 8.63 1.875 9.115 1.935 ;
      RECT 8.815 0.255 9.115 0.585 ;
      RECT 8.82 2.105 9.115 2.465 ;
      RECT 8.945 0.585 9.115 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.445 3.995 1.615 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.425 5.375 0.595 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 0.765 6.295 0.935 ;
      RECT 6.125 1.445 6.295 1.615 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 0.765 7.675 0.935 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 0.425 8.135 0.595 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
    LAYER met1 ;
      RECT 3.765 1.415 4.055 1.46 ;
      RECT 3.765 1.46 6.355 1.6 ;
      RECT 3.765 1.6 4.055 1.645 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.78 7.735 0.92 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 0.395 5.435 0.44 ;
      RECT 5.145 0.44 8.195 0.58 ;
      RECT 5.145 0.58 5.435 0.625 ;
      RECT 6.065 0.735 6.355 0.78 ;
      RECT 6.065 0.92 6.355 0.965 ;
      RECT 6.065 1.415 6.355 1.46 ;
      RECT 6.065 1.6 6.355 1.645 ;
      RECT 7.445 0.735 7.735 0.78 ;
      RECT 7.445 0.92 7.735 0.965 ;
      RECT 7.905 0.395 8.195 0.44 ;
      RECT 7.905 0.58 8.195 0.625 ;
  END
END sky130_fd_sc_hd__xor3_2
MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.525 1.075 8.935 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705 0.995 7.875 1.445 ;
        RECT 7.705 1.445 8.285 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.88 0.995 3.515 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.35 0.765 0.66 ;
        RECT 0.595 0.66 1.605 0.83 ;
        RECT 0.595 0.83 1.535 0.925 ;
        RECT 0.695 1.44 1.42 1.455 ;
        RECT 0.695 1.455 1.705 2.045 ;
        RECT 0.695 2.045 0.865 2.465 ;
        RECT 1.105 0.925 1.42 1.44 ;
        RECT 1.435 0.35 1.605 0.66 ;
        RECT 1.535 2.045 1.705 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.175 0.085 0.345 0.545 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.855 0.085 2.025 0.525 ;
        RECT 4.95 0.085 5.12 0.885 ;
        RECT 8.995 0.085 9.165 0.565 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.235 -0.085 0.405 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.275 2.135 0.445 2.635 ;
        RECT 1.035 2.215 1.365 2.635 ;
        RECT 1.875 2.215 2.205 2.635 ;
        RECT 4.705 2.235 5.035 2.635 ;
        RECT 8.915 2.275 9.245 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.82 0.965 2.045 1.325 ;
      RECT 1.875 0.695 2.365 0.865 ;
      RECT 1.875 0.865 2.045 0.965 ;
      RECT 1.875 1.325 2.045 1.875 ;
      RECT 1.875 1.875 2.545 2.045 ;
      RECT 2.195 0.255 3.76 0.425 ;
      RECT 2.195 0.425 2.365 0.695 ;
      RECT 2.37 1.535 3.855 1.705 ;
      RECT 2.375 2.045 2.545 2.235 ;
      RECT 2.375 2.235 3.915 2.405 ;
      RECT 2.54 0.595 2.71 1.535 ;
      RECT 2.89 1.895 4.195 2.065 ;
      RECT 2.99 0.655 4.1 0.825 ;
      RECT 3.41 0.425 3.76 0.455 ;
      RECT 3.685 0.995 4.055 1.325 ;
      RECT 3.685 1.325 3.855 1.535 ;
      RECT 3.93 0.255 4.78 0.425 ;
      RECT 3.93 0.425 4.1 0.655 ;
      RECT 4.025 1.525 4.555 1.695 ;
      RECT 4.025 1.695 4.195 1.895 ;
      RECT 4.13 2.235 4.535 2.405 ;
      RECT 4.27 0.595 4.44 1.375 ;
      RECT 4.27 1.375 4.555 1.525 ;
      RECT 4.365 1.895 5.54 2.065 ;
      RECT 4.365 2.065 4.535 2.235 ;
      RECT 4.61 0.425 4.78 1.035 ;
      RECT 4.61 1.035 4.865 1.04 ;
      RECT 4.61 1.04 4.88 1.045 ;
      RECT 4.61 1.045 4.89 1.05 ;
      RECT 4.61 1.05 4.895 1.205 ;
      RECT 4.725 1.205 4.895 1.895 ;
      RECT 5.125 1.445 5.54 1.715 ;
      RECT 5.3 0.415 5.54 1.445 ;
      RECT 5.37 2.065 5.54 2.275 ;
      RECT 5.37 2.275 8.465 2.445 ;
      RECT 5.715 0.265 6.13 0.485 ;
      RECT 5.715 0.485 5.935 0.595 ;
      RECT 5.715 0.595 5.885 2.105 ;
      RECT 6.075 0.72 6.47 0.825 ;
      RECT 6.075 0.825 6.275 0.89 ;
      RECT 6.075 0.89 6.245 2.275 ;
      RECT 6.105 0.655 6.47 0.72 ;
      RECT 6.3 0.32 6.47 0.655 ;
      RECT 6.415 1.445 7.195 1.615 ;
      RECT 6.415 1.615 6.83 2.045 ;
      RECT 6.43 0.995 6.855 1.27 ;
      RECT 6.64 0.63 6.855 0.995 ;
      RECT 7.025 0.255 8.17 0.425 ;
      RECT 7.025 0.425 7.195 1.445 ;
      RECT 7.365 0.595 7.535 1.935 ;
      RECT 7.365 1.935 9.675 2.105 ;
      RECT 7.705 0.425 8.17 0.465 ;
      RECT 8.045 0.73 8.25 0.945 ;
      RECT 8.045 0.945 8.355 1.275 ;
      RECT 8.455 1.495 9.275 1.705 ;
      RECT 8.495 0.295 8.785 0.735 ;
      RECT 8.495 0.735 9.275 0.75 ;
      RECT 8.535 0.75 9.275 0.905 ;
      RECT 9.105 0.905 9.275 0.995 ;
      RECT 9.105 0.995 9.335 1.325 ;
      RECT 9.105 1.325 9.275 1.495 ;
      RECT 9.19 1.875 9.675 1.935 ;
      RECT 9.415 0.255 9.675 0.585 ;
      RECT 9.415 2.105 9.675 2.465 ;
      RECT 9.505 0.585 9.675 1.875 ;
    LAYER mcon ;
      RECT 4.385 1.445 4.555 1.615 ;
      RECT 5.305 0.765 5.475 0.935 ;
      RECT 5.765 0.425 5.935 0.595 ;
      RECT 6.685 0.765 6.855 0.935 ;
      RECT 6.685 1.445 6.855 1.615 ;
      RECT 8.065 0.765 8.235 0.935 ;
      RECT 8.525 0.425 8.695 0.595 ;
    LAYER met1 ;
      RECT 4.325 1.415 4.615 1.46 ;
      RECT 4.325 1.46 6.915 1.6 ;
      RECT 4.325 1.6 4.615 1.645 ;
      RECT 5.245 0.735 5.535 0.78 ;
      RECT 5.245 0.78 8.295 0.92 ;
      RECT 5.245 0.92 5.535 0.965 ;
      RECT 5.705 0.395 5.995 0.44 ;
      RECT 5.705 0.44 8.755 0.58 ;
      RECT 5.705 0.58 5.995 0.625 ;
      RECT 6.625 0.735 6.915 0.78 ;
      RECT 6.625 0.92 6.915 0.965 ;
      RECT 6.625 1.415 6.915 1.46 ;
      RECT 6.625 1.6 6.915 1.645 ;
      RECT 8.005 0.735 8.295 0.78 ;
      RECT 8.005 0.92 8.295 0.965 ;
      RECT 8.465 0.395 8.755 0.44 ;
      RECT 8.465 0.58 8.755 0.625 ;
  END
END sky130_fd_sc_hd__xor3_4
MACRO sky130_fd_sc_hd__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.105 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.055 2.155 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.055 3.075 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.055 4.385 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.085 1.055 5.895 1.315 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.485 5.895 1.725 ;
        RECT 2.415 1.725 2.665 2.125 ;
        RECT 3.335 1.725 3.505 2.465 ;
        RECT 4.515 1.725 4.825 2.465 ;
        RECT 4.555 0.655 5.895 0.885 ;
        RECT 4.555 0.885 4.915 1.485 ;
        RECT 5.495 1.725 5.895 2.465 ;
        RECT 5.515 0.255 5.895 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.255 0.485 0.655 ;
      RECT 0.085 0.655 4.385 0.885 ;
      RECT 0.085 1.485 2.225 1.725 ;
      RECT 0.085 1.725 0.465 2.465 ;
      RECT 0.635 1.895 0.965 2.635 ;
      RECT 0.655 0.085 0.985 0.485 ;
      RECT 1.135 1.725 1.305 2.465 ;
      RECT 1.155 0.255 1.325 0.655 ;
      RECT 1.475 1.895 1.805 2.295 ;
      RECT 1.475 2.295 3.165 2.465 ;
      RECT 1.495 0.085 1.825 0.485 ;
      RECT 1.975 1.725 2.225 2.125 ;
      RECT 1.995 0.255 2.165 0.655 ;
      RECT 2.335 0.085 3.105 0.485 ;
      RECT 2.835 1.895 3.165 2.295 ;
      RECT 3.275 0.255 3.445 0.655 ;
      RECT 3.615 0.255 5.345 0.485 ;
      RECT 3.675 1.895 4.345 2.635 ;
      RECT 4.995 1.895 5.325 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__o311ai_2
MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.775 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.055 3.615 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.055 5.885 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.055 7.695 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.865 1.055 9.09 1.315 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.241000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055 1.485 9.575 1.725 ;
        RECT 4.055 1.725 4.305 2.115 ;
        RECT 4.975 1.725 5.145 2.115 ;
        RECT 5.815 1.725 6.005 2.465 ;
        RECT 6.675 1.725 6.845 2.465 ;
        RECT 7.515 1.725 7.685 2.465 ;
        RECT 7.895 0.655 9.575 0.885 ;
        RECT 8.355 1.725 8.525 2.465 ;
        RECT 9.195 1.725 9.575 2.465 ;
        RECT 9.26 0.885 9.575 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.085 0.085 0.505 0.885 ;
      RECT 0.085 1.485 3.865 1.725 ;
      RECT 0.085 1.725 0.405 2.465 ;
      RECT 0.595 1.895 0.925 2.635 ;
      RECT 0.675 0.255 0.845 0.655 ;
      RECT 0.675 0.655 7.385 0.885 ;
      RECT 1.015 0.085 1.345 0.485 ;
      RECT 1.095 1.725 1.265 2.465 ;
      RECT 1.435 1.895 1.765 2.635 ;
      RECT 1.515 0.255 1.685 0.655 ;
      RECT 1.855 0.085 2.185 0.485 ;
      RECT 1.935 1.725 2.105 2.465 ;
      RECT 2.275 1.895 2.605 2.295 ;
      RECT 2.275 2.295 5.645 2.465 ;
      RECT 2.355 0.255 2.525 0.655 ;
      RECT 2.695 0.085 3.025 0.485 ;
      RECT 2.775 1.725 2.945 2.115 ;
      RECT 3.115 1.895 3.445 2.295 ;
      RECT 3.195 0.255 3.365 0.655 ;
      RECT 3.535 0.085 3.885 0.485 ;
      RECT 3.615 1.725 3.865 2.115 ;
      RECT 4.055 0.255 4.225 0.655 ;
      RECT 4.395 0.085 4.725 0.485 ;
      RECT 4.475 1.895 4.805 2.295 ;
      RECT 4.895 0.255 5.065 0.655 ;
      RECT 5.235 0.085 5.585 0.485 ;
      RECT 5.315 1.895 5.645 2.295 ;
      RECT 5.755 0.255 9.575 0.485 ;
      RECT 6.175 1.895 6.505 2.635 ;
      RECT 7.015 1.895 7.345 2.635 ;
      RECT 7.555 0.485 7.725 0.885 ;
      RECT 7.855 1.895 8.185 2.635 ;
      RECT 8.695 1.895 9.025 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__o311ai_4
MACRO sky130_fd_sc_hd__o311ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.78 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.26 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 0.995 1.78 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.32 2.2 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.83 0.995 3.135 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.942000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 1.495 3.135 1.665 ;
        RECT 1.43 1.665 1.98 2.465 ;
        RECT 2.445 0.255 3.135 0.825 ;
        RECT 2.445 0.825 2.66 1.495 ;
        RECT 2.65 1.665 3.135 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.57 0.825 ;
      RECT 0.085 1.495 0.78 2.635 ;
      RECT 0.74 0.255 0.91 0.655 ;
      RECT 0.74 0.655 1.75 0.825 ;
      RECT 1.08 0.085 1.41 0.485 ;
      RECT 1.58 0.255 1.75 0.655 ;
      RECT 2.15 1.835 2.48 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o311ai_1
MACRO sky130_fd_sc_hd__o311ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.57 0.995 ;
        RECT 0.085 0.995 0.78 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.26 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 0.995 1.78 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.26 2.2 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.83 0.765 3.135 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.604000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 1.495 3.135 1.665 ;
        RECT 1.43 1.665 1.98 2.465 ;
        RECT 2.445 0.255 3.135 0.595 ;
        RECT 2.445 0.595 2.66 1.495 ;
        RECT 2.65 1.665 3.135 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.57 0.595 ;
      RECT 0.085 1.795 0.78 2.635 ;
      RECT 0.74 0.255 0.91 0.655 ;
      RECT 0.74 0.655 1.75 0.825 ;
      RECT 1.08 0.085 1.41 0.485 ;
      RECT 1.58 0.255 1.75 0.655 ;
      RECT 2.15 1.835 2.48 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o311ai_0
MACRO sky130_fd_sc_hd__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.765 2.155 0.995 ;
        RECT 1.965 0.995 2.31 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.75 1.705 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.24 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.62 0.995 3.095 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.995 3.535 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.454000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.395 0.67 ;
        RECT 0.085 0.67 0.255 1.785 ;
        RECT 0.085 1.785 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.425 0.995 0.735 1.325 ;
      RECT 0.565 0.655 1.26 0.825 ;
      RECT 0.565 0.825 0.735 0.995 ;
      RECT 0.565 1.325 0.735 1.495 ;
      RECT 0.565 1.495 3.505 1.665 ;
      RECT 0.59 0.085 0.92 0.465 ;
      RECT 0.595 2.175 0.84 2.635 ;
      RECT 1.015 1.835 2.575 2.005 ;
      RECT 1.015 2.005 1.265 2.465 ;
      RECT 1.09 0.255 2.495 0.425 ;
      RECT 1.09 0.425 1.26 0.655 ;
      RECT 1.455 2.255 2.125 2.635 ;
      RECT 2.325 0.425 2.495 0.655 ;
      RECT 2.325 0.655 3.505 0.825 ;
      RECT 2.325 2.005 2.575 2.465 ;
      RECT 2.765 0.085 3.095 0.485 ;
      RECT 3.335 0.255 3.505 0.655 ;
      RECT 3.335 1.665 3.505 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a311o_1
MACRO sky130_fd_sc_hd__a311o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.605 2.62 0.995 ;
        RECT 2.44 0.995 2.675 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.605 2.165 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.71 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.995 3.235 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695 0.995 4.005 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.295 0.845 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.085 0.345 0.885 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 1.015 0.085 1.345 0.465 ;
      RECT 1.015 0.655 1.695 0.825 ;
      RECT 1.015 0.825 1.185 1.495 ;
      RECT 1.015 1.495 3.965 1.665 ;
      RECT 1.16 1.835 1.38 2.635 ;
      RECT 1.525 0.255 2.96 0.425 ;
      RECT 1.525 0.425 1.695 0.655 ;
      RECT 1.59 1.835 3.025 2.005 ;
      RECT 1.59 2.005 1.84 2.465 ;
      RECT 2.125 2.255 2.455 2.635 ;
      RECT 2.715 2.005 3.025 2.465 ;
      RECT 2.79 0.425 2.96 0.655 ;
      RECT 2.79 0.655 3.965 0.825 ;
      RECT 3.22 0.085 3.55 0.485 ;
      RECT 3.795 0.255 3.965 0.655 ;
      RECT 3.795 1.665 3.965 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__a311o_2
MACRO sky130_fd_sc_hd__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.075 7.275 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255 1.075 6.04 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.515 1.075 4.945 1.285 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.505 1.285 ;
        RECT 1.06 1.285 1.255 1.625 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.745 0.35 1.625 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.904000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 0.295 2.545 0.465 ;
        RECT 2.295 0.465 2.465 0.715 ;
        RECT 2.295 0.715 3.305 0.885 ;
        RECT 2.715 1.545 3.885 1.715 ;
        RECT 2.91 0.885 3.105 1.545 ;
        RECT 3.055 0.295 3.385 0.465 ;
        RECT 3.135 0.465 3.305 0.715 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.095 0.085 0.345 0.565 ;
      RECT 0.175 1.795 0.345 2.295 ;
      RECT 0.175 2.295 2.025 2.465 ;
      RECT 0.515 0.295 0.845 0.465 ;
      RECT 0.515 1.955 0.845 2.125 ;
      RECT 0.595 0.465 0.765 0.715 ;
      RECT 0.595 0.715 2.025 0.885 ;
      RECT 0.595 0.885 0.765 1.955 ;
      RECT 1.015 0.085 1.185 0.545 ;
      RECT 1.015 1.795 1.185 2.295 ;
      RECT 1.355 0.295 1.685 0.465 ;
      RECT 1.435 0.465 1.605 0.715 ;
      RECT 1.435 1.455 2.385 1.625 ;
      RECT 1.435 1.625 1.605 2.125 ;
      RECT 1.855 0.085 2.025 0.545 ;
      RECT 1.855 0.885 2.025 1.075 ;
      RECT 1.855 1.075 2.705 1.245 ;
      RECT 1.855 1.795 2.025 2.295 ;
      RECT 2.195 1.625 2.385 1.915 ;
      RECT 2.195 1.915 6.765 2.085 ;
      RECT 2.295 2.255 2.625 2.635 ;
      RECT 2.715 0.085 2.885 0.545 ;
      RECT 3.135 2.255 3.465 2.635 ;
      RECT 3.275 1.075 4.32 1.245 ;
      RECT 3.555 0.085 4.065 0.545 ;
      RECT 3.975 2.255 4.305 2.635 ;
      RECT 4.15 1.245 4.32 1.455 ;
      RECT 4.15 1.455 6.685 1.625 ;
      RECT 4.275 0.295 4.605 0.465 ;
      RECT 4.355 0.465 4.525 0.715 ;
      RECT 4.355 0.715 6.005 0.885 ;
      RECT 4.475 1.795 4.645 1.915 ;
      RECT 4.475 2.085 4.645 2.465 ;
      RECT 4.775 0.085 4.945 0.545 ;
      RECT 4.815 2.255 5.175 2.635 ;
      RECT 5.255 0.255 7.27 0.425 ;
      RECT 5.255 0.425 6.345 0.465 ;
      RECT 5.375 1.795 5.545 1.915 ;
      RECT 5.375 2.085 5.545 2.465 ;
      RECT 5.675 0.645 6.005 0.715 ;
      RECT 5.715 2.255 6.045 2.635 ;
      RECT 6.175 0.465 6.345 0.885 ;
      RECT 6.515 0.645 6.845 0.825 ;
      RECT 6.515 0.825 6.685 1.455 ;
      RECT 6.595 1.795 6.765 1.915 ;
      RECT 6.595 2.085 6.765 2.465 ;
      RECT 6.935 0.425 7.27 0.5 ;
      RECT 6.935 1.795 7.27 2.635 ;
      RECT 7.015 0.5 7.27 0.905 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__a311o_4
MACRO sky130_fd_sc_hd__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.255 2.265 1.415 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615 0.815 1.785 1.615 ;
        RECT 1.615 1.615 2.625 1.785 ;
        RECT 2.435 0.255 2.625 1.615 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.105 1.325 ;
        RECT 0.935 1.325 1.105 2.295 ;
        RECT 0.935 2.295 2.965 2.465 ;
        RECT 2.795 1.44 3.545 1.63 ;
        RECT 2.795 1.63 2.965 2.295 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.255 0.345 0.825 ;
        RECT 0.09 0.825 0.26 1.495 ;
        RECT 0.09 1.495 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.42 -0.085 0.59 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.085 0.845 0.485 ;
      RECT 0.515 0.655 1.445 0.825 ;
      RECT 0.515 0.825 0.685 0.995 ;
      RECT 0.595 1.495 0.765 2.635 ;
      RECT 1.27 0.255 1.8 0.62 ;
      RECT 1.27 0.62 1.445 0.655 ;
      RECT 1.275 0.825 1.445 1.955 ;
      RECT 1.275 1.955 2.4 2.125 ;
      RECT 2.805 0.085 3.315 0.62 ;
      RECT 2.825 0.895 4.055 1.065 ;
      RECT 3.135 1.875 3.305 2.635 ;
      RECT 3.535 0.29 3.78 0.895 ;
      RECT 3.54 1.875 4.055 2.285 ;
      RECT 3.715 1.065 4.055 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__mux2_1
MACRO sky130_fd_sc_hd__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815 0.765 2.445 1.28 ;
        RECT 2.275 1.28 2.445 1.315 ;
        RECT 2.275 1.315 3.09 1.625 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625 0.735 3.09 1.025 ;
        RECT 2.9 0.42 3.09 0.735 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.36 0.755 3.55 1.625 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.765 0.75 ;
        RECT 0.515 0.75 0.685 1.595 ;
        RECT 0.515 1.595 0.825 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.085 0.345 0.885 ;
      RECT 0.09 1.495 0.345 2.635 ;
      RECT 0.855 0.995 1.165 1.325 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 0.995 0.635 1.605 0.805 ;
      RECT 0.995 0.805 1.165 0.995 ;
      RECT 0.995 1.325 1.165 1.835 ;
      RECT 0.995 1.835 1.655 2.005 ;
      RECT 1.025 2.175 1.315 2.635 ;
      RECT 1.335 0.995 1.505 1.495 ;
      RECT 1.335 1.495 1.995 1.665 ;
      RECT 1.435 0.295 2.73 0.465 ;
      RECT 1.435 0.465 1.605 0.635 ;
      RECT 1.485 2.005 1.655 2.255 ;
      RECT 1.485 2.255 2.795 2.425 ;
      RECT 1.825 1.665 1.995 1.835 ;
      RECT 1.825 1.835 4.05 2.005 ;
      RECT 3.325 2.175 3.545 2.635 ;
      RECT 3.35 0.085 3.55 0.585 ;
      RECT 3.715 2.005 4.05 2.465 ;
      RECT 3.72 0.255 4.05 1.835 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__mux2_2
MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.995 1.75 1.615 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.435 1.325 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.74 1.325 ;
        RECT 0.57 0.635 2.85 0.805 ;
        RECT 0.57 0.805 0.74 0.995 ;
        RECT 2.68 0.805 2.85 0.995 ;
        RECT 2.68 0.995 3.395 1.325 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.915 0.255 4.085 0.635 ;
        RECT 3.915 0.635 5.43 0.805 ;
        RECT 3.915 1.575 5.43 1.745 ;
        RECT 3.915 1.745 4.085 2.465 ;
        RECT 4.755 0.255 4.925 0.635 ;
        RECT 4.755 1.745 4.925 2.465 ;
        RECT 5.2 0.805 5.43 1.575 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.09 0.295 0.345 0.625 ;
      RECT 0.09 0.625 0.26 1.495 ;
      RECT 0.09 1.495 1.08 1.665 ;
      RECT 0.09 1.665 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 1.835 0.82 2.635 ;
      RECT 0.91 0.995 1.08 1.495 ;
      RECT 0.99 1.935 1.34 2.275 ;
      RECT 0.99 2.275 2.77 2.445 ;
      RECT 1.53 1.935 3.245 2.105 ;
      RECT 1.975 0.295 3.23 0.465 ;
      RECT 1.98 1.595 3.735 1.765 ;
      RECT 3.06 0.465 3.23 0.655 ;
      RECT 3.06 0.655 3.735 0.825 ;
      RECT 3.075 2.105 3.245 2.465 ;
      RECT 3.415 0.085 3.745 0.465 ;
      RECT 3.415 2.255 3.745 2.635 ;
      RECT 3.565 0.825 3.735 1.075 ;
      RECT 3.565 1.075 5.03 1.245 ;
      RECT 3.565 1.245 3.735 1.595 ;
      RECT 3.565 1.765 3.735 1.785 ;
      RECT 4.255 0.085 4.585 0.465 ;
      RECT 4.255 1.915 4.585 2.635 ;
      RECT 5.095 0.085 5.425 0.465 ;
      RECT 5.095 1.915 5.425 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__mux2_4
MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.18 0.645 6.895 0.815 ;
        RECT 5.18 0.815 5.35 1.325 ;
        RECT 5.305 0.425 5.89 0.645 ;
        RECT 6.725 0.815 6.895 0.995 ;
        RECT 6.725 0.995 7.195 1.165 ;
        RECT 7.025 1.165 7.195 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.29 1.105 4.475 1.275 ;
        RECT 4.305 0.995 4.475 1.105 ;
        RECT 4.305 1.275 4.475 1.325 ;
      LAYER mcon ;
        RECT 4.29 1.105 4.46 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.96 0.995 8.245 1.325 ;
      LAYER mcon ;
        RECT 7.96 1.105 8.13 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.23 1.075 4.52 1.12 ;
        RECT 4.23 1.12 8.19 1.26 ;
        RECT 4.23 1.26 4.52 1.305 ;
        RECT 7.9 1.075 8.19 1.12 ;
        RECT 7.9 1.26 8.19 1.305 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.739500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795 0.995 3.965 1.495 ;
        RECT 3.795 1.495 6.035 1.665 ;
        RECT 5.67 0.995 6.035 1.495 ;
      LAYER mcon ;
        RECT 5.67 1.445 5.84 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.215 0.995 9.51 1.615 ;
      LAYER mcon ;
        RECT 9.34 1.445 9.51 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.61 1.415 5.9 1.46 ;
        RECT 5.61 1.46 9.57 1.6 ;
        RECT 5.61 1.6 5.9 1.645 ;
        RECT 9.28 1.415 9.57 1.46 ;
        RECT 9.28 1.6 9.57 1.645 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 0.635 3.285 0.805 ;
        RECT 0.595 0.805 0.815 1.575 ;
        RECT 0.595 1.575 3.285 1.745 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 0.295 1.605 0.635 ;
        RECT 1.435 1.745 1.605 2.465 ;
        RECT 2.275 0.255 2.445 0.635 ;
        RECT 2.275 1.745 2.445 2.465 ;
        RECT 3.115 0.295 3.285 0.635 ;
        RECT 3.115 1.745 3.285 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.09 0.085 0.425 0.465 ;
      RECT 0.09 1.915 0.425 2.635 ;
      RECT 0.935 0.085 1.265 0.465 ;
      RECT 0.935 1.915 1.265 2.635 ;
      RECT 0.985 1.075 3.625 1.245 ;
      RECT 1.775 0.085 2.105 0.465 ;
      RECT 1.775 1.915 2.105 2.635 ;
      RECT 2.615 0.085 2.945 0.465 ;
      RECT 2.615 1.915 2.945 2.635 ;
      RECT 3.455 0.085 3.785 0.465 ;
      RECT 3.455 0.635 4.92 0.805 ;
      RECT 3.455 0.805 3.625 1.075 ;
      RECT 3.455 1.245 3.625 1.835 ;
      RECT 3.455 1.835 8.225 2.005 ;
      RECT 3.455 2.255 3.785 2.635 ;
      RECT 3.955 0.295 5.125 0.465 ;
      RECT 3.955 2.255 5.905 2.425 ;
      RECT 4.75 0.805 4.92 0.935 ;
      RECT 6.06 0.085 6.39 0.465 ;
      RECT 6.075 2.175 6.245 2.635 ;
      RECT 6.345 0.995 6.515 1.495 ;
      RECT 6.345 1.495 8.855 1.665 ;
      RECT 6.48 2.255 8.645 2.425 ;
      RECT 6.575 0.295 7.865 0.465 ;
      RECT 7.115 0.635 7.67 0.805 ;
      RECT 7.5 0.805 7.67 0.935 ;
      RECT 8.685 0.645 9.485 0.815 ;
      RECT 8.685 0.815 8.855 1.495 ;
      RECT 8.685 1.665 8.855 1.915 ;
      RECT 8.685 1.915 9.485 2.085 ;
      RECT 8.815 0.085 9.145 0.465 ;
      RECT 8.815 2.255 9.145 2.635 ;
      RECT 9.315 0.295 9.485 0.645 ;
      RECT 9.315 1.795 9.485 1.915 ;
      RECT 9.315 2.085 9.485 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.75 0.765 4.92 0.935 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.5 0.765 7.67 0.935 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 4.69 0.735 4.98 0.78 ;
      RECT 4.69 0.78 7.73 0.92 ;
      RECT 4.69 0.92 4.98 0.965 ;
      RECT 7.44 0.735 7.73 0.78 ;
      RECT 7.44 0.92 7.73 0.965 ;
  END
END sky130_fd_sc_hd__mux2_8
MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.23 0.26 3.56 0.735 ;
        RECT 3.23 0.735 6.815 0.905 ;
        RECT 3.23 1.445 6.815 1.615 ;
        RECT 3.23 1.615 3.56 2.465 ;
        RECT 4.07 0.26 4.4 0.735 ;
        RECT 4.07 1.615 4.4 2.465 ;
        RECT 4.91 0.26 5.24 0.735 ;
        RECT 4.91 1.615 5.24 2.465 ;
        RECT 5.75 0.26 6.08 0.735 ;
        RECT 5.75 1.615 6.08 2.465 ;
        RECT 6.435 0.905 6.815 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.095 0.26 0.425 0.735 ;
      RECT 0.095 0.735 0.78 0.905 ;
      RECT 0.095 1.445 0.78 1.615 ;
      RECT 0.095 1.615 0.425 2.16 ;
      RECT 0.595 0.085 0.765 0.565 ;
      RECT 0.595 1.785 0.765 2.635 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 0.995 1.04 1.325 ;
      RECT 0.61 1.325 0.78 1.445 ;
      RECT 1 0.26 1.38 0.825 ;
      RECT 1 1.545 1.38 2.465 ;
      RECT 1.21 0.825 1.38 1.075 ;
      RECT 1.21 1.075 2.72 1.275 ;
      RECT 1.21 1.275 1.38 1.545 ;
      RECT 1.55 0.26 1.88 0.735 ;
      RECT 1.55 0.735 3.06 0.905 ;
      RECT 1.55 1.445 3.06 1.615 ;
      RECT 1.55 1.615 1.88 2.465 ;
      RECT 2.05 0.085 2.22 0.565 ;
      RECT 2.05 1.785 2.22 2.635 ;
      RECT 2.39 0.26 2.72 0.735 ;
      RECT 2.39 1.615 2.72 2.465 ;
      RECT 2.89 0.085 3.06 0.565 ;
      RECT 2.89 0.905 3.06 1.075 ;
      RECT 2.89 1.075 5.36 1.275 ;
      RECT 2.89 1.275 3.06 1.445 ;
      RECT 2.89 1.785 3.06 2.635 ;
      RECT 3.73 0.085 3.9 0.565 ;
      RECT 3.73 1.835 3.9 2.635 ;
      RECT 4.57 0.085 4.74 0.565 ;
      RECT 4.57 1.835 4.74 2.635 ;
      RECT 5.41 0.085 5.58 0.565 ;
      RECT 5.41 1.835 5.58 2.635 ;
      RECT 6.25 0.085 6.42 0.565 ;
      RECT 6.25 1.835 6.42 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
  END
END sky130_fd_sc_hd__bufbuf_8
MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.255 5.485 0.26 ;
        RECT 5.235 0.26 5.565 0.735 ;
        RECT 5.235 0.735 11.875 0.905 ;
        RECT 5.235 1.445 11.875 1.615 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 6.075 0.26 6.405 0.735 ;
        RECT 6.075 1.615 6.405 2.465 ;
        RECT 6.155 0.255 6.325 0.26 ;
        RECT 6.915 0.26 7.245 0.735 ;
        RECT 6.915 1.615 7.245 2.465 ;
        RECT 6.995 0.255 7.165 0.26 ;
        RECT 7.755 0.26 8.085 0.735 ;
        RECT 7.755 1.615 8.085 2.465 ;
        RECT 8.595 0.26 8.925 0.735 ;
        RECT 8.595 1.615 8.925 2.465 ;
        RECT 9.435 0.26 9.765 0.735 ;
        RECT 9.435 1.615 9.765 2.465 ;
        RECT 10.275 0.26 10.605 0.735 ;
        RECT 10.275 1.615 10.605 2.465 ;
        RECT 11.115 0.26 11.445 0.735 ;
        RECT 11.115 1.615 11.445 2.465 ;
        RECT 11.62 0.905 11.875 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.15 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.175 0.085 0.345 0.905 ;
      RECT 0.175 1.445 0.345 2.635 ;
      RECT 0.515 0.26 0.845 0.905 ;
      RECT 0.515 1.445 0.845 2.465 ;
      RECT 0.61 0.905 0.845 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.845 1.445 ;
      RECT 1.035 0.26 1.365 0.735 ;
      RECT 1.035 0.735 2.545 0.905 ;
      RECT 1.035 1.445 2.545 1.615 ;
      RECT 1.035 1.615 1.365 2.465 ;
      RECT 1.535 0.085 1.705 0.565 ;
      RECT 1.535 1.785 1.705 2.635 ;
      RECT 1.875 0.26 2.205 0.735 ;
      RECT 1.875 1.615 2.205 2.465 ;
      RECT 2.375 0.085 2.545 0.565 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 4.685 1.275 ;
      RECT 2.375 1.275 2.545 1.445 ;
      RECT 2.375 1.785 2.545 2.635 ;
      RECT 2.715 0.26 3.045 0.735 ;
      RECT 2.715 0.735 5.065 0.905 ;
      RECT 2.715 1.445 5.065 1.615 ;
      RECT 2.715 1.615 3.045 2.465 ;
      RECT 3.215 0.085 3.385 0.565 ;
      RECT 3.215 1.835 3.385 2.635 ;
      RECT 3.555 0.26 3.885 0.735 ;
      RECT 3.555 1.615 3.885 2.465 ;
      RECT 4.055 0.085 4.225 0.565 ;
      RECT 4.055 1.835 4.225 2.635 ;
      RECT 4.395 0.26 4.725 0.735 ;
      RECT 4.395 1.615 4.725 2.465 ;
      RECT 4.89 0.905 5.065 1.075 ;
      RECT 4.89 1.075 11.45 1.275 ;
      RECT 4.89 1.275 5.065 1.445 ;
      RECT 4.895 0.085 5.065 0.565 ;
      RECT 4.895 1.835 5.065 2.635 ;
      RECT 5.735 0.085 5.905 0.565 ;
      RECT 5.735 1.835 5.905 2.635 ;
      RECT 6.575 0.085 6.745 0.565 ;
      RECT 6.575 1.835 6.745 2.635 ;
      RECT 7.415 0.085 7.585 0.565 ;
      RECT 7.415 1.835 7.585 2.635 ;
      RECT 8.255 0.085 8.425 0.565 ;
      RECT 8.255 1.835 8.425 2.635 ;
      RECT 9.095 0.085 9.265 0.565 ;
      RECT 9.095 1.835 9.265 2.635 ;
      RECT 9.935 0.085 10.105 0.565 ;
      RECT 9.935 1.835 10.105 2.635 ;
      RECT 10.775 0.085 10.945 0.565 ;
      RECT 10.775 1.835 10.945 2.635 ;
      RECT 11.615 0.085 11.785 0.565 ;
      RECT 11.615 1.835 11.785 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
  END
END sky130_fd_sc_hd__bufbuf_16
MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 0.995 1.24 1.615 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.495 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.25 1.055 5.58 1.675 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.8 1.055 5.045 1.675 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265 0.995 3.565 1.995 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 0.995 6.345 1.675 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315 0.255 9.575 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.175 0.26 0.345 0.635 ;
      RECT 0.175 0.635 1.185 0.805 ;
      RECT 0.175 1.795 1.705 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 1.015 0.255 2.09 0.425 ;
      RECT 1.015 0.425 1.185 0.635 ;
      RECT 1.015 2.135 1.185 2.295 ;
      RECT 1.015 2.295 2.545 2.465 ;
      RECT 1.41 0.595 1.75 0.765 ;
      RECT 1.41 0.765 1.7 0.935 ;
      RECT 1.41 0.935 1.58 1.455 ;
      RECT 1.41 1.455 2.045 1.625 ;
      RECT 1.535 1.965 1.705 2.125 ;
      RECT 1.875 1.625 2.045 1.955 ;
      RECT 1.875 1.955 2.205 2.125 ;
      RECT 1.92 0.425 2.09 0.76 ;
      RECT 2.08 1.105 2.62 1.285 ;
      RECT 2.26 0.43 2.62 1.105 ;
      RECT 2.26 1.285 2.62 1.395 ;
      RECT 2.26 1.395 3.065 1.625 ;
      RECT 2.375 1.795 2.545 2.295 ;
      RECT 2.715 1.625 3.065 2.465 ;
      RECT 2.8 0.085 3.09 0.805 ;
      RECT 3.235 2.255 3.565 2.635 ;
      RECT 3.38 0.255 4.98 0.425 ;
      RECT 3.38 0.425 3.55 0.795 ;
      RECT 3.72 0.595 4.05 0.845 ;
      RECT 3.735 0.845 4.05 0.92 ;
      RECT 3.735 0.92 3.905 1.445 ;
      RECT 3.735 1.445 4.495 1.615 ;
      RECT 3.825 1.785 3.995 2.295 ;
      RECT 3.825 2.295 4.835 2.465 ;
      RECT 4.075 1.095 4.405 1.105 ;
      RECT 4.075 1.105 4.46 1.265 ;
      RECT 4.165 1.615 4.495 2.125 ;
      RECT 4.22 0.595 4.39 0.715 ;
      RECT 4.22 0.715 5.74 0.885 ;
      RECT 4.22 0.885 4.39 0.925 ;
      RECT 4.29 1.265 4.46 1.275 ;
      RECT 4.625 0.425 4.98 0.465 ;
      RECT 4.665 1.915 5.73 2.085 ;
      RECT 4.665 2.085 4.835 2.295 ;
      RECT 5.06 2.255 5.39 2.635 ;
      RECT 5.15 0.085 5.32 0.545 ;
      RECT 5.495 0.295 5.74 0.715 ;
      RECT 5.56 2.085 5.73 2.465 ;
      RECT 5.98 2.255 6.33 2.635 ;
      RECT 6.01 0.085 6.34 0.465 ;
      RECT 6.5 2.135 6.685 2.465 ;
      RECT 6.51 0.325 6.685 0.655 ;
      RECT 6.515 0.655 6.685 1.105 ;
      RECT 6.515 1.105 6.805 1.275 ;
      RECT 6.515 1.275 6.685 2.135 ;
      RECT 6.98 0.765 7.22 0.935 ;
      RECT 6.98 0.935 7.15 2.135 ;
      RECT 6.98 2.135 7.19 2.465 ;
      RECT 7.03 0.255 7.2 0.415 ;
      RECT 7.03 0.415 7.56 0.585 ;
      RECT 7.36 2.255 7.69 2.295 ;
      RECT 7.36 2.295 8.645 2.465 ;
      RECT 7.39 0.585 7.56 1.755 ;
      RECT 7.39 1.755 8.175 1.985 ;
      RECT 7.73 0.255 8.725 0.425 ;
      RECT 7.73 0.425 7.9 0.585 ;
      RECT 7.845 1.985 8.175 2.125 ;
      RECT 7.97 0.765 8.385 0.925 ;
      RECT 7.97 0.925 8.38 0.935 ;
      RECT 8.19 1.105 8.645 1.275 ;
      RECT 8.21 0.595 8.385 0.765 ;
      RECT 8.475 1.665 9.125 1.835 ;
      RECT 8.475 1.835 8.645 2.295 ;
      RECT 8.555 0.425 8.725 0.715 ;
      RECT 8.555 0.715 9.125 0.885 ;
      RECT 8.815 2.255 9.145 2.635 ;
      RECT 8.895 0.085 9.065 0.545 ;
      RECT 8.955 0.885 9.125 1.665 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.45 1.105 2.62 1.275 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.29 1.105 4.46 1.275 ;
      RECT 4.325 1.785 4.495 1.955 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.635 1.105 6.805 1.275 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.05 0.765 7.22 0.935 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.555 1.785 7.725 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.475 1.105 8.645 1.275 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 8.2 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 2.39 1.075 2.68 1.12 ;
      RECT 2.39 1.12 4.52 1.26 ;
      RECT 2.39 1.26 2.68 1.305 ;
      RECT 4.23 1.075 4.52 1.12 ;
      RECT 4.23 1.26 4.52 1.305 ;
      RECT 4.265 1.755 4.555 1.8 ;
      RECT 4.265 1.8 7.785 1.94 ;
      RECT 4.265 1.94 4.555 1.985 ;
      RECT 6.575 1.075 6.865 1.12 ;
      RECT 6.575 1.12 8.705 1.26 ;
      RECT 6.575 1.26 6.865 1.305 ;
      RECT 6.99 0.735 7.28 0.78 ;
      RECT 6.99 0.92 7.28 0.965 ;
      RECT 7.495 1.755 7.785 1.8 ;
      RECT 7.495 1.94 7.785 1.985 ;
      RECT 7.91 0.735 8.2 0.78 ;
      RECT 7.91 0.92 8.2 0.965 ;
      RECT 8.415 1.075 8.705 1.12 ;
      RECT 8.415 1.26 8.705 1.305 ;
  END
END sky130_fd_sc_hd__mux4_1
MACRO sky130_fd_sc_hd__mux4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535 0.375 6.845 0.995 ;
        RECT 6.535 0.995 6.945 1.075 ;
        RECT 6.635 1.075 6.945 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.715 5.115 1.395 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 0.765 1.235 1.095 ;
        RECT 1.02 0.395 1.235 0.765 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.715 2.615 1.015 ;
        RECT 2.41 1.015 2.615 1.32 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.975 0.325 1.745 ;
      LAYER mcon ;
        RECT 0.145 1.445 0.315 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.005 1.445 1.39 1.615 ;
        RECT 1.22 1.285 1.39 1.445 ;
      LAYER mcon ;
        RECT 1.065 1.445 1.235 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.125 1.245 6.465 1.645 ;
      LAYER mcon ;
        RECT 6.125 1.445 6.295 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.415 0.375 1.46 ;
        RECT 0.085 1.46 6.355 1.6 ;
        RECT 0.085 1.6 0.375 1.645 ;
        RECT 1.005 1.415 1.295 1.46 ;
        RECT 1.005 1.6 1.295 1.645 ;
        RECT 6.065 1.415 6.355 1.46 ;
        RECT 6.065 1.6 6.355 1.645 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 0.715 3.075 1.32 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.355 1.835 7.765 2.455 ;
        RECT 7.435 0.265 7.765 0.725 ;
        RECT 7.455 1.495 7.765 1.835 ;
        RECT 7.595 0.725 7.765 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.665 0.805 ;
      RECT 0.175 1.915 1.9 1.955 ;
      RECT 0.175 1.955 0.665 2.085 ;
      RECT 0.175 2.085 0.345 2.375 ;
      RECT 0.495 0.805 0.665 1.785 ;
      RECT 0.495 1.785 1.9 1.915 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 1.405 0.705 1.73 1.035 ;
      RECT 1.41 2.125 2.24 2.295 ;
      RECT 1.47 0.365 2.07 0.535 ;
      RECT 1.56 1.035 1.73 1.575 ;
      RECT 1.56 1.575 1.9 1.785 ;
      RECT 1.9 0.535 2.07 1.235 ;
      RECT 1.9 1.235 2.24 1.405 ;
      RECT 2.07 1.405 2.24 2.125 ;
      RECT 2.45 0.085 2.78 0.545 ;
      RECT 2.595 2.055 2.825 2.635 ;
      RECT 2.97 1.785 3.315 1.955 ;
      RECT 2.985 0.295 3.415 0.465 ;
      RECT 3.145 1.49 3.415 1.66 ;
      RECT 3.145 1.66 3.315 1.785 ;
      RECT 3.245 0.465 3.415 1.06 ;
      RECT 3.245 1.06 3.48 1.39 ;
      RECT 3.245 1.39 3.415 1.49 ;
      RECT 3.305 2.125 3.82 2.295 ;
      RECT 3.565 1.81 3.82 2.125 ;
      RECT 3.585 0.345 3.82 0.675 ;
      RECT 3.65 0.675 3.82 1.81 ;
      RECT 3.99 0.345 4.18 2.125 ;
      RECT 3.99 2.125 4.515 2.295 ;
      RECT 4.395 0.255 4.6 0.585 ;
      RECT 4.395 0.585 4.565 1.565 ;
      RECT 4.395 1.565 5.495 1.735 ;
      RECT 4.395 1.735 4.585 1.895 ;
      RECT 4.755 2.005 5.1 2.635 ;
      RECT 4.795 0.085 5.125 0.545 ;
      RECT 5.325 0.295 6.22 0.465 ;
      RECT 5.325 0.465 5.495 1.565 ;
      RECT 5.325 1.735 5.495 2.155 ;
      RECT 5.325 2.155 6.275 2.325 ;
      RECT 5.665 0.705 6.285 1.035 ;
      RECT 5.665 1.035 5.955 1.985 ;
      RECT 6.525 2.125 6.845 2.295 ;
      RECT 6.675 1.495 7.285 1.665 ;
      RECT 6.675 1.665 6.845 2.125 ;
      RECT 7.015 0.085 7.265 0.815 ;
      RECT 7.015 1.835 7.185 2.635 ;
      RECT 7.115 0.995 7.425 1.325 ;
      RECT 7.115 1.325 7.285 1.495 ;
      RECT 7.935 0.085 8.19 0.885 ;
      RECT 7.935 1.495 8.185 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 1.785 1.695 1.955 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.125 2.155 2.295 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.125 3.535 2.295 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.125 4.455 2.295 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 1.785 5.835 1.955 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.125 6.755 2.295 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
    LAYER met1 ;
      RECT 1.465 1.755 1.755 1.8 ;
      RECT 1.465 1.8 5.895 1.94 ;
      RECT 1.465 1.94 1.755 1.985 ;
      RECT 1.925 2.095 2.215 2.14 ;
      RECT 1.925 2.14 3.595 2.28 ;
      RECT 1.925 2.28 2.215 2.325 ;
      RECT 3.305 2.095 3.595 2.14 ;
      RECT 3.305 2.28 3.595 2.325 ;
      RECT 4.225 2.095 4.515 2.14 ;
      RECT 4.225 2.14 6.815 2.28 ;
      RECT 4.225 2.28 4.515 2.325 ;
      RECT 5.605 1.755 5.895 1.8 ;
      RECT 5.605 1.94 5.895 1.985 ;
      RECT 6.525 2.095 6.815 2.14 ;
      RECT 6.525 2.28 6.815 2.325 ;
  END
END sky130_fd_sc_hd__mux4_2
MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.54 0.375 6.85 0.995 ;
        RECT 6.54 0.995 6.95 1.075 ;
        RECT 6.64 1.075 6.95 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.75 0.715 5.12 1.395 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 0.765 1.24 1.095 ;
        RECT 1.025 0.395 1.24 0.765 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245 0.715 2.62 1.015 ;
        RECT 2.415 1.015 2.62 1.32 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.975 0.33 1.745 ;
      LAYER mcon ;
        RECT 0.15 1.445 0.32 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.01 1.445 1.395 1.615 ;
        RECT 1.225 1.285 1.395 1.445 ;
      LAYER mcon ;
        RECT 1.07 1.445 1.24 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.13 1.245 6.47 1.645 ;
      LAYER mcon ;
        RECT 6.13 1.445 6.3 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.415 0.38 1.46 ;
        RECT 0.085 1.46 6.36 1.6 ;
        RECT 0.085 1.6 0.38 1.645 ;
        RECT 1.01 1.415 1.3 1.46 ;
        RECT 1.01 1.6 1.3 1.645 ;
        RECT 6.07 1.415 6.36 1.46 ;
        RECT 6.07 1.6 6.36 1.645 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.79 0.715 3.08 1.32 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.36 1.835 7.77 2.455 ;
        RECT 7.44 0.265 7.77 0.725 ;
        RECT 7.46 1.495 7.77 1.835 ;
        RECT 7.6 0.725 7.77 1.065 ;
        RECT 7.6 1.065 8.685 1.305 ;
        RECT 7.6 1.305 7.77 1.495 ;
        RECT 8.36 0.265 8.685 1.065 ;
        RECT 8.36 1.305 8.685 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.135 0.345 0.345 0.635 ;
      RECT 0.135 0.635 0.67 0.805 ;
      RECT 0.135 1.915 1.905 1.955 ;
      RECT 0.135 1.955 0.67 2.085 ;
      RECT 0.135 2.085 0.345 2.375 ;
      RECT 0.5 0.805 0.67 1.785 ;
      RECT 0.5 1.785 1.905 1.915 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 1.41 0.705 1.735 1.035 ;
      RECT 1.415 2.125 2.245 2.295 ;
      RECT 1.475 0.365 2.075 0.535 ;
      RECT 1.565 1.035 1.735 1.575 ;
      RECT 1.565 1.575 1.905 1.785 ;
      RECT 1.905 0.535 2.075 1.235 ;
      RECT 1.905 1.235 2.245 1.405 ;
      RECT 2.075 1.405 2.245 2.125 ;
      RECT 2.455 0.085 2.785 0.545 ;
      RECT 2.6 2.055 2.83 2.635 ;
      RECT 2.975 1.785 3.32 1.955 ;
      RECT 2.99 0.295 3.42 0.465 ;
      RECT 3.15 1.49 3.42 1.66 ;
      RECT 3.15 1.66 3.32 1.785 ;
      RECT 3.25 0.465 3.42 1.06 ;
      RECT 3.25 1.06 3.485 1.39 ;
      RECT 3.25 1.39 3.42 1.49 ;
      RECT 3.31 2.125 3.825 2.295 ;
      RECT 3.575 1.81 3.825 2.125 ;
      RECT 3.59 0.345 3.825 0.675 ;
      RECT 3.655 0.675 3.825 1.81 ;
      RECT 3.995 0.345 4.185 2.125 ;
      RECT 3.995 2.125 4.52 2.295 ;
      RECT 4.4 0.255 4.605 0.585 ;
      RECT 4.4 0.585 4.57 1.565 ;
      RECT 4.4 1.565 5.5 1.735 ;
      RECT 4.4 1.735 4.59 1.895 ;
      RECT 4.76 2.005 5.105 2.635 ;
      RECT 4.8 0.085 5.13 0.545 ;
      RECT 5.33 0.295 6.225 0.465 ;
      RECT 5.33 0.465 5.5 1.565 ;
      RECT 5.33 1.735 5.5 2.155 ;
      RECT 5.33 2.155 6.28 2.325 ;
      RECT 5.67 0.705 6.29 1.035 ;
      RECT 5.67 1.035 5.96 1.985 ;
      RECT 6.53 2.125 6.85 2.295 ;
      RECT 6.68 1.495 7.29 1.665 ;
      RECT 6.68 1.665 6.85 2.125 ;
      RECT 7.02 0.085 7.27 0.815 ;
      RECT 7.02 1.835 7.19 2.635 ;
      RECT 7.12 0.995 7.43 1.325 ;
      RECT 7.12 1.325 7.29 1.495 ;
      RECT 7.94 0.085 8.19 0.885 ;
      RECT 7.94 1.495 8.19 2.635 ;
      RECT 8.855 0.085 9.105 0.885 ;
      RECT 8.855 1.495 9.105 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.53 1.785 1.7 1.955 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.99 2.125 2.16 2.295 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.37 2.125 3.54 2.295 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.29 2.125 4.46 2.295 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.67 1.785 5.84 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.59 2.125 6.76 2.295 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
    LAYER met1 ;
      RECT 1.47 1.755 1.76 1.8 ;
      RECT 1.47 1.8 5.9 1.94 ;
      RECT 1.47 1.94 1.76 1.985 ;
      RECT 1.93 2.095 2.22 2.14 ;
      RECT 1.93 2.14 3.6 2.28 ;
      RECT 1.93 2.28 2.22 2.325 ;
      RECT 3.31 2.095 3.6 2.14 ;
      RECT 3.31 2.28 3.6 2.325 ;
      RECT 4.23 2.095 4.52 2.14 ;
      RECT 4.23 2.14 6.82 2.28 ;
      RECT 4.23 2.28 4.52 2.325 ;
      RECT 5.61 1.755 5.9 1.8 ;
      RECT 5.61 1.94 5.9 1.985 ;
      RECT 6.53 2.095 6.82 2.14 ;
      RECT 6.53 2.28 6.82 2.325 ;
  END
END sky130_fd_sc_hd__mux4_4
MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 5.965 1.445 8.265 1.615 ;
        RECT 8.095 1.075 9.575 1.275 ;
        RECT 8.095 1.275 8.265 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935 0.995 5.285 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415 0.995 3.765 1.325 ;
        RECT 3.595 1.325 3.765 1.445 ;
        RECT 3.595 1.445 5.795 1.615 ;
        RECT 5.465 1.075 5.795 1.445 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.335 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.905 ;
        RECT 0.575 1.445 1.705 1.615 ;
        RECT 0.575 1.615 0.825 2.125 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 1.615 1.665 2.125 ;
        RECT 1.505 0.905 1.705 1.095 ;
        RECT 1.505 1.095 3.245 1.275 ;
        RECT 1.505 1.275 1.705 1.445 ;
        RECT 3.075 0.645 5.68 0.735 ;
        RECT 3.075 0.735 7.765 0.82 ;
        RECT 3.075 0.82 3.245 1.095 ;
        RECT 5.51 0.82 6.46 0.905 ;
        RECT 6.29 0.645 7.765 0.735 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.09 1.445 0.405 2.295 ;
      RECT 0.09 2.295 2.125 2.465 ;
      RECT 0.115 0.085 0.365 0.895 ;
      RECT 0.995 1.785 1.245 2.295 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.875 0.085 2.045 0.645 ;
      RECT 1.875 0.645 2.905 0.925 ;
      RECT 1.875 1.445 3.03 1.615 ;
      RECT 1.875 1.615 2.125 2.295 ;
      RECT 2.235 0.255 5.585 0.425 ;
      RECT 2.235 0.425 2.61 0.475 ;
      RECT 2.315 1.795 2.565 2.215 ;
      RECT 2.315 2.215 6.005 2.465 ;
      RECT 2.735 0.595 2.905 0.645 ;
      RECT 2.735 1.615 3.03 1.835 ;
      RECT 2.735 1.835 5.585 2.045 ;
      RECT 3.035 0.425 5.585 0.475 ;
      RECT 5.755 1.785 8.605 2.045 ;
      RECT 5.755 2.045 6.005 2.215 ;
      RECT 5.835 0.085 6.005 0.555 ;
      RECT 6.175 0.255 8.185 0.475 ;
      RECT 6.175 2.215 8.185 2.635 ;
      RECT 7.935 0.475 8.185 0.725 ;
      RECT 7.935 0.725 9.025 0.905 ;
      RECT 8.355 0.085 8.525 0.555 ;
      RECT 8.355 2.045 8.525 2.465 ;
      RECT 8.435 1.445 9.405 1.615 ;
      RECT 8.435 1.615 8.605 1.785 ;
      RECT 8.695 0.255 9.025 0.725 ;
      RECT 8.775 1.795 8.945 2.635 ;
      RECT 9.155 1.615 9.405 2.465 ;
      RECT 9.195 0.085 9.365 0.905 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__a221oi_4
MACRO sky130_fd_sc_hd__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.675 2.2 1.075 ;
        RECT 1.945 1.075 2.275 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 0.995 2.755 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.695 1.285 ;
        RECT 1.415 0.675 1.695 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.075 1.055 1.285 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.285 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.767000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.17 0.255 0.345 0.735 ;
        RECT 0.17 0.735 1.235 0.905 ;
        RECT 0.175 1.455 2.3 1.495 ;
        RECT 0.175 1.495 3.135 1.625 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 1.065 0.255 2.58 0.505 ;
        RECT 1.065 0.505 1.235 0.735 ;
        RECT 2.15 1.625 3.135 1.665 ;
        RECT 2.38 0.505 2.58 0.655 ;
        RECT 2.38 0.655 3.135 0.825 ;
        RECT 2.925 0.825 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.515 1.795 0.765 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.025 1.835 ;
      RECT 1.015 1.835 2.625 2.045 ;
      RECT 1.015 2.045 1.24 2.125 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 1.875 2.215 2.205 2.635 ;
      RECT 2.375 2.045 2.625 2.465 ;
      RECT 2.75 0.085 3.08 0.485 ;
      RECT 2.795 1.875 3.125 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a221oi_1
MACRO sky130_fd_sc_hd__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 4.48 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435 1.075 3.765 1.445 ;
        RECT 3.435 1.445 4.82 1.615 ;
        RECT 4.65 1.075 5.435 1.275 ;
        RECT 4.65 1.275 4.82 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 2.765 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 2.04 1.445 ;
        RECT 1.505 1.445 3.265 1.615 ;
        RECT 2.935 1.075 3.265 1.445 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.42 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.305 0.855 0.725 ;
        RECT 0.525 0.725 4.395 0.865 ;
        RECT 0.605 0.865 4.395 0.905 ;
        RECT 0.605 0.905 0.855 2.125 ;
        RECT 2.285 0.645 2.635 0.725 ;
        RECT 4.065 0.645 4.395 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.09 1.795 0.435 2.295 ;
      RECT 0.09 2.295 1.275 2.465 ;
      RECT 0.105 0.085 0.355 0.895 ;
      RECT 1.025 0.085 1.715 0.555 ;
      RECT 1.025 1.495 1.275 1.785 ;
      RECT 1.025 1.785 3.015 1.955 ;
      RECT 1.025 1.955 1.275 2.295 ;
      RECT 1.505 2.125 1.755 2.295 ;
      RECT 1.505 2.295 3.475 2.465 ;
      RECT 1.885 0.255 3.055 0.475 ;
      RECT 1.925 1.955 2.175 2.125 ;
      RECT 2.345 2.125 2.595 2.295 ;
      RECT 2.765 1.955 3.015 2.125 ;
      RECT 3.225 1.785 5.195 1.955 ;
      RECT 3.225 1.955 3.475 2.295 ;
      RECT 3.27 0.085 3.44 0.555 ;
      RECT 3.645 0.255 4.815 0.475 ;
      RECT 3.685 2.125 3.935 2.635 ;
      RECT 4.105 1.955 4.355 2.465 ;
      RECT 4.525 2.125 4.775 2.635 ;
      RECT 4.565 0.475 4.815 0.905 ;
      RECT 4.985 0.085 5.155 0.905 ;
      RECT 4.99 1.455 5.195 1.785 ;
      RECT 4.99 1.955 5.195 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__a221oi_2
MACRO sky130_fd_sc_hd__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.745 0.41 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.125 2.29 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 0.305 2.22 0.765 ;
        RECT 2.01 0.765 2.42 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.795 3.16 2.465 ;
        RECT 2.915 0.255 3.16 0.715 ;
        RECT 2.99 0.715 3.16 0.925 ;
        RECT 2.99 0.925 3.595 1.445 ;
        RECT 2.99 1.445 3.16 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.085 0.355 0.575 ;
      RECT 0.085 1.575 0.4 2.635 ;
      RECT 0.58 0.305 0.855 1.015 ;
      RECT 0.58 1.015 1.415 1.245 ;
      RECT 0.58 1.245 0.855 1.905 ;
      RECT 1.03 2.13 1.645 2.635 ;
      RECT 1.05 1.425 2.82 1.595 ;
      RECT 1.05 1.595 1.285 1.96 ;
      RECT 1.055 0.305 1.84 0.57 ;
      RECT 1.455 1.765 1.785 1.955 ;
      RECT 1.455 1.955 1.645 2.13 ;
      RECT 1.585 0.57 1.84 1.425 ;
      RECT 2.01 1.595 2.2 1.89 ;
      RECT 2.41 0.085 2.74 0.58 ;
      RECT 2.46 1.79 2.675 2.635 ;
      RECT 2.59 0.995 2.82 1.425 ;
      RECT 3.33 0.085 3.595 0.745 ;
      RECT 3.33 1.625 3.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__and3b_2
MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715 0.615 3.995 1.705 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.02 0.725 1.235 1.34 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.715 1.34 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.535 3.535 1.705 ;
        RECT 2.285 0.515 2.475 0.615 ;
        RECT 2.285 0.615 3.535 0.845 ;
        RECT 3.145 0.255 3.335 0.615 ;
        RECT 3.27 0.845 3.535 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.15 0.255 0.635 0.355 ;
      RECT 0.15 0.355 1.6 0.545 ;
      RECT 0.15 0.545 0.635 0.805 ;
      RECT 0.15 0.805 0.37 1.495 ;
      RECT 0.15 1.495 0.51 2.165 ;
      RECT 0.54 0.995 0.85 1.325 ;
      RECT 0.68 1.325 0.85 1.875 ;
      RECT 0.68 1.875 4.445 2.105 ;
      RECT 0.73 2.275 1.18 2.635 ;
      RECT 1.28 1.525 2.055 1.695 ;
      RECT 1.42 0.545 1.6 0.615 ;
      RECT 1.42 0.615 2.115 0.805 ;
      RECT 1.745 2.275 2.075 2.635 ;
      RECT 1.78 0.085 2.11 0.445 ;
      RECT 1.885 0.805 2.115 1.02 ;
      RECT 1.885 1.02 3.1 1.355 ;
      RECT 1.885 1.355 2.055 1.525 ;
      RECT 2.645 0.085 2.975 0.445 ;
      RECT 2.645 2.275 2.98 2.635 ;
      RECT 3.505 0.085 3.835 0.445 ;
      RECT 3.505 2.275 3.835 2.635 ;
      RECT 4.165 0.425 4.445 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__and3b_4
MACRO sky130_fd_sc_hd__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.955 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.79 2.125 2.265 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.305 2.185 0.725 ;
        RECT 1.985 0.725 2.395 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.86 1.765 3.135 2.465 ;
        RECT 2.875 0.255 3.135 0.735 ;
        RECT 2.965 0.735 3.135 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.085 0.085 0.345 0.905 ;
      RECT 0.085 2.125 0.345 2.635 ;
      RECT 0.515 0.485 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.39 1.245 ;
      RECT 0.595 1.245 0.765 2.465 ;
      RECT 1.005 1.425 2.795 1.595 ;
      RECT 1.005 1.595 1.255 1.96 ;
      RECT 1.005 2.13 1.62 2.635 ;
      RECT 1.025 0.305 1.815 0.57 ;
      RECT 1.425 1.765 1.755 1.955 ;
      RECT 1.425 1.955 1.62 2.13 ;
      RECT 1.56 0.57 1.815 1.425 ;
      RECT 1.975 1.595 2.69 1.89 ;
      RECT 2.375 0.085 2.705 0.545 ;
      RECT 2.435 2.09 2.65 2.635 ;
      RECT 2.565 0.995 2.795 1.425 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__and3b_1
MACRO sky130_fd_sc_hd__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.81 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 1.075 1.75 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.735 ;
        RECT 0.535 0.735 2.135 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.375 1.445 2.135 1.665 ;
        RECT 1.375 1.665 1.705 2.125 ;
        RECT 1.92 0.905 2.135 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.09 1.455 1.205 1.665 ;
      RECT 0.09 1.665 0.365 2.465 ;
      RECT 0.535 1.835 0.865 2.635 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.035 1.665 1.205 2.295 ;
      RECT 1.035 2.295 2.175 2.465 ;
      RECT 1.875 0.085 2.165 0.555 ;
      RECT 1.875 1.835 2.175 2.295 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nor2_2
MACRO sky130_fd_sc_hd__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.8 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.12 1.075 3.485 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 4.055 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 1.445 4.055 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
        RECT 3.655 0.905 4.055 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.09 1.455 2.125 1.665 ;
      RECT 0.09 1.665 0.365 2.465 ;
      RECT 0.535 1.835 0.865 2.635 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.375 1.835 1.625 2.635 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.89 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 3.475 1.915 3.89 2.295 ;
      RECT 3.555 0.085 3.84 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__nor2_4
MACRO sky130_fd_sc_hd__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.075 1.295 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.775 1.665 ;
        RECT 0.095 1.665 0.425 2.45 ;
        RECT 0.515 0.255 0.845 0.895 ;
        RECT 0.605 0.895 0.775 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.105 0.085 0.345 0.895 ;
      RECT 0.955 1.495 1.285 2.635 ;
      RECT 1.015 0.085 1.285 0.895 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__nor2_1
MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 3.53 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.8 1.075 6.54 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 7.275 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 3.935 1.445 7.275 1.615 ;
        RECT 3.935 1.615 4.185 2.125 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 4.775 1.615 5.025 2.125 ;
        RECT 5.575 0.255 5.905 0.725 ;
        RECT 5.615 1.615 5.865 2.125 ;
        RECT 6.415 0.255 6.745 0.725 ;
        RECT 6.455 1.615 6.705 2.125 ;
        RECT 6.71 0.905 7.275 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.09 1.455 3.765 1.665 ;
      RECT 0.09 1.665 0.405 2.465 ;
      RECT 0.575 1.835 0.825 2.635 ;
      RECT 0.995 1.665 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.835 1.665 2.635 ;
      RECT 1.835 1.665 2.085 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.255 1.835 2.505 2.635 ;
      RECT 2.675 1.665 2.925 2.465 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 3.095 1.835 3.345 2.635 ;
      RECT 3.515 1.665 3.765 2.295 ;
      RECT 3.515 2.295 7.125 2.465 ;
      RECT 3.555 0.085 3.725 0.555 ;
      RECT 4.355 1.785 4.605 2.295 ;
      RECT 4.395 0.085 4.565 0.555 ;
      RECT 5.195 1.785 5.445 2.295 ;
      RECT 5.235 0.085 5.405 0.555 ;
      RECT 6.035 1.785 6.285 2.295 ;
      RECT 6.075 0.085 6.245 0.555 ;
      RECT 6.875 1.785 7.125 2.295 ;
      RECT 6.915 0.085 7.205 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__nor2_8
MACRO sky130_fd_sc_hd__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425 0.995 1.755 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.732000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.13 1.495 2.675 1.665 ;
        RECT 1.13 1.665 1.46 2.465 ;
        RECT 2.085 0.255 2.675 0.485 ;
        RECT 2.085 1.665 2.675 2.465 ;
        RECT 2.385 0.485 2.675 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.085 0.445 0.51 0.655 ;
      RECT 0.085 0.655 2.215 0.825 ;
      RECT 0.085 0.825 0.255 1.595 ;
      RECT 0.085 1.595 0.51 1.925 ;
      RECT 0.71 0.085 1.04 0.485 ;
      RECT 0.71 1.495 0.96 2.635 ;
      RECT 1.63 1.835 1.915 2.635 ;
      RECT 2.045 0.825 2.215 1.325 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__nand3b_1
MACRO sky130_fd_sc_hd__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.27 1.075 4.48 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 6.5 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.965 0.905 ;
        RECT 1.455 1.445 6.505 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 3.465 2.005 ;
        RECT 2.295 2.005 2.625 2.465 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 2.795 1.075 3.1 1.445 ;
        RECT 3.135 2.005 3.465 2.465 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.285 0.905 ;
      RECT 0.085 0.905 0.26 1.445 ;
      RECT 0.085 1.445 0.425 2.465 ;
      RECT 0.595 0.085 0.845 0.545 ;
      RECT 0.595 1.445 1.285 2.635 ;
      RECT 1.005 0.905 1.285 1.075 ;
      RECT 1.005 1.075 2.625 1.275 ;
      RECT 1.035 0.255 4.725 0.465 ;
      RECT 1.955 1.835 2.125 2.635 ;
      RECT 2.795 2.175 2.965 2.635 ;
      RECT 3.135 0.635 4.725 0.715 ;
      RECT 3.135 0.715 6.505 0.905 ;
      RECT 3.635 1.835 3.805 2.635 ;
      RECT 4.475 1.835 5.165 2.635 ;
      RECT 4.915 0.085 5.165 0.545 ;
      RECT 5.335 0.255 5.665 0.715 ;
      RECT 5.835 0.085 6.005 0.545 ;
      RECT 5.835 1.835 6.005 2.635 ;
      RECT 6.175 0.255 6.505 0.715 ;
      RECT 6.675 0.085 7.005 0.905 ;
      RECT 6.675 1.445 7.005 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__nand3b_4
MACRO sky130_fd_sc_hd__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.075 3.14 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.74 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.785 4.05 1.955 ;
        RECT 1.06 1.955 2.23 2.005 ;
        RECT 1.06 2.005 1.39 2.465 ;
        RECT 1.9 2.005 2.23 2.465 ;
        RECT 3.26 0.635 4.05 0.905 ;
        RECT 3.26 1.955 4.05 2.005 ;
        RECT 3.26 2.005 3.51 2.465 ;
        RECT 3.85 0.905 4.05 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.09 0.255 0.41 0.655 ;
      RECT 0.09 0.655 0.26 1.445 ;
      RECT 0.09 1.445 3.65 1.615 ;
      RECT 0.09 1.615 0.26 2.065 ;
      RECT 0.09 2.065 0.41 2.465 ;
      RECT 0.58 0.085 0.89 0.905 ;
      RECT 0.58 1.835 0.89 2.635 ;
      RECT 1.06 0.255 1.39 0.715 ;
      RECT 1.06 0.715 2.75 0.905 ;
      RECT 1.56 0.085 1.81 0.545 ;
      RECT 1.56 2.175 1.73 2.635 ;
      RECT 2 0.255 4.05 0.465 ;
      RECT 2 0.635 2.75 0.715 ;
      RECT 2.4 2.175 2.65 2.635 ;
      RECT 2.84 2.175 3.09 2.635 ;
      RECT 2.92 0.465 3.09 0.905 ;
      RECT 3.32 1.075 3.65 1.445 ;
      RECT 3.76 2.175 4.05 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__nand3b_2
MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.45 1.675 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.42 1.8 1.695 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 0.42 2.295 1.695 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 0.665 2.825 1.695 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255 0.295 3.59 0.34 ;
        RECT 3.255 0.34 3.595 0.805 ;
        RECT 3.335 1.495 3.595 2.465 ;
        RECT 3.425 0.805 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.17 0.255 0.345 0.655 ;
      RECT 0.17 0.655 0.8 0.825 ;
      RECT 0.17 1.845 0.8 2.015 ;
      RECT 0.17 2.015 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.195 0.845 2.635 ;
      RECT 0.63 0.825 0.8 0.995 ;
      RECT 0.63 0.995 0.98 1.325 ;
      RECT 0.63 1.325 0.8 1.845 ;
      RECT 1.09 0.255 1.32 0.585 ;
      RECT 1.15 0.585 1.32 1.875 ;
      RECT 1.15 1.875 3.165 2.045 ;
      RECT 1.15 2.045 1.32 2.465 ;
      RECT 1.555 2.225 2.225 2.635 ;
      RECT 2.44 2.045 2.61 2.465 ;
      RECT 2.755 0.085 3.085 0.465 ;
      RECT 2.81 2.225 3.14 2.635 ;
      RECT 2.995 0.995 3.255 1.325 ;
      RECT 2.995 1.325 3.165 1.875 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__and4b_1
MACRO sky130_fd_sc_hd__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.44 0.765 0.79 1.635 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.735 4.145 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345 0.755 3.555 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.085 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 0.65 2.08 0.82 ;
        RECT 0.98 0.82 1.26 1.545 ;
        RECT 0.98 1.545 2.16 1.715 ;
        RECT 1.07 0.255 1.24 0.65 ;
        RECT 1.91 0.255 2.08 0.65 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.26 1.915 ;
      RECT 0.085 1.915 4.9 2.085 ;
      RECT 0.085 2.085 0.345 2.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 0.57 0.085 0.9 0.47 ;
      RECT 1.41 0.085 1.74 0.47 ;
      RECT 1.41 2.255 1.74 2.635 ;
      RECT 1.44 1.075 2.55 1.245 ;
      RECT 2.25 2.255 2.58 2.635 ;
      RECT 2.285 0.085 2.615 0.445 ;
      RECT 2.38 0.615 2.965 0.785 ;
      RECT 2.38 0.785 2.55 1.075 ;
      RECT 2.38 1.245 2.55 1.545 ;
      RECT 2.38 1.545 4.545 1.715 ;
      RECT 2.795 0.3 4.965 0.47 ;
      RECT 2.795 0.47 2.965 0.615 ;
      RECT 3.475 2.255 3.805 2.635 ;
      RECT 4.39 0.47 4.965 0.81 ;
      RECT 4.635 2.255 4.965 2.635 ;
      RECT 4.73 0.995 4.9 1.915 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__and4b_4
MACRO sky130_fd_sc_hd__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.74 0.335 1.63 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.42 1.745 1.745 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 0.42 2.275 1.695 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.645 2.775 1.615 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.503250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 0.255 3.545 0.64 ;
        RECT 3.26 0.64 4.055 0.825 ;
        RECT 3.34 1.535 4.055 1.745 ;
        RECT 3.34 1.745 3.545 2.465 ;
        RECT 3.425 0.825 4.055 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.095 0.085 0.425 0.465 ;
      RECT 0.175 1.83 0.805 2 ;
      RECT 0.175 2 0.345 2.465 ;
      RECT 0.515 2.195 0.845 2.635 ;
      RECT 0.595 0.255 0.805 0.585 ;
      RECT 0.635 0.585 0.805 0.995 ;
      RECT 0.635 0.995 0.975 1.325 ;
      RECT 0.635 1.325 0.805 1.83 ;
      RECT 1.015 1.66 1.315 1.915 ;
      RECT 1.015 1.915 3.165 1.965 ;
      RECT 1.015 1.965 2.61 2.085 ;
      RECT 1.015 2.085 1.185 2.465 ;
      RECT 1.095 0.255 1.315 0.585 ;
      RECT 1.145 0.585 1.315 1.66 ;
      RECT 1.555 2.255 2.225 2.635 ;
      RECT 2.44 1.795 3.165 1.915 ;
      RECT 2.44 2.085 2.61 2.465 ;
      RECT 2.76 0.085 3.09 0.465 ;
      RECT 2.84 2.195 3.17 2.635 ;
      RECT 2.995 0.995 3.255 1.325 ;
      RECT 2.995 1.325 3.165 1.795 ;
      RECT 3.715 0.085 4.05 0.465 ;
      RECT 3.715 1.915 4.05 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__and4b_2
MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.315 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.085 1.315 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 1.835 2.17 2.005 ;
        RECT 1 2.005 1.33 2.465 ;
        RECT 1.42 0.255 2.17 0.545 ;
        RECT 1.8 0.545 2.17 1.835 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.09 0.525 0.36 0.735 ;
      RECT 0.09 0.735 1.425 0.905 ;
      RECT 0.09 1.495 1.425 1.665 ;
      RECT 0.09 1.665 0.37 1.825 ;
      RECT 0.58 0.085 0.91 0.545 ;
      RECT 0.58 1.835 0.83 2.635 ;
      RECT 1.255 0.905 1.425 1.075 ;
      RECT 1.255 1.075 1.63 1.325 ;
      RECT 1.255 1.325 1.425 1.495 ;
      RECT 1.5 2.175 1.715 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nand2b_1
MACRO sky130_fd_sc_hd__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.075 4.94 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.64 0.905 ;
        RECT 1.455 1.445 4.32 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.64 2.465 ;
        RECT 2.375 0.905 2.64 1.445 ;
        RECT 3.15 1.665 3.48 2.465 ;
        RECT 3.99 1.665 4.32 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.25 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.06 0.085 ;
      RECT 0 2.635 5.06 2.805 ;
      RECT 0.09 0.255 0.425 0.715 ;
      RECT 0.09 0.715 0.78 0.905 ;
      RECT 0.09 1.445 0.78 1.665 ;
      RECT 0.09 1.665 0.425 2.465 ;
      RECT 0.595 0.085 0.79 0.545 ;
      RECT 0.595 1.835 1.285 2.635 ;
      RECT 0.61 0.905 0.78 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.78 1.445 ;
      RECT 0.97 1.445 1.285 1.835 ;
      RECT 1.035 0.255 3.06 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 1.955 1.835 2.125 2.635 ;
      RECT 2.81 0.465 3.06 0.715 ;
      RECT 2.81 0.715 4.85 0.905 ;
      RECT 2.81 1.835 2.98 2.635 ;
      RECT 3.23 0.085 3.4 0.545 ;
      RECT 3.57 0.255 3.9 0.715 ;
      RECT 3.65 1.835 3.82 2.635 ;
      RECT 4.07 0.085 4.31 0.545 ;
      RECT 4.52 0.255 4.85 0.715 ;
      RECT 4.52 1.495 4.85 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
  END
END sky130_fd_sc_hd__nand2b_4
MACRO sky130_fd_sc_hd__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 0.995 0.8 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.135 1.275 ;
        RECT 1.99 1.275 2.18 1.655 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.775500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.835 2.635 2.005 ;
        RECT 1.035 2.005 1.365 2.465 ;
        RECT 1.525 0.635 1.855 0.805 ;
        RECT 1.53 0.805 1.855 0.905 ;
        RECT 1.53 0.905 1.81 1.835 ;
        RECT 2.28 2.005 2.635 2.465 ;
        RECT 2.36 1.495 2.635 1.835 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.11 0.51 0.345 0.84 ;
      RECT 0.11 0.84 0.28 1.495 ;
      RECT 0.11 1.495 1.36 1.665 ;
      RECT 0.11 1.665 0.41 1.86 ;
      RECT 0.515 0.085 0.845 0.825 ;
      RECT 0.58 1.835 0.835 2.635 ;
      RECT 1.03 1.075 1.36 1.495 ;
      RECT 1.08 0.255 2.275 0.465 ;
      RECT 1.08 0.465 1.355 0.905 ;
      RECT 1.535 2.175 2.11 2.635 ;
      RECT 2.025 0.465 2.275 0.695 ;
      RECT 2.025 0.695 3.135 0.905 ;
      RECT 2.445 0.085 2.615 0.525 ;
      RECT 2.785 0.255 3.135 0.695 ;
      RECT 2.805 1.495 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__nand2b_2
MACRO sky130_fd_sc_hd__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.075 1.055 1.325 ;
        RECT 0.595 1.325 0.83 2.05 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305 0.265 2.635 0.735 ;
        RECT 2.305 0.735 4.055 0.905 ;
        RECT 2.345 1.455 4.055 1.625 ;
        RECT 2.345 1.625 2.595 2.465 ;
        RECT 3.145 0.265 3.475 0.735 ;
        RECT 3.185 1.625 3.435 2.465 ;
        RECT 3.765 0.905 4.055 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.255 0.425 0.725 ;
      RECT 0.085 0.725 2.09 0.905 ;
      RECT 0.085 1.495 0.425 2.295 ;
      RECT 0.085 2.295 1.265 2.465 ;
      RECT 0.595 0.085 0.765 0.555 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 1 1.495 2.09 1.665 ;
      RECT 1 1.665 1.265 2.295 ;
      RECT 1.435 0.085 2.135 0.555 ;
      RECT 1.435 1.835 2.135 2.635 ;
      RECT 1.87 0.905 2.09 1.075 ;
      RECT 1.87 1.075 3.595 1.245 ;
      RECT 1.87 1.245 2.09 1.495 ;
      RECT 2.765 1.795 3.015 2.635 ;
      RECT 2.805 0.085 2.975 0.555 ;
      RECT 3.605 1.795 3.855 2.635 ;
      RECT 3.645 0.085 3.815 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__or3_4
MACRO sky130_fd_sc_hd__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.43 1.325 ;
        RECT 0.605 1.325 0.83 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.28 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.435 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 0.415 2.215 0.76 ;
        RECT 1.94 1.495 2.215 2.465 ;
        RECT 2.045 0.76 2.215 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.105 0.305 0.36 0.655 ;
      RECT 0.105 0.655 1.77 0.825 ;
      RECT 0.105 1.495 0.435 1.785 ;
      RECT 0.105 1.785 1.27 1.955 ;
      RECT 0.53 0.085 0.86 0.485 ;
      RECT 1.03 0.305 1.2 0.655 ;
      RECT 1.1 1.495 1.77 1.665 ;
      RECT 1.1 1.665 1.27 1.785 ;
      RECT 1.37 0.085 1.75 0.485 ;
      RECT 1.45 1.835 1.73 2.635 ;
      RECT 1.6 0.825 1.77 0.995 ;
      RECT 1.6 0.995 1.875 1.325 ;
      RECT 1.6 1.325 1.77 1.495 ;
      RECT 2.385 0.085 2.675 0.915 ;
      RECT 2.385 1.43 2.675 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__or3_2
MACRO sky130_fd_sc_hd__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.6 0.995 1.425 1.325 ;
        RECT 0.6 1.325 0.795 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.275 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.43 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.415 2.21 0.76 ;
        RECT 1.935 1.495 2.21 2.465 ;
        RECT 2.04 0.76 2.21 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.1 0.305 0.355 0.655 ;
      RECT 0.1 0.655 1.765 0.825 ;
      RECT 0.105 1.495 0.43 1.785 ;
      RECT 0.105 1.785 1.275 1.955 ;
      RECT 0.525 0.085 0.855 0.485 ;
      RECT 1.025 0.305 1.195 0.655 ;
      RECT 1.105 1.495 1.765 1.665 ;
      RECT 1.105 1.665 1.275 1.785 ;
      RECT 1.365 0.085 1.745 0.485 ;
      RECT 1.445 1.835 1.725 2.635 ;
      RECT 1.595 0.825 1.765 0.995 ;
      RECT 1.595 0.995 1.87 1.325 ;
      RECT 1.595 1.325 1.765 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__or3_1
MACRO sky130_fd_sc_hd__dlymetal6s2s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s2s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.57 1.7 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 0.255 1.67 0.825 ;
        RECT 1.245 1.495 2.15 1.675 ;
        RECT 1.245 1.675 1.67 2.465 ;
        RECT 1.32 0.825 1.67 0.995 ;
        RECT 1.32 0.995 2.15 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.12 -0.085 0.29 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.255 0.52 0.655 ;
      RECT 0.085 0.655 1.075 0.825 ;
      RECT 0.085 1.87 1.075 2.04 ;
      RECT 0.085 2.04 0.52 2.465 ;
      RECT 0.69 0.085 1.075 0.485 ;
      RECT 0.69 2.21 1.075 2.635 ;
      RECT 0.74 0.825 1.075 0.995 ;
      RECT 0.74 0.995 1.15 1.325 ;
      RECT 0.74 1.325 1.075 1.87 ;
      RECT 1.84 1.845 2.67 2.04 ;
      RECT 1.84 2.04 2.115 2.465 ;
      RECT 1.86 0.255 2.115 0.655 ;
      RECT 1.86 0.655 2.67 0.825 ;
      RECT 2.285 0.085 2.67 0.485 ;
      RECT 2.285 2.21 2.67 2.635 ;
      RECT 2.32 0.825 2.67 0.995 ;
      RECT 2.32 0.995 2.745 1.325 ;
      RECT 2.32 1.325 2.67 1.845 ;
      RECT 2.84 0.255 3.085 0.825 ;
      RECT 2.84 1.495 3.565 1.675 ;
      RECT 2.84 1.675 3.085 2.465 ;
      RECT 2.915 0.825 3.085 0.995 ;
      RECT 2.915 0.995 3.565 1.495 ;
      RECT 3.275 0.255 3.53 0.655 ;
      RECT 3.275 0.655 4.085 0.825 ;
      RECT 3.275 1.845 4.085 2.04 ;
      RECT 3.275 2.04 3.53 2.465 ;
      RECT 3.7 0.085 4.085 0.485 ;
      RECT 3.7 2.21 4.085 2.635 ;
      RECT 3.735 0.825 4.085 0.995 ;
      RECT 3.735 0.995 4.16 1.325 ;
      RECT 3.735 1.325 4.085 1.845 ;
      RECT 4.255 0.255 4.515 0.825 ;
      RECT 4.255 1.495 4.515 2.465 ;
      RECT 4.33 0.825 4.515 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__dlymetal6s2s_1
MACRO sky130_fd_sc_hd__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.375000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.375000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_1
MACRO sky130_fd_sc_hd__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.835000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.775000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.835000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_2
MACRO sky130_fd_sc_hd__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.18 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 4.07 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 1.075 5.705 1.285 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875 1.075 7.295 1.285 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 7.735 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 4.415 0.255 4.745 0.725 ;
        RECT 5.255 0.255 5.585 0.725 ;
        RECT 6.095 0.255 6.425 0.725 ;
        RECT 6.135 1.455 7.735 1.625 ;
        RECT 6.135 1.625 6.385 2.125 ;
        RECT 6.935 0.255 7.265 0.725 ;
        RECT 6.975 1.625 7.225 2.125 ;
        RECT 7.465 0.905 7.735 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.01 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.82 0.085 ;
      RECT 0 2.635 7.82 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.09 1.455 2.085 1.625 ;
      RECT 0.09 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.795 1.665 2.635 ;
      RECT 1.835 1.625 2.085 2.295 ;
      RECT 1.835 2.295 3.82 2.465 ;
      RECT 1.875 0.085 2.045 0.555 ;
      RECT 2.255 1.455 5.545 1.625 ;
      RECT 2.255 1.625 2.505 2.125 ;
      RECT 2.675 1.795 2.925 2.295 ;
      RECT 2.715 0.085 2.885 0.555 ;
      RECT 3.095 1.625 3.345 2.125 ;
      RECT 3.515 1.795 3.82 2.295 ;
      RECT 3.555 0.085 4.245 0.555 ;
      RECT 4.005 1.795 4.285 2.295 ;
      RECT 4.005 2.295 7.645 2.465 ;
      RECT 4.455 1.625 4.705 2.125 ;
      RECT 4.875 1.795 5.125 2.295 ;
      RECT 4.915 0.085 5.085 0.555 ;
      RECT 5.295 1.625 5.545 2.125 ;
      RECT 5.715 1.795 5.965 2.295 ;
      RECT 5.755 0.085 5.925 0.555 ;
      RECT 6.555 1.795 6.805 2.295 ;
      RECT 6.595 0.085 6.765 0.555 ;
      RECT 7.395 1.795 7.645 2.295 ;
      RECT 7.435 0.085 7.605 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
  END
END sky130_fd_sc_hd__nor4_4
MACRO sky130_fd_sc_hd__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.2 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 1.94 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 3.105 1.285 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.34 1.075 3.925 1.285 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 4.515 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.615 0.255 3.945 0.725 ;
        RECT 3.655 1.455 4.515 1.625 ;
        RECT 3.655 1.625 3.905 2.125 ;
        RECT 4.18 0.905 4.515 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.065 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 1.875 0.085 2.605 0.555 ;
      RECT 2.395 1.455 3.485 1.625 ;
      RECT 2.395 1.625 2.645 2.125 ;
      RECT 2.815 1.795 3.065 2.295 ;
      RECT 3.235 1.625 3.485 2.295 ;
      RECT 3.235 2.295 4.325 2.465 ;
      RECT 3.275 0.085 3.445 0.555 ;
      RECT 4.075 1.795 4.325 2.295 ;
      RECT 4.115 0.085 4.405 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__nor4_2
MACRO sky130_fd_sc_hd__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.655 2.215 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 1.075 1.695 1.245 ;
        RECT 1.455 1.245 1.695 2.45 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 0.995 1.075 1.415 ;
        RECT 0.845 1.415 1.285 1.615 ;
        RECT 1.03 1.615 1.285 2.45 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.335 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.672750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.495 0.675 1.665 ;
        RECT 0.09 1.665 0.425 2.45 ;
        RECT 0.505 0.645 0.86 0.655 ;
        RECT 0.505 0.655 1.705 0.825 ;
        RECT 0.505 0.825 0.675 1.495 ;
        RECT 0.595 0.385 0.86 0.645 ;
        RECT 1.535 0.385 1.705 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.49 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.3 0.085 ;
      RECT 0 2.635 2.3 2.805 ;
      RECT 0.085 0.085 0.345 0.575 ;
      RECT 1.035 0.085 1.365 0.485 ;
      RECT 1.875 0.085 2.205 0.485 ;
      RECT 1.955 1.835 2.215 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
  END
END sky130_fd_sc_hd__nor4_1
MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 1.055 5.47 1.36 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265 1.055 4.97 1.36 ;
        RECT 4.68 1.36 4.97 1.53 ;
        RECT 4.68 1.53 6.355 1.7 ;
        RECT 5.64 1.055 6.355 1.53 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765 1.055 4.095 1.36 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 1.055 3.575 1.355 ;
        RECT 2.78 1.355 3.15 1.695 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 1.765 0.885 ;
        RECT 0.085 0.885 0.735 1.46 ;
        RECT 0.085 1.46 1.75 1.665 ;
        RECT 0.68 0.255 0.895 0.655 ;
        RECT 0.68 0.655 1.765 0.715 ;
        RECT 0.68 1.665 0.895 2.465 ;
        RECT 1.565 0.255 1.765 0.655 ;
        RECT 1.565 1.665 1.75 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.085 0.085 0.51 0.545 ;
      RECT 0.085 1.835 0.51 2.635 ;
      RECT 0.905 1.055 2.61 1.29 ;
      RECT 1.065 0.085 1.395 0.485 ;
      RECT 1.065 1.835 1.395 2.635 ;
      RECT 1.92 1.46 2.25 2.635 ;
      RECT 1.935 0.085 2.25 0.885 ;
      RECT 2.44 0.255 3.57 0.465 ;
      RECT 2.44 0.635 3.21 0.885 ;
      RECT 2.44 0.885 2.61 1.055 ;
      RECT 2.44 1.29 2.61 1.87 ;
      RECT 2.44 1.87 4.09 2.07 ;
      RECT 2.44 2.07 2.61 2.465 ;
      RECT 2.78 2.24 3.11 2.635 ;
      RECT 3.32 1.53 4.51 1.7 ;
      RECT 3.38 0.465 3.57 0.635 ;
      RECT 3.38 0.635 6.355 0.885 ;
      RECT 3.76 0.085 4.09 0.445 ;
      RECT 3.76 2.07 4.09 2.465 ;
      RECT 4.26 0.255 4.43 0.635 ;
      RECT 4.26 1.7 4.51 2.465 ;
      RECT 4.6 0.085 4.93 0.445 ;
      RECT 4.68 1.87 5.72 2.07 ;
      RECT 4.68 2.07 4.85 2.465 ;
      RECT 5.02 2.24 5.35 2.635 ;
      RECT 5.1 0.255 5.27 0.635 ;
      RECT 5.44 0.085 5.77 0.445 ;
      RECT 5.52 2.07 5.72 2.465 ;
      RECT 5.89 1.87 6.355 2.465 ;
      RECT 5.94 0.255 6.355 0.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.125 4.455 2.295 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.125 6.295 2.295 ;
      RECT 6.125 2.635 6.295 2.805 ;
    LAYER met1 ;
      RECT 4.225 2.095 4.515 2.14 ;
      RECT 4.225 2.14 6.355 2.28 ;
      RECT 4.225 2.28 4.515 2.325 ;
      RECT 6.065 2.095 6.355 2.14 ;
      RECT 6.065 2.28 6.355 2.325 ;
  END
END sky130_fd_sc_hd__o31a_4
MACRO sky130_fd_sc_hd__o31a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.995 1.76 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.995 2.19 1.325 ;
        RECT 1.99 1.325 2.19 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 0.995 2.64 2.125 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.255 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.577500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.86 1.295 ;
        RECT 0.55 0.265 0.99 0.825 ;
        RECT 0.55 0.825 0.86 1.075 ;
        RECT 0.55 1.295 0.86 1.835 ;
        RECT 0.55 1.835 0.99 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.085 0.085 0.38 0.905 ;
      RECT 0.085 1.465 0.38 2.635 ;
      RECT 1.03 0.995 1.2 1.445 ;
      RECT 1.03 1.445 1.82 1.615 ;
      RECT 1.16 0.085 1.61 0.825 ;
      RECT 1.165 1.785 1.48 2.635 ;
      RECT 1.65 1.615 1.82 2.295 ;
      RECT 1.65 2.295 3.08 2.465 ;
      RECT 1.78 0.255 1.95 0.655 ;
      RECT 1.78 0.655 2.94 0.825 ;
      RECT 2.12 0.085 2.54 0.485 ;
      RECT 2.71 0.255 2.94 0.655 ;
      RECT 2.83 1.495 3.595 1.665 ;
      RECT 2.83 1.665 3.08 2.295 ;
      RECT 3.11 0.255 3.595 0.825 ;
      RECT 3.255 1.835 3.59 2.635 ;
      RECT 3.425 0.825 3.595 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o31a_2
MACRO sky130_fd_sc_hd__o31a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.295 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.995 1.725 1.325 ;
        RECT 1.525 1.325 1.725 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.995 2.175 2.125 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 0.995 2.795 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.594000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.265 0.525 0.825 ;
        RECT 0.085 0.825 0.395 1.835 ;
        RECT 0.085 1.835 0.525 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.565 0.995 0.735 1.445 ;
      RECT 0.565 1.445 1.355 1.615 ;
      RECT 0.695 0.085 1.145 0.825 ;
      RECT 0.7 1.785 1.015 2.635 ;
      RECT 1.185 1.615 1.355 2.295 ;
      RECT 1.185 2.295 2.615 2.465 ;
      RECT 1.315 0.255 1.485 0.655 ;
      RECT 1.315 0.655 2.475 0.825 ;
      RECT 1.655 0.085 2.075 0.485 ;
      RECT 2.245 0.255 2.475 0.655 ;
      RECT 2.365 1.495 3.135 1.665 ;
      RECT 2.365 1.665 2.615 2.295 ;
      RECT 2.645 0.255 3.135 0.825 ;
      RECT 2.795 1.835 3.125 2.635 ;
      RECT 2.965 0.825 3.135 1.495 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o31a_1
MACRO sky130_fd_sc_hd__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.485 0.995 5.845 1.62 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.765 0.78 1.635 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 0.755 3.545 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 0.995 3.08 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 0.65 2.08 0.82 ;
        RECT 0.96 0.82 1.24 1.545 ;
        RECT 0.96 1.545 2.16 1.715 ;
        RECT 1.07 0.255 1.24 0.65 ;
        RECT 1.91 0.255 2.08 0.65 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.17 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.98 0.085 ;
      RECT 0 2.635 5.98 2.805 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.26 1.915 ;
      RECT 0.085 1.915 4.49 2.085 ;
      RECT 0.085 2.085 0.345 2.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 0.57 0.085 0.9 0.47 ;
      RECT 1.41 0.085 1.74 0.47 ;
      RECT 1.41 1.075 2.5 1.245 ;
      RECT 1.41 2.255 1.74 2.635 ;
      RECT 2.25 2.255 2.58 2.635 ;
      RECT 2.27 0.085 2.6 0.445 ;
      RECT 2.33 0.615 2.94 0.785 ;
      RECT 2.33 0.785 2.5 1.075 ;
      RECT 2.33 1.245 2.5 1.545 ;
      RECT 2.33 1.545 4.15 1.715 ;
      RECT 2.77 0.3 4.61 0.47 ;
      RECT 2.77 0.47 2.94 0.615 ;
      RECT 3.33 2.255 3.66 2.635 ;
      RECT 3.73 0.995 3.9 1.155 ;
      RECT 3.73 1.155 4.49 1.325 ;
      RECT 4.255 0.47 4.61 0.81 ;
      RECT 4.32 1.325 4.49 1.915 ;
      RECT 4.36 2.255 5.37 2.635 ;
      RECT 4.95 0.655 5.805 0.825 ;
      RECT 4.95 0.825 5.12 1.915 ;
      RECT 4.95 1.915 5.805 2.085 ;
      RECT 4.975 0.085 5.305 0.465 ;
      RECT 5.635 0.255 5.805 0.655 ;
      RECT 5.635 2.085 5.805 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
  END
END sky130_fd_sc_hd__and4bb_4
MACRO sky130_fd_sc_hd__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.625 0.775 1.955 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.765 0.815 0.945 ;
        RECT 0.605 0.945 1.225 1.115 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.415 3.08 0.995 ;
        RECT 2.895 0.995 3.125 1.325 ;
        RECT 2.895 1.325 3.08 1.635 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.42 3.545 0.995 ;
        RECT 3.35 0.995 3.605 1.325 ;
        RECT 3.35 1.325 3.545 1.635 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.425400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255 0.255 4.515 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.285 ;
      RECT 0.085 1.285 1.215 1.455 ;
      RECT 0.085 1.455 0.255 2.135 ;
      RECT 0.085 2.135 0.345 2.465 ;
      RECT 0.655 0.085 0.985 0.465 ;
      RECT 0.655 2.255 0.985 2.635 ;
      RECT 1.045 1.455 1.215 1.575 ;
      RECT 1.045 1.575 1.625 1.745 ;
      RECT 1.165 0.255 2.645 0.425 ;
      RECT 1.165 0.425 1.565 0.755 ;
      RECT 1.225 1.915 1.965 2.085 ;
      RECT 1.225 2.085 1.415 2.465 ;
      RECT 1.395 0.755 1.565 1.235 ;
      RECT 1.395 1.235 1.965 1.405 ;
      RECT 1.665 2.255 1.995 2.635 ;
      RECT 1.755 0.595 2.305 0.925 ;
      RECT 1.795 1.405 1.965 1.915 ;
      RECT 2.135 0.925 2.305 1.915 ;
      RECT 2.135 1.915 4.085 2.085 ;
      RECT 2.205 2.085 2.375 2.465 ;
      RECT 2.475 0.425 2.645 1.325 ;
      RECT 2.57 2.255 2.9 2.635 ;
      RECT 3.16 2.085 3.33 2.465 ;
      RECT 3.755 0.085 4.085 0.465 ;
      RECT 3.755 2.255 4.085 2.635 ;
      RECT 3.915 0.995 4.085 1.915 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__and4bb_1
MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.33 1.635 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.765 4.175 1.305 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.91 0.42 3.175 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.425 3.655 1.405 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.545 1.32 1.715 ;
        RECT 1.015 0.255 1.24 1.545 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.67 0.805 ;
      RECT 0.175 1.885 1.925 2.055 ;
      RECT 0.175 2.055 0.345 2.465 ;
      RECT 0.5 0.805 0.67 1.885 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.255 0.845 2.635 ;
      RECT 1.41 0.085 1.74 0.465 ;
      RECT 1.415 0.635 2.405 0.805 ;
      RECT 1.415 0.805 1.585 1.325 ;
      RECT 1.49 2.255 2.16 2.635 ;
      RECT 1.755 0.995 2.065 1.325 ;
      RECT 1.755 1.325 1.925 1.885 ;
      RECT 2.01 0.255 2.18 0.635 ;
      RECT 2.235 0.805 2.405 1.915 ;
      RECT 2.235 1.915 3.415 2.085 ;
      RECT 2.395 2.085 2.565 2.465 ;
      RECT 2.575 1.4 2.745 1.575 ;
      RECT 2.575 1.575 3.755 1.745 ;
      RECT 2.735 2.255 3.075 2.635 ;
      RECT 3.245 2.085 3.415 2.465 ;
      RECT 3.585 1.745 3.755 1.915 ;
      RECT 3.585 1.915 4.515 2.085 ;
      RECT 3.755 2.255 4.085 2.635 ;
      RECT 3.835 0.085 4.085 0.585 ;
      RECT 4.255 0.255 4.515 0.585 ;
      RECT 4.255 2.085 4.515 2.465 ;
      RECT 4.345 0.585 4.515 1.915 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__and4bb_2
MACRO sky130_fd_sc_hd__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.52 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.01 1.24 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 0.995 3.07 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245 0.995 2.61 1.615 ;
        RECT 2.44 0.425 2.61 0.995 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.515500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 1.785 1.945 1.955 ;
        RECT 1.42 1.955 1.785 2.465 ;
        RECT 1.775 0.255 2.205 0.825 ;
        RECT 1.775 0.825 1.945 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.095 0.085 0.425 0.825 ;
      RECT 0.095 1.805 0.425 2.635 ;
      RECT 0.595 0.255 0.765 0.66 ;
      RECT 0.595 0.66 1.58 0.83 ;
      RECT 0.875 1.445 1.58 1.615 ;
      RECT 0.875 1.615 1.205 2.465 ;
      RECT 0.935 0.085 1.605 0.49 ;
      RECT 1.41 0.83 1.58 1.445 ;
      RECT 1.955 2.235 2.285 2.465 ;
      RECT 2.115 1.785 3.13 1.955 ;
      RECT 2.115 1.955 2.285 2.235 ;
      RECT 2.455 2.135 2.705 2.635 ;
      RECT 2.795 0.085 3.125 0.825 ;
      RECT 2.875 1.955 3.13 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a2bb2oi_1
MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.31 1.075 4.205 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.455 1.075 5.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.71 1.445 ;
        RECT 0.085 1.445 2.03 1.615 ;
        RECT 1.7 1.075 2.03 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.075 1.48 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.645 1.4 0.725 ;
        RECT 1.07 0.725 2.66 0.905 ;
        RECT 2.33 0.255 2.66 0.725 ;
        RECT 2.37 0.905 2.66 1.66 ;
        RECT 2.37 1.66 2.62 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.27 1.785 2.2 1.955 ;
      RECT 0.27 1.955 0.52 2.465 ;
      RECT 0.31 0.085 0.48 0.895 ;
      RECT 0.65 0.255 1.82 0.475 ;
      RECT 0.65 0.475 0.9 0.895 ;
      RECT 0.69 2.135 0.94 2.635 ;
      RECT 1.11 1.955 1.36 2.465 ;
      RECT 1.53 2.135 1.78 2.635 ;
      RECT 1.95 1.955 2.2 2.295 ;
      RECT 1.95 2.295 3.04 2.465 ;
      RECT 1.99 0.085 2.16 0.555 ;
      RECT 2.79 1.795 3.04 2.295 ;
      RECT 2.83 0.085 3.52 0.555 ;
      RECT 2.83 0.995 3.12 1.325 ;
      RECT 2.95 0.725 4.86 0.905 ;
      RECT 2.95 0.905 3.12 0.995 ;
      RECT 2.95 1.325 3.12 1.445 ;
      RECT 2.95 1.445 4.82 1.615 ;
      RECT 3.31 1.785 4.4 1.965 ;
      RECT 3.31 1.965 3.56 2.465 ;
      RECT 3.69 0.255 4.02 0.725 ;
      RECT 3.73 2.135 3.98 2.635 ;
      RECT 4.15 1.965 4.4 2.295 ;
      RECT 4.15 2.295 5.24 2.465 ;
      RECT 4.19 0.085 4.36 0.555 ;
      RECT 4.53 0.255 4.86 0.725 ;
      RECT 4.57 1.615 4.82 2.125 ;
      RECT 4.99 1.455 5.24 2.295 ;
      RECT 5.03 0.085 5.2 0.905 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2
MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945 1.075 7.32 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595 1.075 9.045 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 1.555 1.285 ;
        RECT 1.385 1.285 1.555 1.445 ;
        RECT 1.385 1.445 3.575 1.615 ;
        RECT 3.245 1.075 3.575 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725 1.075 3.075 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 0.645 2.995 0.725 ;
        RECT 1.775 0.725 5.045 0.905 ;
        RECT 3.745 0.905 3.915 1.415 ;
        RECT 3.745 1.415 4.965 1.615 ;
        RECT 3.875 0.275 4.205 0.725 ;
        RECT 3.915 1.615 4.165 2.125 ;
        RECT 4.715 0.275 5.045 0.725 ;
        RECT 4.745 1.615 4.965 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.085 1.455 1.215 1.625 ;
      RECT 0.085 1.625 0.425 2.465 ;
      RECT 0.175 0.085 0.345 0.895 ;
      RECT 0.515 0.255 0.845 0.725 ;
      RECT 0.515 0.725 1.605 0.905 ;
      RECT 0.595 1.795 0.805 2.635 ;
      RECT 0.975 1.625 1.215 1.795 ;
      RECT 0.975 1.795 3.745 1.965 ;
      RECT 0.975 1.965 1.215 2.465 ;
      RECT 1.015 0.085 1.185 0.555 ;
      RECT 1.355 0.255 3.365 0.475 ;
      RECT 1.355 0.475 1.605 0.725 ;
      RECT 1.395 2.135 1.645 2.635 ;
      RECT 1.815 1.965 2.065 2.465 ;
      RECT 2.235 2.135 2.485 2.635 ;
      RECT 2.655 1.965 2.905 2.465 ;
      RECT 3.075 2.135 3.325 2.635 ;
      RECT 3.495 1.965 3.745 2.295 ;
      RECT 3.495 2.295 5.465 2.465 ;
      RECT 3.535 0.085 3.705 0.555 ;
      RECT 4.085 1.075 5.725 1.245 ;
      RECT 4.335 1.795 4.575 2.295 ;
      RECT 4.375 0.085 4.545 0.555 ;
      RECT 5.135 1.455 5.465 2.295 ;
      RECT 5.215 0.085 5.905 0.555 ;
      RECT 5.555 0.735 9.575 0.905 ;
      RECT 5.555 0.905 5.725 1.075 ;
      RECT 5.655 1.455 7.625 1.625 ;
      RECT 5.655 1.625 5.985 2.465 ;
      RECT 6.075 0.255 6.405 0.725 ;
      RECT 6.075 0.725 8.925 0.735 ;
      RECT 6.155 1.795 6.365 2.635 ;
      RECT 6.54 1.625 6.78 2.465 ;
      RECT 6.575 0.085 6.745 0.555 ;
      RECT 6.915 0.255 7.245 0.725 ;
      RECT 6.955 1.795 7.205 2.635 ;
      RECT 7.375 1.625 7.625 2.295 ;
      RECT 7.375 2.295 9.31 2.465 ;
      RECT 7.415 0.085 7.585 0.555 ;
      RECT 7.755 0.255 8.085 0.725 ;
      RECT 7.795 1.455 9.575 1.625 ;
      RECT 7.795 1.625 8.045 2.125 ;
      RECT 8.215 1.795 8.465 2.295 ;
      RECT 8.255 0.085 8.425 0.555 ;
      RECT 8.595 0.255 8.925 0.725 ;
      RECT 8.635 1.625 8.885 2.125 ;
      RECT 9.06 1.795 9.31 2.295 ;
      RECT 9.095 0.085 9.265 0.555 ;
      RECT 9.215 0.905 9.575 1.455 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4
MACRO sky130_fd_sc_hd__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.78 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 2.625 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.87 1.075 4.23 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 5.26 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305 0.255 6.635 0.715 ;
        RECT 6.305 0.715 8.135 0.905 ;
        RECT 6.305 1.495 8.135 1.665 ;
        RECT 6.305 1.665 6.635 2.465 ;
        RECT 7.145 0.255 7.475 0.715 ;
        RECT 7.145 1.665 7.475 2.465 ;
        RECT 7.645 0.905 8.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 8.47 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 8.28 0.085 ;
      RECT 0 2.635 8.28 2.805 ;
      RECT 0.085 0.255 0.345 0.635 ;
      RECT 0.085 0.635 2.965 0.885 ;
      RECT 0.085 1.445 1.265 1.665 ;
      RECT 0.085 1.665 0.425 2.465 ;
      RECT 0.515 0.085 2.545 0.465 ;
      RECT 0.595 1.835 0.765 2.635 ;
      RECT 0.935 1.665 1.265 2.295 ;
      RECT 0.935 2.295 2.105 2.465 ;
      RECT 1.435 1.445 2.625 1.69 ;
      RECT 1.435 1.69 1.605 2.045 ;
      RECT 1.775 1.86 2.105 2.295 ;
      RECT 2.295 1.69 2.625 2.295 ;
      RECT 2.295 2.295 3.465 2.465 ;
      RECT 2.715 0.255 5.695 0.465 ;
      RECT 2.715 0.465 2.965 0.635 ;
      RECT 2.795 1.105 3.645 1.275 ;
      RECT 2.795 1.275 2.965 2.045 ;
      RECT 3.135 1.445 3.465 2.295 ;
      RECT 3.455 0.635 5.775 0.805 ;
      RECT 3.455 0.805 3.645 1.105 ;
      RECT 3.655 1.445 3.985 1.785 ;
      RECT 3.655 1.785 4.825 1.955 ;
      RECT 3.655 1.955 3.985 2.465 ;
      RECT 4.155 2.125 4.325 2.635 ;
      RECT 4.4 0.805 4.62 1.445 ;
      RECT 4.4 1.445 5.195 1.615 ;
      RECT 4.495 1.955 4.825 2.285 ;
      RECT 4.495 2.285 5.695 2.465 ;
      RECT 5.025 1.615 5.195 2.115 ;
      RECT 5.365 1.445 5.695 2.285 ;
      RECT 5.52 0.805 5.775 1.075 ;
      RECT 5.52 1.075 7.475 1.245 ;
      RECT 5.52 1.245 6.135 1.265 ;
      RECT 5.965 0.085 6.135 0.885 ;
      RECT 5.965 1.835 6.135 2.635 ;
      RECT 6.805 0.085 6.975 0.545 ;
      RECT 6.805 1.835 6.975 2.635 ;
      RECT 7.645 0.085 7.9 0.545 ;
      RECT 7.645 1.835 7.9 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
  END
END sky130_fd_sc_hd__o32a_4
MACRO sky130_fd_sc_hd__o32a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 0.995 1.175 1.075 ;
        RECT 1.005 1.075 1.255 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.995 1.81 1.325 ;
        RECT 1.485 1.325 1.81 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 0.995 2.255 1.66 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.995 3.595 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.795 1.66 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.595 0.825 ;
        RECT 0.085 0.825 0.26 1.495 ;
        RECT 0.085 1.495 0.47 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.14 -0.085 0.31 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.445 0.995 0.635 1.075 ;
      RECT 0.445 1.075 0.81 1.325 ;
      RECT 0.64 1.325 0.81 1.495 ;
      RECT 0.64 1.495 1.315 1.665 ;
      RECT 0.685 1.835 0.975 2.635 ;
      RECT 0.765 0.085 0.935 0.645 ;
      RECT 1.14 0.255 1.47 0.655 ;
      RECT 1.14 0.655 2.54 0.825 ;
      RECT 1.145 1.665 1.315 2.295 ;
      RECT 1.145 2.295 2.51 2.465 ;
      RECT 1.645 0.085 1.975 0.485 ;
      RECT 2.18 1.835 3.135 2.085 ;
      RECT 2.18 2.085 2.51 2.295 ;
      RECT 2.21 0.255 3.595 0.465 ;
      RECT 2.21 0.465 2.54 0.655 ;
      RECT 2.71 0.635 3.135 0.825 ;
      RECT 2.965 0.825 3.135 1.835 ;
      RECT 3.305 0.465 3.595 0.735 ;
      RECT 3.305 1.495 3.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__o32a_1
MACRO sky130_fd_sc_hd__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.715 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.16 1.615 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.995 2.635 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695 1.075 4.055 1.245 ;
        RECT 3.725 1.245 4.055 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.91 0.995 3.155 1.615 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.085 0.085 0.345 0.885 ;
      RECT 0.085 1.495 0.345 2.635 ;
      RECT 1.015 0.995 1.325 1.785 ;
      RECT 1.015 1.785 3.525 1.955 ;
      RECT 1.015 2.125 1.525 2.635 ;
      RECT 1.095 0.085 1.425 0.825 ;
      RECT 1.695 0.255 2.025 0.655 ;
      RECT 1.695 0.655 3.025 0.825 ;
      RECT 2.195 0.085 2.525 0.485 ;
      RECT 2.695 0.255 4.055 0.425 ;
      RECT 2.695 0.425 3.025 0.655 ;
      RECT 2.695 1.955 3.025 2.465 ;
      RECT 3.195 0.595 3.525 0.825 ;
      RECT 3.325 0.825 3.525 1.785 ;
      RECT 3.695 0.425 4.055 0.905 ;
      RECT 3.695 1.495 4.055 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__o32a_2
MACRO sky130_fd_sc_hd__sedfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.48 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755 0.305 13.085 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.8 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.885 1.435 ;
        RECT -0.19 1.435 13.99 2.91 ;
        RECT 7.2 1.305 13.99 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.8 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 13.8 0.085 ;
      RECT 0 2.635 13.8 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 5.665 2.175 6.01 2.635 ;
      RECT 5.76 0.085 6.01 0.905 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.245 0.085 8.64 0.56 ;
      RECT 8.425 1.835 8.66 2.635 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 9.37 2.105 9.66 2.635 ;
      RECT 9.465 0.085 9.74 0.615 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.28 2.135 11.54 2.635 ;
      RECT 11.35 0.085 11.665 0.615 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
      RECT 12.35 0.085 12.585 0.9 ;
      RECT 12.35 1.465 12.585 2.635 ;
      RECT 13.255 0.085 13.515 0.9 ;
      RECT 13.255 1.465 13.515 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12 0.765 12.17 0.935 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_2
MACRO sky130_fd_sc_hd__sedfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.4 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755 0.305 13.085 1.07 ;
        RECT 12.755 1.07 13.925 1.295 ;
        RECT 12.755 1.295 13.085 2.42 ;
        RECT 13.595 0.305 13.925 1.07 ;
        RECT 13.595 1.295 13.925 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.72 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.885 1.435 ;
        RECT -0.19 1.435 14.91 2.91 ;
        RECT 7.2 1.305 14.91 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.72 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 14.72 0.085 ;
      RECT 0 2.635 14.72 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 5.665 2.175 6.01 2.635 ;
      RECT 5.76 0.085 6.01 0.905 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.245 0.085 8.64 0.56 ;
      RECT 8.425 1.835 8.66 2.635 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 9.37 2.105 9.66 2.635 ;
      RECT 9.465 0.085 9.74 0.615 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.28 2.135 11.54 2.635 ;
      RECT 11.35 0.085 11.665 0.615 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
      RECT 12.35 0.085 12.585 0.9 ;
      RECT 12.35 1.465 12.585 2.635 ;
      RECT 13.255 0.085 13.425 0.9 ;
      RECT 13.255 1.465 13.425 2.635 ;
      RECT 14.095 0.085 14.355 1.28 ;
      RECT 14.095 1.465 14.355 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12 0.765 12.17 0.935 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.485 2.635 13.655 2.805 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.945 2.635 14.115 2.805 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 14.405 2.635 14.575 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_4
MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765 0.305 13.095 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.885 1.435 ;
        RECT -0.19 1.435 13.53 2.91 ;
        RECT 7.2 1.305 13.53 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 13.34 0.085 ;
      RECT 0 2.635 13.34 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.235 0.085 2.565 0.515 ;
      RECT 2.235 1.89 2.565 2.635 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.185 0.085 3.515 0.61 ;
      RECT 3.265 1.825 3.46 2.635 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 5.665 2.175 6.01 2.635 ;
      RECT 5.76 0.085 6.01 0.905 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.245 0.085 8.64 0.56 ;
      RECT 8.425 1.835 8.66 2.635 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 9.37 2.105 9.66 2.635 ;
      RECT 9.465 0.085 9.74 0.615 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.28 2.135 11.54 2.635 ;
      RECT 11.35 0.085 11.665 0.615 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
      RECT 12.35 0.085 12.595 0.9 ;
      RECT 12.35 1.465 12.595 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 12 0.765 12.17 0.935 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 12.105 2.635 12.275 2.805 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.565 2.635 12.735 2.805 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 13.025 2.635 13.195 2.805 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_1
MACRO sky130_fd_sc_hd__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.47 1.315 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.255 1.185 0.735 ;
        RECT 1.015 0.735 2.025 0.905 ;
        RECT 1.015 1.445 2.025 1.615 ;
        RECT 1.015 1.615 1.185 2.465 ;
        RECT 1.53 0.905 2.025 1.445 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 1.615 2.025 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.095 1.485 0.81 1.655 ;
      RECT 0.095 1.655 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 0.81 0.905 ;
      RECT 0.525 0.085 0.765 0.565 ;
      RECT 0.595 1.835 0.835 2.635 ;
      RECT 0.64 0.905 0.81 1.075 ;
      RECT 0.64 1.075 1.14 1.245 ;
      RECT 0.64 1.245 0.81 1.485 ;
      RECT 1.355 0.085 1.685 0.565 ;
      RECT 1.355 1.835 1.685 2.635 ;
      RECT 2.195 0.085 2.525 0.885 ;
      RECT 2.195 1.485 2.525 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__buf_4
MACRO sky130_fd_sc_hd__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.28 1.075 1.185 1.315 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.255 1.865 0.735 ;
        RECT 1.695 0.735 3.545 0.905 ;
        RECT 1.695 1.445 3.545 1.615 ;
        RECT 1.695 1.615 1.865 2.465 ;
        RECT 2.21 0.905 3.545 1.445 ;
        RECT 2.535 0.255 2.705 0.735 ;
        RECT 2.535 1.615 2.705 2.465 ;
        RECT 3.375 0.255 3.545 0.735 ;
        RECT 3.375 1.615 3.545 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.33 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.14 0.085 ;
      RECT 0 2.635 4.14 2.805 ;
      RECT 0.435 0.085 0.605 0.565 ;
      RECT 0.435 1.485 0.605 2.635 ;
      RECT 0.775 0.255 1.105 0.735 ;
      RECT 0.775 0.735 1.525 0.905 ;
      RECT 0.775 1.485 1.525 1.655 ;
      RECT 0.775 1.655 1.105 2.465 ;
      RECT 1.275 0.085 1.445 0.565 ;
      RECT 1.275 1.835 1.515 2.635 ;
      RECT 1.355 0.905 1.525 1.075 ;
      RECT 1.355 1.075 1.825 1.245 ;
      RECT 1.355 1.245 1.525 1.485 ;
      RECT 2.035 0.085 2.365 0.565 ;
      RECT 2.035 1.835 2.365 2.635 ;
      RECT 2.875 0.085 3.205 0.565 ;
      RECT 2.875 1.835 3.205 2.635 ;
      RECT 3.715 0.085 4.045 0.885 ;
      RECT 3.715 1.485 4.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
  END
END sky130_fd_sc_hd__buf_6
MACRO sky130_fd_sc_hd__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 4.29 0.905 4.545 1.445 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.375 1.615 4.545 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.515 0.085 0.845 0.565 ;
      RECT 0.595 1.835 0.765 2.635 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.355 0.085 1.685 0.565 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
      RECT 1.435 1.835 1.605 2.635 ;
      RECT 2.195 0.085 2.525 0.565 ;
      RECT 2.195 1.835 2.525 2.635 ;
      RECT 3.035 0.085 3.365 0.565 ;
      RECT 3.035 1.835 3.365 2.635 ;
      RECT 3.875 0.085 4.205 0.565 ;
      RECT 3.875 1.835 4.205 2.635 ;
      RECT 4.715 0.085 5.045 0.885 ;
      RECT 4.715 1.485 5.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__buf_8
MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.44 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 0.255 1.315 0.83 ;
        RECT 1.06 1.56 1.315 2.465 ;
        RECT 1.145 0.83 1.315 1.56 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.03 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.84 0.085 ;
      RECT 0 2.635 1.84 2.805 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.89 0.805 ;
      RECT 0.175 1.535 0.89 1.705 ;
      RECT 0.175 1.705 0.345 2.465 ;
      RECT 0.56 0.085 0.89 0.465 ;
      RECT 0.56 1.875 0.89 2.635 ;
      RECT 0.72 0.805 0.89 0.995 ;
      RECT 0.72 0.995 0.975 1.325 ;
      RECT 0.72 1.325 0.89 1.535 ;
      RECT 1.49 0.085 1.75 0.925 ;
      RECT 1.49 1.485 1.75 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
  END
END sky130_fd_sc_hd__buf_2
MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.985 0.445 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.56 1.295 2.465 ;
        RECT 1.035 0.255 1.295 0.76 ;
        RECT 1.115 0.76 1.295 1.56 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.085 0.325 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.57 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.38 0.085 ;
      RECT 0 2.635 1.38 2.805 ;
      RECT 0.165 1.535 0.84 1.705 ;
      RECT 0.165 1.705 0.345 2.465 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.525 0.085 0.855 0.465 ;
      RECT 0.525 1.875 0.855 2.635 ;
      RECT 0.67 0.805 0.84 1.06 ;
      RECT 0.67 1.06 0.945 1.39 ;
      RECT 0.67 1.39 0.84 1.535 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
  END
END sky130_fd_sc_hd__buf_1
MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 2.485 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035 0.255 3.285 0.26 ;
        RECT 3.035 0.26 3.365 0.735 ;
        RECT 3.035 0.735 10.035 0.905 ;
        RECT 3.035 1.445 10.035 1.615 ;
        RECT 3.035 1.615 3.365 2.465 ;
        RECT 3.875 0.26 4.205 0.735 ;
        RECT 3.875 1.615 4.205 2.465 ;
        RECT 3.955 0.255 4.125 0.26 ;
        RECT 4.715 0.26 5.045 0.735 ;
        RECT 4.715 1.615 5.045 2.465 ;
        RECT 4.795 0.255 4.965 0.26 ;
        RECT 5.555 0.26 5.885 0.735 ;
        RECT 5.555 1.615 5.885 2.465 ;
        RECT 6.395 0.26 6.725 0.735 ;
        RECT 6.395 1.615 6.725 2.465 ;
        RECT 7.235 0.26 7.565 0.735 ;
        RECT 7.235 1.615 7.565 2.465 ;
        RECT 8.075 0.26 8.405 0.735 ;
        RECT 8.075 1.615 8.405 2.465 ;
        RECT 8.915 0.26 9.245 0.735 ;
        RECT 8.915 1.615 9.245 2.465 ;
        RECT 9.655 0.905 10.035 1.445 ;
        RECT 9.76 0.365 10.035 0.735 ;
        RECT 9.76 1.615 10.035 2.36 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.175 0.085 0.345 0.905 ;
      RECT 0.175 1.445 0.345 2.635 ;
      RECT 0.515 0.26 0.845 0.735 ;
      RECT 0.515 0.735 2.865 0.905 ;
      RECT 0.515 1.445 2.865 1.615 ;
      RECT 0.515 1.615 0.845 2.465 ;
      RECT 1.015 0.085 1.185 0.565 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.355 0.26 1.685 0.735 ;
      RECT 1.355 1.615 1.685 2.465 ;
      RECT 1.855 0.085 2.025 0.565 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.195 0.26 2.525 0.735 ;
      RECT 2.195 1.615 2.525 2.465 ;
      RECT 2.69 0.905 2.865 1.075 ;
      RECT 2.69 1.075 9.41 1.275 ;
      RECT 2.69 1.275 2.865 1.445 ;
      RECT 2.695 0.085 2.865 0.565 ;
      RECT 2.695 1.835 2.865 2.635 ;
      RECT 3.535 0.085 3.705 0.565 ;
      RECT 3.535 1.835 3.705 2.635 ;
      RECT 4.375 0.085 4.545 0.565 ;
      RECT 4.375 1.835 4.545 2.635 ;
      RECT 5.215 0.085 5.385 0.565 ;
      RECT 5.215 1.835 5.385 2.635 ;
      RECT 6.055 0.085 6.225 0.565 ;
      RECT 6.055 1.835 6.225 2.635 ;
      RECT 6.895 0.085 7.065 0.565 ;
      RECT 6.895 1.835 7.065 2.635 ;
      RECT 7.735 0.085 7.905 0.565 ;
      RECT 7.735 1.835 7.905 2.635 ;
      RECT 8.575 0.085 8.745 0.565 ;
      RECT 8.575 1.835 8.745 2.635 ;
      RECT 9.415 0.085 9.585 0.565 ;
      RECT 9.415 1.835 9.585 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__buf_16
MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 1.66 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.255 2.445 0.735 ;
        RECT 2.275 0.735 6.645 0.905 ;
        RECT 2.275 1.445 6.645 1.615 ;
        RECT 2.275 1.615 2.445 2.465 ;
        RECT 3.115 0.255 3.285 0.735 ;
        RECT 3.115 1.615 3.285 2.465 ;
        RECT 3.955 0.255 4.125 0.735 ;
        RECT 3.955 1.615 4.125 2.465 ;
        RECT 4.71 0.905 6.645 1.445 ;
        RECT 4.795 0.255 4.965 0.735 ;
        RECT 4.795 1.615 4.965 2.465 ;
        RECT 5.635 0.255 5.805 0.735 ;
        RECT 5.635 1.615 5.805 2.465 ;
        RECT 6.475 0.255 6.645 0.735 ;
        RECT 6.475 1.615 6.645 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.57 -0.085 0.74 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 0.095 0.085 0.425 0.565 ;
      RECT 0.175 1.835 0.345 2.635 ;
      RECT 0.515 1.445 2.015 1.615 ;
      RECT 0.515 1.615 0.845 2.465 ;
      RECT 0.595 0.255 0.765 0.735 ;
      RECT 0.595 0.735 2.015 0.905 ;
      RECT 0.935 0.085 1.265 0.565 ;
      RECT 1.015 1.835 1.185 2.635 ;
      RECT 1.355 1.615 1.685 2.465 ;
      RECT 1.435 0.26 1.605 0.735 ;
      RECT 1.775 0.085 2.105 0.565 ;
      RECT 1.84 0.905 2.015 1.075 ;
      RECT 1.84 1.075 4.465 1.245 ;
      RECT 1.84 1.245 2.015 1.445 ;
      RECT 1.855 1.835 2.025 2.635 ;
      RECT 2.615 0.085 2.945 0.565 ;
      RECT 2.615 1.835 2.945 2.635 ;
      RECT 3.455 0.085 3.785 0.565 ;
      RECT 3.455 1.835 3.785 2.635 ;
      RECT 4.295 0.085 4.625 0.565 ;
      RECT 4.295 1.835 4.625 2.635 ;
      RECT 5.135 0.085 5.465 0.565 ;
      RECT 5.135 1.835 5.465 2.635 ;
      RECT 5.975 0.085 6.305 0.565 ;
      RECT 5.975 1.835 6.305 2.635 ;
      RECT 6.815 0.085 7.145 0.885 ;
      RECT 6.815 1.485 7.145 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
  END
END sky130_fd_sc_hd__buf_12
MACRO sky130_fd_sc_hd__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 0.415 6.355 2.455 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.5 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 1.025 ;
      RECT 3.33 1.025 4.33 1.245 ;
      RECT 3.48 1.245 4.33 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.74 0.085 4.07 0.53 ;
      RECT 3.82 1.535 5.925 1.865 ;
      RECT 3.82 2.135 4.11 2.635 ;
      RECT 4.24 0.255 4.59 0.655 ;
      RECT 4.24 0.655 5.925 0.825 ;
      RECT 4.3 2.135 4.58 2.635 ;
      RECT 4.75 1.865 4.94 2.465 ;
      RECT 5.095 0.085 5.925 0.485 ;
      RECT 5.11 2.135 5.925 2.635 ;
      RECT 5.605 0.825 5.925 1.535 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_1
MACRO sky130_fd_sc_hd__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.255 5.965 0.485 ;
        RECT 5.68 1.875 5.965 2.465 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 0.255 6.775 0.765 ;
        RECT 6.575 1.325 6.775 2.465 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.55 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.96 1.835 2.275 2.635 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.46 1.495 2.145 1.665 ;
      RECT 1.46 1.665 1.79 2.415 ;
      RECT 1.54 0.345 1.71 0.615 ;
      RECT 1.54 0.615 2.145 0.765 ;
      RECT 1.54 0.765 2.345 0.785 ;
      RECT 1.88 0.085 2.21 0.445 ;
      RECT 1.975 0.785 2.345 1.095 ;
      RECT 1.975 1.095 2.145 1.495 ;
      RECT 2.475 1.355 2.76 2.005 ;
      RECT 2.72 0.705 3.1 1.035 ;
      RECT 2.845 0.365 3.505 0.535 ;
      RECT 2.905 2.255 3.655 2.425 ;
      RECT 2.93 1.035 3.1 1.415 ;
      RECT 2.93 1.415 3.27 1.995 ;
      RECT 3.335 0.535 3.505 1.025 ;
      RECT 3.335 1.025 4.315 1.245 ;
      RECT 3.485 1.245 4.315 1.325 ;
      RECT 3.485 1.325 3.655 2.255 ;
      RECT 3.745 0.085 4.075 0.53 ;
      RECT 3.825 1.535 5.625 1.705 ;
      RECT 3.825 1.705 4.945 1.865 ;
      RECT 4.245 0.255 4.595 0.655 ;
      RECT 4.245 0.655 5.625 0.825 ;
      RECT 4.755 1.865 4.945 2.465 ;
      RECT 5.1 0.085 5.44 0.485 ;
      RECT 5.455 0.825 5.625 1.535 ;
      RECT 6.135 0.085 6.405 0.595 ;
      RECT 6.945 0.085 7.275 0.595 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.475 1.785 2.645 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.935 1.445 3.105 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.165 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.705 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.415 1.755 2.705 1.8 ;
      RECT 2.415 1.94 2.705 1.985 ;
      RECT 2.875 1.415 3.165 1.46 ;
      RECT 2.875 1.6 3.165 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_4
MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595 0.255 5.925 0.485 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 1.425 6.355 1.5 ;
        RECT 5.755 1.5 5.925 1.875 ;
        RECT 5.76 1.415 6.355 1.425 ;
        RECT 5.765 1.41 6.355 1.415 ;
        RECT 5.77 0.865 6.355 0.89 ;
        RECT 5.775 1.385 6.355 1.41 ;
        RECT 5.785 0.89 6.355 1.385 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.48 0.995 5.17 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 6.63 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.44 0.085 ;
      RECT 0 2.635 6.44 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.875 0.085 2.205 0.445 ;
      RECT 1.955 1.835 2.27 2.635 ;
      RECT 1.96 0.785 2.34 1.095 ;
      RECT 1.96 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.675 0.705 3.095 1.145 ;
      RECT 2.775 2.255 3.605 2.425 ;
      RECT 2.81 0.365 3.5 0.535 ;
      RECT 2.925 1.145 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 1.025 ;
      RECT 3.33 1.025 4.31 1.245 ;
      RECT 3.435 1.245 4.31 1.325 ;
      RECT 3.435 1.325 3.605 2.255 ;
      RECT 3.735 0.085 4.07 0.53 ;
      RECT 3.8 2.135 4.11 2.635 ;
      RECT 3.82 1.535 5.585 1.705 ;
      RECT 3.82 1.705 4.92 1.865 ;
      RECT 4.24 0.255 4.59 0.655 ;
      RECT 4.24 0.655 5.585 0.825 ;
      RECT 4.28 2.135 4.56 2.635 ;
      RECT 4.73 1.865 4.92 2.465 ;
      RECT 5.09 1.875 5.46 2.635 ;
      RECT 5.095 0.085 5.425 0.485 ;
      RECT 5.35 0.995 5.615 1.325 ;
      RECT 5.415 0.825 5.585 0.995 ;
      RECT 5.415 1.325 5.585 1.535 ;
      RECT 6.095 0.085 6.355 0.595 ;
      RECT 6.095 1.67 6.355 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_2
MACRO sky130_fd_sc_hd__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.18 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
      LAYER mcon ;
        RECT 6.865 0.765 7.035 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
      LAYER mcon ;
        RECT 9.69 1.105 9.86 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.5 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215 -0.01 0.235 0.015 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 1.97 1.425 ;
        RECT -0.19 1.425 11.69 2.91 ;
        RECT 4.405 1.305 11.69 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.5 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.5 0.085 ;
      RECT 0 2.635 11.5 2.805 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.53 2.135 0.86 2.635 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.875 0.085 2.205 0.56 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.32 2.04 2.49 2.635 ;
      RECT 2.395 0.085 2.725 0.825 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.3 2.275 4.63 2.635 ;
      RECT 4.445 0.085 4.775 0.54 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.41 2.355 6.74 2.635 ;
      RECT 6.915 0.085 7.245 0.545 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.375 2.175 7.745 2.635 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.085 0.085 9.255 0.525 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.36 2.195 9.61 2.635 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.12 2.255 10.45 2.635 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.72 0.085 10.89 0.545 ;
      RECT 10.72 1.495 10.97 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.675 1.785 0.845 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.145 1.105 1.315 1.275 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.445 1.785 8.615 1.955 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
    LAYER met1 ;
      RECT 0.615 1.755 0.915 1.8 ;
      RECT 0.615 1.8 8.675 1.94 ;
      RECT 0.615 1.94 0.915 1.985 ;
      RECT 1.085 1.075 1.375 1.12 ;
      RECT 1.085 1.12 8.635 1.26 ;
      RECT 1.085 1.26 1.375 1.305 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtn_1
MACRO sky130_fd_sc_hd__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.43 1.075 3.76 1.445 ;
        RECT 3.43 1.445 4.815 1.615 ;
        RECT 4.645 1.075 5.435 1.275 ;
        RECT 4.645 1.275 4.815 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.98 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.02 1.075 2.035 1.445 ;
        RECT 1.02 1.445 3.26 1.615 ;
        RECT 2.93 1.075 3.26 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 2.76 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.52 0.645 0.85 0.865 ;
        RECT 0.56 1.445 0.85 1.785 ;
        RECT 0.56 1.785 4.35 1.955 ;
        RECT 0.56 1.955 0.81 2.465 ;
        RECT 0.605 0.865 0.85 1.445 ;
        RECT 2.34 1.955 2.59 2.125 ;
        RECT 4.1 1.955 4.35 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.1 0.255 1.27 0.475 ;
      RECT 0.1 0.475 0.35 0.895 ;
      RECT 0.14 1.455 0.39 2.635 ;
      RECT 0.98 2.125 1.75 2.635 ;
      RECT 1.02 0.475 1.27 0.645 ;
      RECT 1.02 0.645 3.05 0.905 ;
      RECT 1.46 0.255 3.55 0.475 ;
      RECT 1.92 2.125 2.17 2.295 ;
      RECT 1.92 2.295 3.01 2.465 ;
      RECT 2.76 2.125 3.01 2.295 ;
      RECT 3.18 2.125 3.51 2.635 ;
      RECT 3.22 0.475 3.55 0.735 ;
      RECT 3.22 0.735 5.23 0.905 ;
      RECT 3.68 2.125 3.93 2.295 ;
      RECT 3.68 2.295 4.77 2.465 ;
      RECT 3.72 0.085 3.89 0.555 ;
      RECT 4.06 0.255 4.39 0.725 ;
      RECT 4.06 0.725 5.23 0.735 ;
      RECT 4.52 1.785 4.77 2.295 ;
      RECT 4.56 0.085 4.73 0.555 ;
      RECT 4.9 0.255 5.23 0.725 ;
      RECT 4.985 1.455 5.19 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__o221ai_2
MACRO sky130_fd_sc_hd__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165 1.075 2.505 1.245 ;
        RECT 2.295 1.245 2.505 1.445 ;
        RECT 2.295 1.445 2.675 1.615 ;
        RECT 2.465 1.615 2.675 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.995 1.355 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.985 1.325 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.465 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.899000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.345 0.645 ;
        RECT 0.085 0.645 0.84 0.825 ;
        RECT 0.085 1.495 2.125 1.705 ;
        RECT 0.085 1.705 0.365 2.465 ;
        RECT 0.635 0.825 0.84 1.495 ;
        RECT 1.735 1.705 2.125 1.785 ;
        RECT 1.735 1.785 2.245 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.515 0.305 1.775 0.475 ;
      RECT 0.55 1.875 1.34 2.635 ;
      RECT 1.01 0.645 2.22 0.695 ;
      RECT 1.01 0.695 3.135 0.825 ;
      RECT 1.945 0.28 2.22 0.645 ;
      RECT 2.105 0.825 3.135 0.865 ;
      RECT 2.455 0.085 2.625 0.525 ;
      RECT 2.795 0.28 3.135 0.695 ;
      RECT 2.875 1.455 3.135 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__o221ai_1
MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 5.965 1.445 8.42 1.615 ;
        RECT 8.155 1.075 9.575 1.275 ;
        RECT 8.155 1.275 8.42 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.36 1.075 4.505 1.275 ;
        RECT 4.335 1.275 4.505 1.495 ;
        RECT 4.335 1.495 5.795 1.665 ;
        RECT 5.465 1.075 5.795 1.495 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675 0.995 5.285 1.325 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.75 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.645 2.125 0.865 ;
        RECT 0.575 1.445 4.165 1.615 ;
        RECT 0.575 1.615 0.825 2.465 ;
        RECT 1.415 1.615 2.125 1.955 ;
        RECT 1.415 1.955 1.665 2.465 ;
        RECT 1.92 0.865 2.125 1.445 ;
        RECT 3.995 1.615 4.165 1.835 ;
        RECT 3.995 1.835 7.725 1.955 ;
        RECT 3.995 1.955 6.885 2.005 ;
        RECT 3.995 2.005 4.285 2.125 ;
        RECT 4.875 2.005 5.085 2.125 ;
        RECT 5.965 1.785 7.725 1.835 ;
        RECT 6.675 2.005 6.885 2.125 ;
        RECT 7.475 1.955 7.725 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.115 0.255 5.585 0.475 ;
      RECT 0.115 0.475 0.365 0.895 ;
      RECT 0.155 1.485 0.405 2.635 ;
      RECT 0.995 1.825 1.245 2.635 ;
      RECT 1.835 2.125 2.605 2.635 ;
      RECT 2.315 0.645 6.085 0.735 ;
      RECT 2.315 0.735 9.445 0.82 ;
      RECT 2.775 1.785 3.825 1.955 ;
      RECT 2.775 1.955 3.025 2.465 ;
      RECT 3.195 2.125 3.445 2.635 ;
      RECT 3.615 1.955 3.825 2.295 ;
      RECT 3.615 2.295 5.585 2.465 ;
      RECT 4.455 2.175 4.705 2.295 ;
      RECT 5.255 2.175 5.585 2.295 ;
      RECT 5.465 0.82 9.445 0.905 ;
      RECT 5.755 0.255 6.085 0.645 ;
      RECT 5.755 2.175 6.005 2.635 ;
      RECT 6.175 2.175 6.505 2.295 ;
      RECT 6.175 2.295 8.145 2.465 ;
      RECT 6.255 0.085 6.425 0.555 ;
      RECT 6.595 0.255 6.925 0.725 ;
      RECT 6.595 0.725 7.765 0.735 ;
      RECT 7.055 2.125 7.305 2.295 ;
      RECT 7.095 0.085 7.265 0.555 ;
      RECT 7.435 0.255 7.765 0.725 ;
      RECT 7.895 1.785 8.985 1.955 ;
      RECT 7.895 1.955 8.145 2.295 ;
      RECT 7.935 0.085 8.105 0.555 ;
      RECT 8.275 0.255 8.605 0.725 ;
      RECT 8.275 0.725 9.445 0.735 ;
      RECT 8.315 2.125 8.565 2.635 ;
      RECT 8.735 1.445 8.985 1.785 ;
      RECT 8.735 1.955 8.985 2.465 ;
      RECT 8.775 0.085 8.945 0.555 ;
      RECT 9.115 0.255 9.445 0.725 ;
      RECT 9.155 1.445 9.405 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
  END
END sky130_fd_sc_hd__o221ai_4
MACRO sky130_fd_sc_hd__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.675 0.255 9.005 0.735 ;
        RECT 8.675 0.735 10.44 0.905 ;
        RECT 8.715 1.455 10.44 1.625 ;
        RECT 8.715 1.625 9.005 2.465 ;
        RECT 9.515 0.255 9.845 0.735 ;
        RECT 9.555 1.625 9.805 2.465 ;
        RECT 10.03 0.905 10.44 1.455 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.77 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.58 0.085 ;
      RECT 0 2.635 10.58 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.04 2.635 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 1.075 ;
      RECT 7.815 1.075 9.845 1.285 ;
      RECT 7.815 1.285 8.16 1.295 ;
      RECT 7.99 1.295 8.16 1.915 ;
      RECT 8.335 0.085 8.505 0.895 ;
      RECT 8.335 1.575 8.505 2.635 ;
      RECT 9.175 0.085 9.345 0.555 ;
      RECT 9.175 1.795 9.345 2.635 ;
      RECT 10.015 0.085 10.185 0.555 ;
      RECT 10.015 1.795 10.185 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_4
MACRO sky130_fd_sc_hd__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.105 0.795 ;
        RECT 8.855 1.445 9.105 2.325 ;
        RECT 8.9 0.795 9.105 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.04 2.635 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.38 0.085 8.685 0.545 ;
      RECT 8.38 1.495 8.685 2.635 ;
      RECT 9.275 0.085 9.525 0.84 ;
      RECT 9.275 1.495 9.525 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_2
MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.11 0.795 ;
        RECT 8.855 1.445 9.11 2.325 ;
        RECT 8.9 0.795 9.11 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
      LAYER mcon ;
        RECT 4.165 0.765 4.335 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
      LAYER mcon ;
        RECT 7.105 1.08 7.275 1.25 ;
        RECT 7.405 0.765 7.575 0.935 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.39 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.2 0.085 ;
      RECT 0 2.635 9.2 2.805 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.545 0.085 1.875 0.445 ;
      RECT 1.85 2.175 2.1 2.635 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 3.99 2.205 4.32 2.635 ;
      RECT 4.475 0.085 4.805 0.545 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 4.955 2.175 5.325 2.635 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.085 6.895 0.525 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 6.94 2.175 7.19 2.635 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.71 2.255 8.04 2.635 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.38 0.085 8.685 0.545 ;
      RECT 8.38 1.495 8.685 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_1
MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.79 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.23 0.305 9.575 0.82 ;
        RECT 9.23 1.505 9.575 2.395 ;
        RECT 9.405 0.82 9.575 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.53 1.055 3.99 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.635 3.25 0.785 ;
        RECT 1.76 0.785 1.99 0.835 ;
        RECT 1.76 0.835 1.93 1.685 ;
        RECT 1.87 0.615 3.25 0.635 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.065 0.785 3.25 1.095 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 9.85 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.52 2.135 0.85 2.635 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.23 0.715 ;
      RECT 1.02 0.715 1.23 2.465 ;
      RECT 1.42 0.26 1.79 0.465 ;
      RECT 1.42 0.465 1.59 1.86 ;
      RECT 1.42 1.86 3.22 2.075 ;
      RECT 1.42 2.075 1.71 2.445 ;
      RECT 1.88 2.245 2.21 2.635 ;
      RECT 1.96 0.085 2.305 0.445 ;
      RECT 2.115 0.96 2.46 1.13 ;
      RECT 2.115 1.13 2.29 1.86 ;
      RECT 2.69 2.245 3.56 2.415 ;
      RECT 2.82 0.275 3.59 0.445 ;
      RECT 3.05 1.305 3.27 1.635 ;
      RECT 3.05 1.635 3.22 1.86 ;
      RECT 3.39 1.825 4.35 1.995 ;
      RECT 3.39 1.995 3.56 2.245 ;
      RECT 3.42 0.445 3.59 0.715 ;
      RECT 3.42 0.715 4.35 0.885 ;
      RECT 3.73 2.165 3.925 2.635 ;
      RECT 3.76 0.085 3.96 0.545 ;
      RECT 4.18 0.285 4.46 0.615 ;
      RECT 4.18 0.615 4.35 0.715 ;
      RECT 4.18 0.885 4.35 1.825 ;
      RECT 4.18 1.995 4.35 2.065 ;
      RECT 4.18 2.065 4.42 2.44 ;
      RECT 4.52 0.78 5.1 1.035 ;
      RECT 4.52 1.035 4.76 1.905 ;
      RECT 4.63 0.705 5.1 0.78 ;
      RECT 4.66 2.19 5.73 2.36 ;
      RECT 4.7 0.365 5.44 0.535 ;
      RECT 4.95 1.655 5.39 2.01 ;
      RECT 5.27 0.535 5.44 1.315 ;
      RECT 5.27 1.315 6.07 1.485 ;
      RECT 5.56 1.485 6.07 1.575 ;
      RECT 5.56 1.575 5.73 2.19 ;
      RECT 5.61 0.765 6.41 1.065 ;
      RECT 5.61 1.065 5.78 1.095 ;
      RECT 5.69 0.085 6.06 0.585 ;
      RECT 5.9 1.245 6.07 1.315 ;
      RECT 5.9 1.835 6.07 2.635 ;
      RECT 6.24 0.365 6.7 0.535 ;
      RECT 6.24 0.535 6.41 0.765 ;
      RECT 6.24 1.065 6.41 2.135 ;
      RECT 6.24 2.135 6.49 2.465 ;
      RECT 6.58 0.705 7.13 1.035 ;
      RECT 6.58 1.245 6.77 1.965 ;
      RECT 6.715 2.165 7.6 2.335 ;
      RECT 6.93 0.365 7.47 0.535 ;
      RECT 6.94 1.035 7.13 1.575 ;
      RECT 6.94 1.575 7.26 1.905 ;
      RECT 7.3 0.535 7.47 0.995 ;
      RECT 7.3 0.995 8.365 1.325 ;
      RECT 7.3 1.325 7.6 1.405 ;
      RECT 7.43 1.405 7.6 2.165 ;
      RECT 7.715 0.085 8.085 0.615 ;
      RECT 7.77 1.575 8.705 1.905 ;
      RECT 7.79 2.135 8.095 2.635 ;
      RECT 8.355 0.3 8.705 0.825 ;
      RECT 8.435 1.905 8.705 2.455 ;
      RECT 8.535 0.825 8.705 0.995 ;
      RECT 8.535 0.995 9.235 1.325 ;
      RECT 8.535 1.325 8.705 1.575 ;
      RECT 8.875 0.085 9.045 0.695 ;
      RECT 8.875 1.625 9.045 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.64 1.785 0.81 1.955 ;
      RECT 1.04 0.765 1.21 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.59 1.785 6.76 1.955 ;
      RECT 6.63 0.765 6.8 0.935 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
    LAYER met1 ;
      RECT 0.58 1.755 0.87 1.8 ;
      RECT 0.58 1.8 6.82 1.94 ;
      RECT 0.58 1.94 0.87 1.985 ;
      RECT 0.98 0.735 1.27 0.78 ;
      RECT 0.98 0.78 6.86 0.92 ;
      RECT 0.98 0.92 1.27 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.53 1.755 6.82 1.8 ;
      RECT 6.53 1.94 6.82 1.985 ;
      RECT 6.57 0.735 6.86 0.78 ;
      RECT 6.57 0.92 6.86 0.965 ;
  END
END sky130_fd_sc_hd__sdfxtp_1
MACRO sky130_fd_sc_hd__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.79 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.26 0.305 9.605 0.82 ;
        RECT 9.26 1.505 9.605 2.395 ;
        RECT 9.435 0.82 9.605 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.53 1.035 4.02 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.25 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.08 0.785 3.25 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.52 2.135 0.85 2.635 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.245 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 1.88 2.245 2.21 2.635 ;
      RECT 1.975 0.085 2.305 0.445 ;
      RECT 2.12 0.955 2.46 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.69 2.245 3.585 2.415 ;
      RECT 2.82 0.275 3.59 0.445 ;
      RECT 3.075 1.355 3.27 1.685 ;
      RECT 3.075 1.685 3.245 1.86 ;
      RECT 3.415 1.825 4.38 1.995 ;
      RECT 3.415 1.995 3.585 2.245 ;
      RECT 3.42 0.445 3.59 0.695 ;
      RECT 3.42 0.695 4.38 0.865 ;
      RECT 3.755 2.165 3.925 2.635 ;
      RECT 3.76 0.085 3.96 0.525 ;
      RECT 4.21 0.365 4.56 0.535 ;
      RECT 4.21 0.535 4.38 0.695 ;
      RECT 4.21 0.865 4.38 1.825 ;
      RECT 4.21 1.995 4.38 2.065 ;
      RECT 4.21 2.065 4.445 2.44 ;
      RECT 4.55 0.705 5.13 1.035 ;
      RECT 4.55 1.035 4.79 1.905 ;
      RECT 4.69 2.19 5.76 2.36 ;
      RECT 4.73 0.365 5.47 0.535 ;
      RECT 4.98 1.655 5.42 2.01 ;
      RECT 5.3 0.535 5.47 1.315 ;
      RECT 5.3 1.315 6.1 1.485 ;
      RECT 5.59 1.485 6.1 1.575 ;
      RECT 5.59 1.575 5.76 2.19 ;
      RECT 5.64 0.765 6.44 1.065 ;
      RECT 5.64 1.065 5.81 1.095 ;
      RECT 5.72 0.085 6.09 0.585 ;
      RECT 5.93 1.245 6.1 1.315 ;
      RECT 5.93 1.835 6.1 2.635 ;
      RECT 6.27 0.365 6.73 0.535 ;
      RECT 6.27 0.535 6.44 0.765 ;
      RECT 6.27 1.065 6.44 2.135 ;
      RECT 6.27 2.135 6.52 2.465 ;
      RECT 6.61 0.705 7.16 1.035 ;
      RECT 6.61 1.245 6.8 1.965 ;
      RECT 6.745 2.165 7.63 2.335 ;
      RECT 6.96 0.365 7.5 0.535 ;
      RECT 6.97 1.035 7.16 1.575 ;
      RECT 6.97 1.575 7.29 1.905 ;
      RECT 7.33 0.535 7.5 0.995 ;
      RECT 7.33 0.995 8.395 1.325 ;
      RECT 7.33 1.325 7.63 1.405 ;
      RECT 7.46 1.405 7.63 2.165 ;
      RECT 7.745 0.085 8.115 0.615 ;
      RECT 7.8 1.575 8.735 1.905 ;
      RECT 7.81 2.135 8.115 2.635 ;
      RECT 8.385 0.3 8.735 0.825 ;
      RECT 8.465 1.905 8.735 2.455 ;
      RECT 8.565 0.825 8.735 0.995 ;
      RECT 8.565 0.995 9.265 1.325 ;
      RECT 8.565 1.325 8.735 1.575 ;
      RECT 8.905 0.085 9.075 0.695 ;
      RECT 8.905 1.625 9.08 2.635 ;
      RECT 9.775 0.085 9.945 0.93 ;
      RECT 9.775 1.405 9.945 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.64 1.785 0.81 1.955 ;
      RECT 1.05 0.765 1.22 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.62 1.785 6.79 1.955 ;
      RECT 6.63 0.765 6.8 0.935 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
    LAYER met1 ;
      RECT 0.58 1.755 0.87 1.8 ;
      RECT 0.58 1.8 6.85 1.94 ;
      RECT 0.58 1.94 0.87 1.985 ;
      RECT 0.99 0.735 1.28 0.78 ;
      RECT 0.99 0.78 6.86 0.92 ;
      RECT 0.99 0.92 1.28 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.56 1.755 6.85 1.8 ;
      RECT 6.56 1.94 6.85 1.985 ;
      RECT 6.57 0.735 6.86 0.78 ;
      RECT 6.57 0.92 6.86 0.965 ;
  END
END sky130_fd_sc_hd__sdfxtp_2
MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.795 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.285 0.305 9.615 0.735 ;
        RECT 9.285 0.735 10.955 0.905 ;
        RECT 9.285 1.505 10.955 1.675 ;
        RECT 9.285 1.675 9.615 2.395 ;
        RECT 10.135 0.305 10.465 0.735 ;
        RECT 10.135 1.675 10.465 2.395 ;
        RECT 10.655 0.905 10.955 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.025 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.255 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.085 0.785 3.255 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.52 2.135 0.85 2.635 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.25 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 1.88 2.245 2.21 2.635 ;
      RECT 1.975 0.085 2.305 0.445 ;
      RECT 2.12 0.955 2.465 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.695 2.245 3.59 2.415 ;
      RECT 2.82 0.275 3.595 0.445 ;
      RECT 3.08 1.355 3.275 1.685 ;
      RECT 3.08 1.685 3.25 1.86 ;
      RECT 3.42 1.825 4.385 1.995 ;
      RECT 3.42 1.995 3.59 2.245 ;
      RECT 3.425 0.445 3.595 0.695 ;
      RECT 3.425 0.695 4.385 0.865 ;
      RECT 3.76 2.165 3.93 2.635 ;
      RECT 3.765 0.085 3.965 0.525 ;
      RECT 4.215 0.365 4.565 0.535 ;
      RECT 4.215 0.535 4.385 0.695 ;
      RECT 4.215 0.865 4.385 1.825 ;
      RECT 4.215 1.995 4.385 2.065 ;
      RECT 4.215 2.065 4.45 2.44 ;
      RECT 4.555 0.705 5.135 1.035 ;
      RECT 4.555 1.035 4.795 1.905 ;
      RECT 4.695 2.19 5.765 2.36 ;
      RECT 4.735 0.365 5.475 0.535 ;
      RECT 4.985 1.655 5.425 2.01 ;
      RECT 5.305 0.535 5.475 1.315 ;
      RECT 5.305 1.315 6.105 1.485 ;
      RECT 5.595 1.485 6.105 1.575 ;
      RECT 5.595 1.575 5.765 2.19 ;
      RECT 5.645 0.765 6.445 1.065 ;
      RECT 5.645 1.065 5.815 1.095 ;
      RECT 5.725 0.085 6.095 0.585 ;
      RECT 5.935 1.245 6.105 1.315 ;
      RECT 5.935 1.835 6.105 2.635 ;
      RECT 6.275 0.365 6.735 0.535 ;
      RECT 6.275 0.535 6.445 0.765 ;
      RECT 6.275 1.065 6.445 2.135 ;
      RECT 6.275 2.135 6.525 2.465 ;
      RECT 6.615 0.705 7.165 1.035 ;
      RECT 6.615 1.245 6.805 1.965 ;
      RECT 6.75 2.165 7.635 2.335 ;
      RECT 6.965 0.365 7.505 0.535 ;
      RECT 6.975 1.035 7.165 1.575 ;
      RECT 6.975 1.575 7.295 1.905 ;
      RECT 7.335 0.535 7.505 0.995 ;
      RECT 7.335 0.995 8.4 1.325 ;
      RECT 7.335 1.325 7.635 1.405 ;
      RECT 7.465 1.405 7.635 2.165 ;
      RECT 7.75 0.085 8.12 0.615 ;
      RECT 7.805 1.575 8.755 1.905 ;
      RECT 7.815 2.135 8.12 2.635 ;
      RECT 8.39 0.3 8.75 0.825 ;
      RECT 8.47 1.905 8.755 2.455 ;
      RECT 8.57 0.825 8.75 1.075 ;
      RECT 8.57 1.075 10.485 1.325 ;
      RECT 8.57 1.325 8.755 1.575 ;
      RECT 8.925 0.085 9.095 0.695 ;
      RECT 8.925 1.625 9.105 2.635 ;
      RECT 9.795 0.085 9.965 0.565 ;
      RECT 9.795 1.845 9.965 2.635 ;
      RECT 10.635 0.085 10.805 0.565 ;
      RECT 10.635 1.845 10.805 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.615 1.785 0.785 1.955 ;
      RECT 1.055 0.765 1.225 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.755 0.765 4.925 0.935 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.215 1.785 5.385 1.955 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.625 0.765 6.795 0.935 ;
      RECT 6.625 1.785 6.795 1.955 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.555 1.755 0.845 1.8 ;
      RECT 0.555 1.8 6.855 1.94 ;
      RECT 0.555 1.94 0.845 1.985 ;
      RECT 0.995 0.735 1.285 0.78 ;
      RECT 0.995 0.78 6.855 0.92 ;
      RECT 0.995 0.92 1.285 0.965 ;
      RECT 4.695 0.735 4.985 0.78 ;
      RECT 4.695 0.92 4.985 0.965 ;
      RECT 5.155 1.755 5.445 1.8 ;
      RECT 5.155 1.94 5.445 1.985 ;
      RECT 6.565 0.735 6.855 0.78 ;
      RECT 6.565 0.92 6.855 0.965 ;
      RECT 6.565 1.755 6.855 1.8 ;
      RECT 6.565 1.94 6.855 1.985 ;
  END
END sky130_fd_sc_hd__sdfxtp_4
MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.795 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.255 0.255 9.585 0.79 ;
        RECT 9.255 0.79 9.615 0.825 ;
        RECT 9.255 1.495 9.615 1.53 ;
        RECT 9.255 1.53 9.585 2.43 ;
        RECT 9.41 0.825 9.615 0.89 ;
        RECT 9.41 1.43 9.615 1.495 ;
        RECT 9.445 0.89 9.615 1.43 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.19 0.265 11.44 0.795 ;
        RECT 11.19 1.445 11.44 2.325 ;
        RECT 11.235 0.795 11.44 1.445 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.035 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.255 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.085 0.785 3.255 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 12.15 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.52 2.135 0.85 2.635 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.25 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 1.88 2.245 2.21 2.635 ;
      RECT 1.975 0.085 2.305 0.445 ;
      RECT 2.12 0.955 2.465 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.695 2.245 3.59 2.415 ;
      RECT 2.82 0.275 3.595 0.445 ;
      RECT 3.08 1.355 3.275 1.685 ;
      RECT 3.08 1.685 3.25 1.86 ;
      RECT 3.42 1.825 4.375 1.995 ;
      RECT 3.42 1.995 3.59 2.245 ;
      RECT 3.425 0.445 3.595 0.695 ;
      RECT 3.425 0.695 4.375 0.865 ;
      RECT 3.76 2.165 3.93 2.635 ;
      RECT 3.765 0.085 3.965 0.525 ;
      RECT 4.205 0.365 4.555 0.535 ;
      RECT 4.205 0.535 4.375 0.695 ;
      RECT 4.205 0.865 4.375 1.825 ;
      RECT 4.205 1.995 4.375 2.065 ;
      RECT 4.205 2.065 4.485 2.44 ;
      RECT 4.545 0.705 5.125 1.035 ;
      RECT 4.545 1.035 4.785 1.905 ;
      RECT 4.685 2.19 5.755 2.36 ;
      RECT 4.725 0.365 5.465 0.535 ;
      RECT 4.975 1.655 5.415 2.01 ;
      RECT 5.295 0.535 5.465 1.315 ;
      RECT 5.295 1.315 6.095 1.485 ;
      RECT 5.585 1.485 6.095 1.575 ;
      RECT 5.585 1.575 5.755 2.19 ;
      RECT 5.635 0.765 6.435 1.065 ;
      RECT 5.635 1.065 5.805 1.095 ;
      RECT 5.715 0.085 6.085 0.585 ;
      RECT 5.925 1.245 6.095 1.315 ;
      RECT 5.925 1.835 6.095 2.635 ;
      RECT 6.265 0.365 6.725 0.535 ;
      RECT 6.265 0.535 6.435 0.765 ;
      RECT 6.265 1.065 6.435 2.135 ;
      RECT 6.265 2.135 6.515 2.465 ;
      RECT 6.605 0.705 7.155 1.035 ;
      RECT 6.605 1.245 6.795 1.965 ;
      RECT 6.74 2.165 7.625 2.335 ;
      RECT 6.955 0.365 7.495 0.535 ;
      RECT 6.965 1.035 7.155 1.575 ;
      RECT 6.965 1.575 7.285 1.905 ;
      RECT 7.325 0.535 7.495 0.995 ;
      RECT 7.325 0.995 8.37 1.325 ;
      RECT 7.325 1.325 7.625 1.405 ;
      RECT 7.455 1.405 7.625 2.165 ;
      RECT 7.74 0.085 8.11 0.615 ;
      RECT 7.795 1.575 8.725 1.905 ;
      RECT 7.805 2.135 8.11 2.635 ;
      RECT 8.36 0.3 8.725 0.825 ;
      RECT 8.395 1.905 8.725 2.455 ;
      RECT 8.54 0.825 8.725 0.995 ;
      RECT 8.54 0.995 9.275 1.325 ;
      RECT 8.54 1.325 8.725 1.575 ;
      RECT 8.895 0.085 9.085 0.695 ;
      RECT 8.895 1.625 9.075 2.635 ;
      RECT 9.755 0.085 9.985 0.69 ;
      RECT 9.765 1.615 9.935 2.635 ;
      RECT 10.205 0.345 10.455 0.995 ;
      RECT 10.205 0.995 11.065 1.325 ;
      RECT 10.205 1.325 10.535 2.425 ;
      RECT 10.69 0.085 11.02 0.805 ;
      RECT 10.715 1.495 11.02 2.635 ;
      RECT 11.61 0.085 11.78 0.955 ;
      RECT 11.61 1.395 11.78 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.05 0.765 1.22 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.625 1.785 6.795 1.955 ;
      RECT 6.64 0.765 6.81 0.935 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 6.855 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 0.99 0.735 1.28 0.78 ;
      RECT 0.99 0.78 6.87 0.92 ;
      RECT 0.99 0.92 1.28 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.565 1.755 6.855 1.8 ;
      RECT 6.565 1.94 6.855 1.985 ;
      RECT 6.58 0.735 6.87 0.78 ;
      RECT 6.58 0.92 6.87 0.965 ;
  END
END sky130_fd_sc_hd__sdfxbp_2
MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 1.355 2.775 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.18 0.305 9.53 0.725 ;
        RECT 9.18 0.725 9.56 0.79 ;
        RECT 9.18 0.79 9.61 0.825 ;
        RECT 9.2 1.505 9.61 1.54 ;
        RECT 9.2 1.54 9.53 2.465 ;
        RECT 9.355 1.43 9.61 1.505 ;
        RECT 9.39 0.825 9.61 1.43 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685 0.265 10.94 0.795 ;
        RECT 10.685 1.445 10.94 2.325 ;
        RECT 10.73 0.795 10.94 1.445 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.055 3.995 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.75 3.235 0.785 ;
        RECT 1.76 0.785 2.01 0.81 ;
        RECT 1.76 0.81 1.99 0.82 ;
        RECT 1.76 0.82 1.975 0.835 ;
        RECT 1.76 0.835 1.97 0.84 ;
        RECT 1.76 0.84 1.965 0.85 ;
        RECT 1.76 0.85 1.96 0.855 ;
        RECT 1.76 0.855 1.955 0.86 ;
        RECT 1.76 0.86 1.95 0.87 ;
        RECT 1.76 0.87 1.945 0.875 ;
        RECT 1.76 0.875 1.94 0.88 ;
        RECT 1.76 0.88 1.93 1.685 ;
        RECT 1.79 0.735 3.235 0.75 ;
        RECT 1.805 0.725 3.235 0.735 ;
        RECT 1.82 0.715 3.235 0.725 ;
        RECT 1.83 0.705 3.235 0.715 ;
        RECT 1.84 0.69 3.235 0.705 ;
        RECT 1.86 0.655 3.235 0.69 ;
        RECT 1.875 0.615 3.235 0.655 ;
        RECT 2.455 0.305 2.63 0.615 ;
        RECT 3.065 0.785 3.235 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 11.23 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0 2.635 11.04 2.805 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.515 0.085 0.845 0.465 ;
      RECT 0.515 2.135 0.845 2.635 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.42 0.255 1.705 0.585 ;
      RECT 1.42 0.585 1.59 1.86 ;
      RECT 1.42 1.86 3.23 2.075 ;
      RECT 1.42 2.075 1.705 2.445 ;
      RECT 1.875 2.245 2.205 2.635 ;
      RECT 1.955 0.085 2.285 0.445 ;
      RECT 2.1 0.955 2.445 1.125 ;
      RECT 2.1 1.125 2.27 1.86 ;
      RECT 2.675 2.245 3.57 2.415 ;
      RECT 2.8 0.275 3.575 0.445 ;
      RECT 3.06 1.355 3.255 1.685 ;
      RECT 3.06 1.685 3.23 1.86 ;
      RECT 3.4 1.825 4.335 1.995 ;
      RECT 3.4 1.995 3.57 2.245 ;
      RECT 3.405 0.445 3.575 0.715 ;
      RECT 3.405 0.715 4.335 0.885 ;
      RECT 3.74 2.165 3.91 2.635 ;
      RECT 3.745 0.085 3.945 0.545 ;
      RECT 4.165 0.365 4.515 0.535 ;
      RECT 4.165 0.535 4.335 0.715 ;
      RECT 4.165 0.885 4.335 1.825 ;
      RECT 4.165 1.995 4.335 2.07 ;
      RECT 4.165 2.07 4.45 2.44 ;
      RECT 4.505 0.705 5.085 1.035 ;
      RECT 4.505 1.035 4.745 1.905 ;
      RECT 4.645 2.19 5.715 2.36 ;
      RECT 4.685 0.365 5.425 0.535 ;
      RECT 4.935 1.655 5.375 2.01 ;
      RECT 5.255 0.535 5.425 1.315 ;
      RECT 5.255 1.315 6.055 1.485 ;
      RECT 5.545 1.485 6.055 1.575 ;
      RECT 5.545 1.575 5.715 2.19 ;
      RECT 5.595 0.765 6.395 1.065 ;
      RECT 5.595 1.065 5.765 1.095 ;
      RECT 5.675 0.085 6.045 0.585 ;
      RECT 5.885 1.245 6.055 1.315 ;
      RECT 5.885 1.835 6.055 2.635 ;
      RECT 6.225 0.365 6.685 0.535 ;
      RECT 6.225 0.535 6.395 0.765 ;
      RECT 6.225 1.065 6.395 2.135 ;
      RECT 6.225 2.135 6.475 2.465 ;
      RECT 6.565 0.705 7.115 1.035 ;
      RECT 6.565 1.245 6.755 1.965 ;
      RECT 6.7 2.165 7.585 2.335 ;
      RECT 6.915 0.365 7.455 0.535 ;
      RECT 6.925 1.035 7.115 1.575 ;
      RECT 6.925 1.575 7.245 1.905 ;
      RECT 7.285 0.535 7.455 0.995 ;
      RECT 7.285 0.995 8.315 1.325 ;
      RECT 7.285 1.325 7.585 1.405 ;
      RECT 7.415 1.405 7.585 2.165 ;
      RECT 7.7 0.085 8.07 0.615 ;
      RECT 7.755 1.575 8.67 1.905 ;
      RECT 7.765 2.135 8.07 2.635 ;
      RECT 8.34 0.3 8.67 0.825 ;
      RECT 8.38 1.905 8.67 2.455 ;
      RECT 8.485 0.825 8.67 0.995 ;
      RECT 8.485 0.995 9.22 1.325 ;
      RECT 8.485 1.325 8.67 1.575 ;
      RECT 8.84 0.085 9.01 0.695 ;
      RECT 8.84 1.625 9.01 2.635 ;
      RECT 9.7 0.345 9.95 0.62 ;
      RECT 9.7 1.685 10.03 2.425 ;
      RECT 9.78 0.62 9.95 0.995 ;
      RECT 9.78 0.995 10.56 1.325 ;
      RECT 9.78 1.325 10.03 1.685 ;
      RECT 10.185 0.085 10.515 0.805 ;
      RECT 10.21 1.495 10.515 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.015 0.765 1.185 0.935 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.165 1.785 5.335 1.955 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.575 1.785 6.745 1.955 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 0.765 6.755 0.935 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 6.805 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 0.955 0.735 1.245 0.78 ;
      RECT 0.955 0.78 6.815 0.92 ;
      RECT 0.955 0.92 1.245 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.105 1.755 5.395 1.8 ;
      RECT 5.105 1.94 5.395 1.985 ;
      RECT 6.515 1.755 6.805 1.8 ;
      RECT 6.515 1.94 6.805 1.985 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
  END
END sky130_fd_sc_hd__sdfxbp_1
MACRO sky130_fd_sc_hd__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465 0.985 3.715 1.445 ;
        RECT 3.465 1.445 5.29 1.675 ;
        RECT 4.895 0.995 5.29 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.97 1.015 4.725 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185 1.03 2.855 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.045 0.455 1.445 ;
        RECT 0.125 1.445 1.8 1.68 ;
        RECT 1.615 1.03 1.975 1.275 ;
        RECT 1.615 1.275 1.8 1.445 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755 1.075 1.425 1.275 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.212750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.255 0.38 0.615 ;
        RECT 0.12 0.615 5.355 0.805 ;
        RECT 0.12 0.805 3.255 0.845 ;
        RECT 0.9 1.85 2.14 2.105 ;
        RECT 1.05 0.255 1.295 0.615 ;
        RECT 1.965 0.255 2.295 0.615 ;
        RECT 1.97 1.445 3.255 1.625 ;
        RECT 1.97 1.625 2.14 1.85 ;
        RECT 2.965 0.275 3.295 0.615 ;
        RECT 3.025 0.845 3.255 1.445 ;
        RECT 5.02 0.295 5.355 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 5.71 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.52 0.085 ;
      RECT 0 2.635 5.52 2.805 ;
      RECT 0.1 1.87 0.46 2.275 ;
      RECT 0.1 2.275 2.185 2.295 ;
      RECT 0.1 2.295 2.985 2.465 ;
      RECT 0.55 0.085 0.88 0.445 ;
      RECT 1.465 0.085 1.795 0.445 ;
      RECT 2.31 1.795 3.335 1.845 ;
      RECT 2.31 1.845 5.4 1.965 ;
      RECT 2.31 1.965 2.64 2.06 ;
      RECT 2.465 0.085 2.795 0.445 ;
      RECT 2.815 2.135 2.985 2.295 ;
      RECT 3.155 1.965 5.4 2.095 ;
      RECT 3.155 2.095 3.52 2.465 ;
      RECT 3.69 2.275 4.02 2.635 ;
      RECT 4.125 0.085 4.455 0.445 ;
      RECT 4.19 2.095 5.4 2.105 ;
      RECT 4.19 2.105 4.4 2.465 ;
      RECT 4.57 2.275 4.9 2.635 ;
      RECT 5.07 2.105 5.4 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
  END
END sky130_fd_sc_hd__a2111oi_2
MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.02 7.745 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.96 1.02 9.99 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955 1.02 5.65 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.02 3.745 1.275 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495 1.02 1.845 1.275 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.009500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.615 7.62 0.785 ;
        RECT 0.145 0.785 0.32 1.475 ;
        RECT 0.145 1.475 1.72 1.655 ;
        RECT 0.53 1.655 1.72 1.685 ;
        RECT 0.53 1.685 0.86 2.085 ;
        RECT 0.615 0.455 0.79 0.615 ;
        RECT 1.39 1.685 1.72 2.085 ;
        RECT 1.46 0.455 1.65 0.615 ;
        RECT 2.4 0.455 2.59 0.615 ;
        RECT 3.26 0.455 3.51 0.615 ;
        RECT 4.18 0.455 4.42 0.615 ;
        RECT 5.09 0.455 5.275 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 10.31 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.12 0.085 ;
      RECT 0 2.635 10.12 2.805 ;
      RECT 0.1 1.835 0.36 2.255 ;
      RECT 0.1 2.255 3.87 2.445 ;
      RECT 0.115 0.085 0.445 0.445 ;
      RECT 0.96 0.085 1.29 0.445 ;
      RECT 1.03 1.855 1.22 2.255 ;
      RECT 1.82 0.085 2.23 0.445 ;
      RECT 1.89 1.855 2.08 2.255 ;
      RECT 2.25 1.475 5.68 1.655 ;
      RECT 2.25 1.655 3.44 1.685 ;
      RECT 2.25 1.685 2.58 2.085 ;
      RECT 2.75 1.855 2.94 2.255 ;
      RECT 2.76 0.085 3.09 0.445 ;
      RECT 3.11 1.685 3.44 2.085 ;
      RECT 3.61 1.835 3.87 2.255 ;
      RECT 3.68 0.085 4.01 0.445 ;
      RECT 4.06 1.835 4.32 2.255 ;
      RECT 4.06 2.255 5.18 2.275 ;
      RECT 4.06 2.275 6.05 2.445 ;
      RECT 4.49 1.655 5.68 1.685 ;
      RECT 4.49 1.685 4.82 2.085 ;
      RECT 4.59 0.085 4.92 0.445 ;
      RECT 4.99 1.855 5.18 2.255 ;
      RECT 5.35 1.685 5.68 2.085 ;
      RECT 5.445 0.085 5.78 0.445 ;
      RECT 5.86 1.445 9.77 1.615 ;
      RECT 5.86 1.615 6.05 2.275 ;
      RECT 5.98 0.275 8.075 0.445 ;
      RECT 6.22 1.785 6.55 2.635 ;
      RECT 6.72 1.615 6.91 2.315 ;
      RECT 7.08 1.805 7.41 2.635 ;
      RECT 7.58 1.615 9.77 1.665 ;
      RECT 7.58 1.665 7.91 2.315 ;
      RECT 7.885 0.445 8.075 0.615 ;
      RECT 7.885 0.615 9.865 0.785 ;
      RECT 8.08 1.895 8.41 2.635 ;
      RECT 8.245 0.085 8.575 0.445 ;
      RECT 8.58 1.665 9.77 1.67 ;
      RECT 8.58 1.67 8.84 2.29 ;
      RECT 8.745 0.3 8.935 0.615 ;
      RECT 9.03 1.915 9.36 2.635 ;
      RECT 9.105 0.085 9.435 0.445 ;
      RECT 9.53 1.67 9.77 2.26 ;
      RECT 9.605 0.29 9.865 0.615 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
  END
END sky130_fd_sc_hd__a2111oi_4
MACRO sky130_fd_sc_hd__a2111oi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.07 2.625 1.4 ;
        RECT 2.355 0.66 2.625 1.07 ;
        RECT 2.355 1.4 2.625 1.735 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795 0.65 3.135 1.735 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.055 1.845 1.735 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.055 1.325 2.36 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.73 0.435 1.655 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.424000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.825 0.785 2.465 ;
        RECT 0.605 0.635 2.04 0.885 ;
        RECT 0.605 0.885 0.785 1.825 ;
        RECT 0.785 0.255 1.04 0.615 ;
        RECT 0.785 0.615 2.04 0.635 ;
        RECT 1.71 0.28 2.04 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.41 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.22 0.085 ;
      RECT 0 2.635 3.22 2.805 ;
      RECT 0.285 0.085 0.615 0.465 ;
      RECT 1.21 0.085 1.54 0.445 ;
      RECT 1.54 1.905 2.87 2.085 ;
      RECT 1.54 2.085 1.87 2.465 ;
      RECT 2.04 2.255 2.37 2.635 ;
      RECT 2.47 0.085 2.8 0.48 ;
      RECT 2.54 2.085 2.87 2.465 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
  END
END sky130_fd_sc_hd__a2111oi_0
MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.725 1.4 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.35 3.09 1.02 ;
        RECT 2.905 1.02 3.54 1.29 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.05 2.27 1.4 ;
        RECT 1.94 1.4 2.215 2.455 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.05 1.77 2.455 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785 1.05 1.235 2.455 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.388750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.7 1.375 0.705 ;
        RECT 0.145 0.705 2.42 0.815 ;
        RECT 0.145 0.815 2.3 0.88 ;
        RECT 0.145 0.88 0.53 2.46 ;
        RECT 1.045 0.26 1.375 0.7 ;
        RECT 2.09 0.305 2.42 0.705 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975 -0.065 2.145 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.315 0.085 0.63 0.525 ;
      RECT 1.55 0.085 1.88 0.535 ;
      RECT 2.395 1.58 3.505 1.75 ;
      RECT 2.395 1.75 2.625 2.46 ;
      RECT 2.8 1.92 3.13 2.635 ;
      RECT 3.27 0.085 3.51 0.76 ;
      RECT 3.31 1.75 3.505 2.46 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a2111oi_1
MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.075 2.69 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.075 4.3 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.445 1.285 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.255 1.285 0.725 ;
        RECT 0.955 0.725 6.76 0.905 ;
        RECT 1.795 0.255 2.125 0.725 ;
        RECT 3.155 0.255 3.485 0.725 ;
        RECT 3.995 0.255 4.325 0.725 ;
        RECT 4.835 0.255 5.165 0.725 ;
        RECT 4.875 1.455 6.76 1.625 ;
        RECT 4.875 1.625 5.125 2.125 ;
        RECT 5.675 0.255 6.005 0.725 ;
        RECT 5.715 1.625 5.965 2.125 ;
        RECT 6.42 0.905 6.76 1.455 ;
        RECT 6.515 0.315 6.76 0.725 ;
        RECT 6.555 1.625 6.76 2.415 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 7.09 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 0.11 0.255 0.445 0.735 ;
      RECT 0.11 0.735 0.785 0.905 ;
      RECT 0.11 1.455 4.705 1.625 ;
      RECT 0.11 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.615 0.085 0.785 0.555 ;
      RECT 0.615 0.905 0.785 1.455 ;
      RECT 0.995 1.795 4.285 1.965 ;
      RECT 0.995 1.965 1.245 2.465 ;
      RECT 1.415 2.135 1.665 2.635 ;
      RECT 1.455 0.085 1.625 0.555 ;
      RECT 1.835 1.965 2.085 2.465 ;
      RECT 2.255 2.135 2.505 2.635 ;
      RECT 2.295 0.085 2.985 0.555 ;
      RECT 2.775 2.135 3.025 2.295 ;
      RECT 2.775 2.295 6.385 2.465 ;
      RECT 3.195 1.965 3.445 2.125 ;
      RECT 3.615 2.135 3.865 2.295 ;
      RECT 3.655 0.085 3.825 0.555 ;
      RECT 4.035 1.965 4.285 2.125 ;
      RECT 4.455 1.795 4.705 2.295 ;
      RECT 4.495 0.085 4.665 0.555 ;
      RECT 4.535 1.075 6.125 1.285 ;
      RECT 4.535 1.285 4.705 1.455 ;
      RECT 5.295 1.795 5.545 2.295 ;
      RECT 5.335 0.085 5.505 0.555 ;
      RECT 6.135 1.795 6.385 2.295 ;
      RECT 6.175 0.085 6.345 0.555 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
  END
END sky130_fd_sc_hd__nor3b_4
MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.64 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.03 1.075 4.515 1.285 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.105 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 2.815 0.905 3.065 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.15 -0.085 0.32 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 4.79 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.6 0.085 ;
      RECT 0 2.635 4.6 2.805 ;
      RECT 0.09 0.085 0.365 0.905 ;
      RECT 0.09 1.455 2.085 1.625 ;
      RECT 0.09 1.625 0.405 2.465 ;
      RECT 0.575 1.795 0.825 2.635 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.035 0.085 1.205 0.555 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.48 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 1.875 0.085 2.605 0.555 ;
      RECT 2.375 1.455 2.645 2.295 ;
      RECT 3.235 1.075 3.86 1.285 ;
      RECT 3.235 1.455 3.48 2.295 ;
      RECT 3.275 0.085 3.48 0.895 ;
      RECT 3.69 0.38 4.045 0.905 ;
      RECT 3.69 0.905 3.86 1.075 ;
      RECT 3.69 1.285 3.86 1.455 ;
      RECT 3.69 1.455 4.045 1.87 ;
      RECT 4.215 0.085 4.505 0.825 ;
      RECT 4.215 1.54 4.465 2.635 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
  END
END sky130_fd_sc_hd__nor3b_2
MACRO sky130_fd_sc_hd__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.815 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.995 1.305 1.615 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.335 1.615 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.716500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 0.655 ;
        RECT 0.085 0.655 1.445 0.825 ;
        RECT 0.085 0.825 0.255 1.445 ;
        RECT 0.085 1.445 0.545 2.455 ;
        RECT 1.275 0.31 1.445 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 2.95 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.76 0.085 ;
      RECT 0 2.635 2.76 2.805 ;
      RECT 0.425 1.075 0.885 1.245 ;
      RECT 0.715 1.245 0.885 1.785 ;
      RECT 0.715 1.785 2.675 1.955 ;
      RECT 0.775 0.085 1.105 0.485 ;
      RECT 1.615 0.085 1.945 0.825 ;
      RECT 1.615 2.125 1.945 2.635 ;
      RECT 2.18 0.405 2.35 0.655 ;
      RECT 2.18 0.655 2.675 0.825 ;
      RECT 2.505 0.825 2.675 1.785 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
  END
END sky130_fd_sc_hd__nor3b_1
MACRO sky130_fd_sc_hd__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a222oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1 2.925 1.33 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1 3.435 1.33 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135 1 2.445 1.33 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 1 1.965 1.33 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1 0.545 1.315 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.715 1 1.085 1.315 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  0.897600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.255 0.425 0.645 ;
        RECT 0.095 0.645 2.645 0.815 ;
        RECT 0.095 1.485 0.425 1.5 ;
        RECT 0.095 1.5 1.425 1.67 ;
        RECT 0.095 1.67 0.425 1.68 ;
        RECT 0.095 1.68 0.345 2.255 ;
        RECT 0.095 2.255 0.425 2.465 ;
        RECT 1.015 1.67 1.185 1.83 ;
        RECT 1.255 0.815 1.48 1.33 ;
        RECT 1.255 1.33 1.425 1.5 ;
        RECT 2.315 0.295 2.645 0.645 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 3.68 0.24 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.19 1.305 3.87 2.91 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.68 0.085 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0.515 1.875 0.845 2.075 ;
      RECT 0.595 2.075 0.765 2.295 ;
      RECT 0.595 2.295 2.185 2.465 ;
      RECT 0.875 0.085 1.605 0.465 ;
      RECT 1.515 1.825 2.015 1.965 ;
      RECT 1.515 1.965 1.97 1.97 ;
      RECT 1.515 1.97 1.935 1.98 ;
      RECT 1.515 1.98 1.915 1.995 ;
      RECT 1.845 1.655 3.595 1.67 ;
      RECT 1.845 1.67 2.685 1.735 ;
      RECT 1.845 1.735 2.605 1.825 ;
      RECT 2.015 2.135 2.185 2.295 ;
      RECT 2.355 1.5 3.595 1.655 ;
      RECT 2.355 1.825 2.605 2.255 ;
      RECT 2.355 2.255 2.685 2.465 ;
      RECT 2.775 1.905 3.105 2.075 ;
      RECT 2.855 2.075 3.025 2.635 ;
      RECT 3.22 1.67 3.595 1.735 ;
      RECT 3.255 0.085 3.585 0.815 ;
      RECT 3.255 2.255 3.595 2.465 ;
      RECT 3.335 1.735 3.595 2.255 ;
    LAYER mcon ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
  END
END sky130_fd_sc_hd__a222oi_1

MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END G_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.220000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 21.490000 145.315000 ;
      RECT 11.095000 145.315000 12.220000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.015000 ;
      RECT 11.275000  26.015000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.575000 ;
      RECT 11.275000  81.575000 23.280000  82.085000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.640000 100.865000 68.495000 101.035000 ;
      RECT 20.640000 101.035000 21.490000 109.275000 ;
      RECT 20.640000 109.275000 68.495000 109.445000 ;
      RECT 20.640000 109.445000 21.490000 117.770000 ;
      RECT 20.640000 117.770000 68.495000 117.940000 ;
      RECT 20.640000 117.940000 21.490000 144.465000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.085000 23.280000  82.180000 ;
      RECT 22.430000  82.180000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.770000  97.890000 23.280000  98.990000 ;
      RECT 22.770000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.015000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.325000 72.000000 195.000000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.950000   3.000000 72.000000   6.330000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   9.705000 11.735000   9.715000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   9.705000 11.735000   9.710000 ;
      RECT 10.710000   9.710000 11.735000   9.715000 ;
      RECT 10.710000   9.715000 11.515000   9.935000 ;
      RECT 10.720000   8.145000 11.720000   8.160000 ;
      RECT 10.780000   9.715000 11.665000   9.785000 ;
      RECT 10.790000   8.075000 11.650000   8.145000 ;
      RECT 10.850000   9.785000 11.595000   9.855000 ;
      RECT 10.860000   8.005000 11.580000   8.075000 ;
      RECT 10.920000   9.855000 11.525000   9.925000 ;
      RECT 10.930000   7.935000 11.510000   8.005000 ;
      RECT 10.930000   7.935000 11.735000   8.160000 ;
      RECT 10.930000   9.925000 11.515000   9.935000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.860000  25.500000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.500000 65.860000  29.820000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.555000 65.720000  29.765000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.820000 64.810000  30.870000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.750000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.750000 65.860000  39.875000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.805000 65.720000  39.820000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.875000 64.885000  40.850000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.730000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.730000 65.860000  49.895000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.785000 65.720000  49.840000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.895000 64.885000  50.870000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.745000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.745000 65.855000  59.880000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.800000 65.715000  59.825000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.880000 64.885000  60.850000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.735000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.735000 65.855000  69.880000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.795000 65.715000  69.825000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.880000 64.885000  70.850000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.550000  74.180000 ;
      RECT 14.030000  73.910000 65.085000  73.980000 ;
      RECT 14.030000  73.980000 65.155000  74.050000 ;
      RECT 14.030000  74.050000 65.225000  74.120000 ;
      RECT 14.030000  74.120000 65.295000  74.180000 ;
      RECT 14.030000  74.180000 65.760000  74.390000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.100000  74.180000 65.350000  74.250000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.170000  74.250000 65.425000  74.320000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.860000  74.490000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.490000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.545000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.820000 ;
      RECT 14.240000  98.840000 75.000000 129.820000 ;
      RECT 14.240000 129.820000 75.000000 130.705000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 139.825000 75.000000 140.710000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 149.825000 75.000000 150.710000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 159.825000 75.000000 160.710000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 169.825000 75.000000 170.710000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 179.825000 75.000000 180.710000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 189.825000 75.000000 190.710000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 134.795000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 144.795000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 154.795000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 164.795000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 174.795000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 184.795000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.520000 130.705000 75.000000 130.845000 ;
      RECT 15.520000 140.710000 75.000000 140.850000 ;
      RECT 15.520000 150.710000 75.000000 150.850000 ;
      RECT 15.520000 160.710000 75.000000 160.850000 ;
      RECT 15.520000 170.710000 75.000000 170.850000 ;
      RECT 15.520000 180.710000 75.000000 180.850000 ;
      RECT 15.520000 190.710000 75.000000 190.850000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.660000 133.770000 75.000000 133.910000 ;
      RECT 15.660000 143.770000 75.000000 143.910000 ;
      RECT 15.660000 153.770000 75.000000 153.910000 ;
      RECT 15.660000 163.770000 75.000000 163.910000 ;
      RECT 15.660000 173.770000 75.000000 173.910000 ;
      RECT 15.660000 183.770000 75.000000 183.910000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.140000   5.235000 17.350000   9.250000 ;
      RECT 17.140000   5.235000 17.490000   9.250000 ;
      RECT 17.140000   9.250000 17.490000   9.600000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.210000   5.165000 17.350000   5.235000 ;
      RECT 17.210000   9.250000 17.350000   9.320000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.280000   5.095000 17.350000   5.165000 ;
      RECT 17.280000   9.320000 17.350000   9.390000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.320000   5.055000 17.490000   5.235000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 65.660000  25.300000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.570000   9.680000 55.880000   9.800000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.580000 193.770000 75.000000 193.910000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.400000  19.930000 53.955000  21.835000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.600000 ;
      RECT 20.775000   1.600000 20.785000   1.760000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.555000  17.775000 53.955000  19.930000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 56.110000  17.775000 ;
      RECT 53.675000   0.000000 53.955000   7.875000 ;
      RECT 53.675000   7.875000 55.760000   9.680000 ;
      RECT 53.815000   8.000000 53.885000   8.070000 ;
      RECT 53.815000   8.070000 53.955000   8.140000 ;
      RECT 53.815000   8.140000 54.025000   8.210000 ;
      RECT 53.815000   8.210000 54.095000   8.280000 ;
      RECT 53.815000   8.280000 54.165000   8.350000 ;
      RECT 53.815000   8.350000 54.235000   8.420000 ;
      RECT 53.815000   8.420000 54.305000   8.490000 ;
      RECT 53.815000   8.490000 54.375000   8.560000 ;
      RECT 53.815000   8.560000 54.445000   8.630000 ;
      RECT 53.815000   8.630000 54.515000   8.700000 ;
      RECT 53.815000   8.700000 54.585000   8.770000 ;
      RECT 53.815000   8.770000 54.655000   8.840000 ;
      RECT 53.815000   8.840000 54.725000   8.910000 ;
      RECT 53.815000   8.910000 54.795000   8.980000 ;
      RECT 53.815000   8.980000 54.865000   9.050000 ;
      RECT 53.815000   9.050000 54.935000   9.120000 ;
      RECT 53.815000   9.120000 55.005000   9.190000 ;
      RECT 53.815000   9.190000 55.075000   9.260000 ;
      RECT 53.815000   9.260000 55.145000   9.330000 ;
      RECT 53.815000   9.330000 55.215000   9.400000 ;
      RECT 53.815000   9.400000 55.285000   9.470000 ;
      RECT 53.815000   9.470000 55.355000   9.540000 ;
      RECT 53.815000   9.540000 55.425000   9.610000 ;
      RECT 53.815000   9.610000 55.495000   9.680000 ;
      RECT 53.815000   9.680000 55.565000   9.750000 ;
      RECT 53.815000   9.750000 55.635000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.030000 ;
      RECT 55.875000  10.030000 56.110000  17.360000 ;
      RECT 68.150000  74.490000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.545000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.865000  73.770000 75.000000  74.490000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.385000 15.205000 171.495000 ;
      RECT 13.300000  94.425000 15.205000 171.595000 ;
      RECT 13.440000  94.145000 15.205000  94.385000 ;
      RECT 13.440000  94.285000 15.205000  94.425000 ;
      RECT 13.580000  94.145000 15.205000  94.285000 ;
      RECT 13.725000  94.000000 15.205000  94.145000 ;
      RECT 13.875000  93.850000 15.350000  94.000000 ;
      RECT 14.025000  93.700000 15.500000  93.850000 ;
      RECT 14.175000  93.550000 15.650000  93.700000 ;
      RECT 14.325000  93.400000 15.800000  93.550000 ;
      RECT 14.475000  93.250000 15.950000  93.400000 ;
      RECT 14.625000  93.100000 16.100000  93.250000 ;
      RECT 14.775000  92.950000 16.250000  93.100000 ;
      RECT 14.925000  92.800000 16.400000  92.950000 ;
      RECT 15.075000  92.650000 16.550000  92.800000 ;
      RECT 15.225000  92.500000 16.700000  92.650000 ;
      RECT 15.375000  92.350000 16.850000  92.500000 ;
      RECT 15.525000  92.200000 17.000000  92.350000 ;
      RECT 15.675000  92.050000 17.150000  92.200000 ;
      RECT 15.825000  91.900000 17.300000  92.050000 ;
      RECT 15.975000  91.750000 17.450000  91.900000 ;
      RECT 16.125000  91.600000 17.600000  91.750000 ;
      RECT 16.275000  91.450000 17.750000  91.600000 ;
      RECT 16.425000  91.300000 17.900000  91.450000 ;
      RECT 16.575000  91.150000 18.050000  91.300000 ;
      RECT 16.725000  91.000000 18.200000  91.150000 ;
      RECT 16.875000  90.850000 18.350000  91.000000 ;
      RECT 17.025000  90.700000 18.500000  90.850000 ;
      RECT 17.175000  90.550000 18.650000  90.700000 ;
      RECT 17.325000  90.400000 18.800000  90.550000 ;
      RECT 17.475000  90.250000 18.950000  90.400000 ;
      RECT 17.625000  90.100000 19.100000  90.250000 ;
      RECT 17.775000  89.950000 19.250000  90.100000 ;
      RECT 17.925000  89.800000 19.400000  89.950000 ;
      RECT 18.075000  89.650000 19.550000  89.800000 ;
      RECT 18.225000  89.500000 19.700000  89.650000 ;
      RECT 18.375000  89.350000 19.850000  89.500000 ;
      RECT 18.525000  89.200000 20.000000  89.350000 ;
      RECT 18.675000  89.050000 20.150000  89.200000 ;
      RECT 18.825000  88.900000 20.300000  89.050000 ;
      RECT 18.975000  88.750000 20.450000  88.900000 ;
      RECT 19.125000  88.600000 20.600000  88.750000 ;
      RECT 19.275000  88.450000 20.750000  88.600000 ;
      RECT 19.425000  88.300000 20.900000  88.450000 ;
      RECT 19.575000  88.150000 21.050000  88.300000 ;
      RECT 19.725000  88.000000 21.200000  88.150000 ;
      RECT 19.875000  87.850000 21.350000  88.000000 ;
      RECT 20.025000  87.700000 21.500000  87.850000 ;
      RECT 20.175000  87.550000 21.650000  87.700000 ;
      RECT 20.325000  87.400000 21.800000  87.550000 ;
      RECT 20.475000  87.250000 21.950000  87.400000 ;
      RECT 20.625000  87.100000 22.100000  87.250000 ;
      RECT 20.775000  86.950000 22.250000  87.100000 ;
      RECT 20.925000  86.800000 22.400000  86.950000 ;
      RECT 21.075000  86.650000 22.550000  86.800000 ;
      RECT 21.225000  86.500000 22.700000  86.650000 ;
      RECT 21.375000  86.350000 22.850000  86.500000 ;
      RECT 21.525000  86.200000 23.000000  86.350000 ;
      RECT 21.675000  86.050000 23.150000  86.200000 ;
      RECT 21.825000  85.900000 23.300000  86.050000 ;
      RECT 21.950000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000 166.935000 25.635000 170.445000 ;
      RECT 22.075000  96.885000 25.635000  96.955000 ;
      RECT 22.100000  85.625000 23.450000  85.775000 ;
      RECT 22.155000 166.935000 25.635000 167.085000 ;
      RECT 22.225000  96.735000 25.635000  96.885000 ;
      RECT 22.250000  85.475000 23.450000  85.625000 ;
      RECT 22.305000 167.085000 25.635000 167.235000 ;
      RECT 22.375000  96.585000 25.635000  96.735000 ;
      RECT 22.400000  85.325000 23.450000  85.475000 ;
      RECT 22.455000 167.235000 25.635000 167.385000 ;
      RECT 22.525000  96.435000 25.635000  96.585000 ;
      RECT 22.550000  85.175000 23.450000  85.325000 ;
      RECT 22.605000 167.385000 25.635000 167.535000 ;
      RECT 22.675000  96.285000 25.635000  96.435000 ;
      RECT 22.700000  85.025000 23.450000  85.175000 ;
      RECT 22.755000 167.535000 25.635000 167.685000 ;
      RECT 22.825000  96.135000 25.635000  96.285000 ;
      RECT 22.850000  84.875000 23.450000  85.025000 ;
      RECT 22.905000 167.685000 25.635000 167.835000 ;
      RECT 22.975000  95.985000 25.635000  96.135000 ;
      RECT 23.000000  84.725000 23.450000  84.875000 ;
      RECT 23.055000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.485000 23.450000  85.900000 ;
      RECT 23.125000  95.835000 25.635000  95.985000 ;
      RECT 23.150000  84.575000 23.450000  84.725000 ;
      RECT 23.205000 167.985000 25.635000 168.135000 ;
      RECT 23.275000  95.685000 25.635000  95.835000 ;
      RECT 23.300000  84.425000 23.450000  84.575000 ;
      RECT 23.355000 168.135000 25.635000 168.285000 ;
      RECT 23.425000  95.535000 25.635000  95.685000 ;
      RECT 23.505000 168.285000 25.635000 168.435000 ;
      RECT 23.575000  95.385000 25.635000  95.535000 ;
      RECT 23.655000 168.435000 25.635000 168.585000 ;
      RECT 23.725000  95.235000 25.635000  95.385000 ;
      RECT 23.805000 168.585000 25.635000 168.735000 ;
      RECT 23.875000  95.085000 25.635000  95.235000 ;
      RECT 23.955000 168.735000 25.635000 168.885000 ;
      RECT 24.025000  94.935000 25.635000  95.085000 ;
      RECT 24.105000 168.885000 25.635000 169.035000 ;
      RECT 24.175000  94.785000 25.635000  94.935000 ;
      RECT 24.255000 169.035000 25.635000 169.185000 ;
      RECT 24.325000  94.635000 25.635000  94.785000 ;
      RECT 24.405000 169.185000 25.635000 169.335000 ;
      RECT 24.475000  94.485000 25.635000  94.635000 ;
      RECT 24.555000 169.335000 25.635000 169.485000 ;
      RECT 24.625000  94.335000 25.635000  94.485000 ;
      RECT 24.625000  94.335000 25.635000  96.955000 ;
      RECT 24.705000 169.485000 25.635000 169.635000 ;
      RECT 24.745000  94.215000 25.635000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.335000 ;
      RECT 24.800000  82.335000 25.150000  82.785000 ;
      RECT 24.855000 169.635000 25.635000 169.785000 ;
      RECT 24.895000  94.065000 25.755000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.335000 ;
      RECT 24.900000  82.335000 25.450000  82.485000 ;
      RECT 24.900000  82.485000 25.300000  82.635000 ;
      RECT 24.900000  82.635000 25.150000  82.785000 ;
      RECT 24.900000  82.785000 25.000000  82.935000 ;
      RECT 25.005000 169.785000 25.635000 169.935000 ;
      RECT 25.045000  93.915000 25.905000  94.065000 ;
      RECT 25.155000 169.935000 25.635000 170.085000 ;
      RECT 25.195000  93.765000 26.055000  93.915000 ;
      RECT 25.305000 170.085000 25.635000 170.235000 ;
      RECT 25.345000  93.615000 26.205000  93.765000 ;
      RECT 25.455000 170.235000 25.635000 170.385000 ;
      RECT 25.495000  93.465000 26.355000  93.615000 ;
      RECT 25.515000 170.445000 25.635000 189.915000 ;
      RECT 25.605000 170.385000 25.635000 170.535000 ;
      RECT 25.645000  93.315000 26.505000  93.465000 ;
      RECT 25.795000  93.165000 26.655000  93.315000 ;
      RECT 25.945000  93.015000 26.805000  93.165000 ;
      RECT 26.095000  92.865000 26.955000  93.015000 ;
      RECT 26.245000  92.715000 27.105000  92.865000 ;
      RECT 26.395000  92.565000 27.255000  92.715000 ;
      RECT 26.545000  92.415000 27.405000  92.565000 ;
      RECT 26.695000  92.265000 27.555000  92.415000 ;
      RECT 26.845000  92.115000 27.705000  92.265000 ;
      RECT 26.995000  91.965000 27.855000  92.115000 ;
      RECT 27.145000  91.815000 28.005000  91.965000 ;
      RECT 27.295000  91.665000 28.155000  91.815000 ;
      RECT 27.445000  91.515000 28.305000  91.665000 ;
      RECT 27.595000  91.365000 28.455000  91.515000 ;
      RECT 27.745000  91.215000 28.605000  91.365000 ;
      RECT 27.895000  91.065000 28.755000  91.215000 ;
      RECT 28.045000  90.915000 28.905000  91.065000 ;
      RECT 28.195000  90.765000 29.055000  90.915000 ;
      RECT 28.345000  90.615000 29.205000  90.765000 ;
      RECT 28.495000  90.465000 29.355000  90.615000 ;
      RECT 28.645000  90.315000 29.505000  90.465000 ;
      RECT 28.795000  90.165000 29.655000  90.315000 ;
      RECT 28.945000  90.015000 29.805000  90.165000 ;
      RECT 29.095000  89.865000 29.955000  90.015000 ;
      RECT 29.245000  89.715000 30.105000  89.865000 ;
      RECT 29.395000  89.565000 30.255000  89.715000 ;
      RECT 29.545000  89.415000 30.405000  89.565000 ;
      RECT 29.695000  89.265000 30.555000  89.415000 ;
      RECT 29.845000  89.115000 30.705000  89.265000 ;
      RECT 29.995000  88.965000 30.855000  89.115000 ;
      RECT 30.145000  88.815000 31.005000  88.965000 ;
      RECT 30.295000  88.665000 31.155000  88.815000 ;
      RECT 30.445000  88.515000 31.305000  88.665000 ;
      RECT 30.595000  88.365000 31.455000  88.515000 ;
      RECT 30.745000  88.215000 31.605000  88.365000 ;
      RECT 30.895000  88.065000 31.755000  88.215000 ;
      RECT 31.045000  87.915000 31.905000  88.065000 ;
      RECT 31.195000  87.765000 32.055000  87.915000 ;
      RECT 31.345000  87.615000 32.205000  87.765000 ;
      RECT 31.495000  87.465000 32.355000  87.615000 ;
      RECT 31.645000  87.315000 32.505000  87.465000 ;
      RECT 31.795000  87.165000 32.655000  87.315000 ;
      RECT 31.945000  87.015000 32.805000  87.165000 ;
      RECT 32.095000  86.865000 32.955000  87.015000 ;
      RECT 32.245000  86.715000 33.105000  86.865000 ;
      RECT 32.395000  86.565000 33.255000  86.715000 ;
      RECT 32.435000  93.555000 40.410000  93.705000 ;
      RECT 32.435000  93.555000 42.435000  95.580000 ;
      RECT 32.435000  93.705000 40.560000  93.855000 ;
      RECT 32.435000  93.855000 40.710000  94.005000 ;
      RECT 32.435000  94.005000 40.860000  94.155000 ;
      RECT 32.435000  94.155000 41.010000  94.305000 ;
      RECT 32.435000  94.305000 41.160000  94.455000 ;
      RECT 32.435000  94.455000 41.310000  94.605000 ;
      RECT 32.435000  94.605000 41.460000  94.755000 ;
      RECT 32.435000  94.755000 41.610000  94.905000 ;
      RECT 32.435000  94.905000 41.760000  95.055000 ;
      RECT 32.435000  95.055000 41.910000  95.205000 ;
      RECT 32.435000  95.205000 42.060000  95.355000 ;
      RECT 32.435000  95.355000 42.210000  95.505000 ;
      RECT 32.435000  95.505000 42.360000  95.580000 ;
      RECT 32.435000  95.580000 35.440000 159.400000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000 159.400000 36.680000 162.405000 ;
      RECT 32.435000 162.405000 42.435000 163.970000 ;
      RECT 32.515000  93.475000 40.330000  93.555000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  85.865000 33.555000  86.415000 ;
      RECT 32.545000  85.865000 33.955000  86.015000 ;
      RECT 32.545000  86.015000 33.805000  86.165000 ;
      RECT 32.545000  86.165000 33.655000  86.315000 ;
      RECT 32.545000  86.315000 33.555000  86.415000 ;
      RECT 32.545000  86.415000 33.405000  86.565000 ;
      RECT 32.570000  84.830000 34.080000  84.855000 ;
      RECT 32.585000 162.405000 42.435000 162.555000 ;
      RECT 32.665000  93.325000 40.180000  93.475000 ;
      RECT 32.720000  84.680000 33.930000  84.830000 ;
      RECT 32.735000 162.555000 42.435000 162.705000 ;
      RECT 32.815000  93.175000 40.030000  93.325000 ;
      RECT 32.870000  84.530000 33.780000  84.680000 ;
      RECT 32.885000 162.705000 42.435000 162.855000 ;
      RECT 32.965000  93.025000 39.880000  93.175000 ;
      RECT 33.020000  84.380000 33.630000  84.530000 ;
      RECT 33.020000  84.380000 34.105000  84.855000 ;
      RECT 33.035000 162.855000 42.435000 163.005000 ;
      RECT 33.115000  92.875000 39.730000  93.025000 ;
      RECT 33.185000 163.005000 42.435000 163.155000 ;
      RECT 33.265000  92.725000 39.580000  92.875000 ;
      RECT 33.335000 163.155000 42.435000 163.305000 ;
      RECT 33.415000  92.575000 39.430000  92.725000 ;
      RECT 33.485000 163.305000 42.435000 163.455000 ;
      RECT 33.565000  92.425000 39.280000  92.575000 ;
      RECT 33.635000 163.455000 42.435000 163.605000 ;
      RECT 33.715000  92.275000 39.130000  92.425000 ;
      RECT 33.785000 163.605000 42.435000 163.755000 ;
      RECT 33.865000  92.125000 38.980000  92.275000 ;
      RECT 33.935000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.905000 42.435000 163.970000 ;
      RECT 34.000000 163.970000 39.110000 167.295000 ;
      RECT 34.015000  91.975000 38.830000  92.125000 ;
      RECT 34.150000 163.970000 42.285000 164.120000 ;
      RECT 34.165000  91.825000 38.680000  91.975000 ;
      RECT 34.300000 164.120000 42.135000 164.270000 ;
      RECT 34.315000  91.675000 38.530000  91.825000 ;
      RECT 34.450000 164.270000 41.985000 164.420000 ;
      RECT 34.465000  91.525000 38.380000  91.675000 ;
      RECT 34.600000 164.420000 41.835000 164.570000 ;
      RECT 34.615000  91.375000 38.230000  91.525000 ;
      RECT 34.750000 164.570000 41.685000 164.720000 ;
      RECT 34.765000  91.225000 38.080000  91.375000 ;
      RECT 34.900000 164.720000 41.535000 164.870000 ;
      RECT 34.915000  91.075000 37.930000  91.225000 ;
      RECT 35.050000 164.870000 41.385000 165.020000 ;
      RECT 35.065000  90.925000 37.780000  91.075000 ;
      RECT 35.200000 165.020000 41.235000 165.170000 ;
      RECT 35.215000  90.775000 37.630000  90.925000 ;
      RECT 35.215000  90.775000 40.410000  93.555000 ;
      RECT 35.350000 165.170000 41.085000 165.320000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.825000 39.435000 161.160000 ;
      RECT 35.500000 165.320000 40.935000 165.470000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.650000 165.470000 40.785000 165.620000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.800000 165.620000 40.635000 165.770000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.950000 165.770000 40.485000 165.920000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.100000 165.920000 40.335000 166.070000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.250000 166.070000 40.185000 166.220000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.400000 166.220000 40.035000 166.370000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.550000 166.370000 39.885000 166.520000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.700000 166.520000 39.735000 166.670000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.850000 166.670000 39.585000 166.820000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 166.820000 39.435000 166.970000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 166.970000 39.285000 167.120000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.940000 ;
      RECT 37.280000  69.890000 50.355000  74.340000 ;
      RECT 37.280000  69.890000 50.455000  70.940000 ;
      RECT 37.280000  70.940000 50.455000  74.340000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 167.120000 39.135000 167.270000 ;
      RECT 37.325000 167.270000 39.110000 167.295000 ;
      RECT 37.325000 167.295000 37.545000 168.860000 ;
      RECT 37.325000 167.295000 38.960000 167.445000 ;
      RECT 37.325000 167.445000 38.810000 167.595000 ;
      RECT 37.325000 167.595000 38.660000 167.745000 ;
      RECT 37.325000 167.745000 38.510000 167.895000 ;
      RECT 37.325000 167.895000 38.360000 168.045000 ;
      RECT 37.325000 168.045000 38.210000 168.195000 ;
      RECT 37.325000 168.195000 38.060000 168.345000 ;
      RECT 37.325000 168.345000 37.910000 168.495000 ;
      RECT 37.325000 168.495000 37.760000 168.645000 ;
      RECT 37.325000 168.645000 37.610000 168.795000 ;
      RECT 37.325000 168.795000 37.460000 168.945000 ;
      RECT 37.325000 168.860000 37.545000 189.915000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.190000  95.580000 42.435000  98.585000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.430000  98.585000 42.435000 162.405000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  87.195000 41.210000  87.610000 ;
      RECT 39.810000  84.830000 41.185000  84.855000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.935000  87.195000 41.210000  87.345000 ;
      RECT 39.960000  84.680000 41.035000  84.830000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 40.085000  87.345000 41.210000  87.495000 ;
      RECT 40.110000  84.530000 40.885000  84.680000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.200000  87.495000 41.210000  87.610000 ;
      RECT 40.200000  87.610000 50.245000  96.645000 ;
      RECT 40.260000  84.380000 40.735000  84.530000 ;
      RECT 40.260000  84.380000 41.210000  84.855000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.350000  87.610000 41.210000  87.760000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.500000  87.760000 41.360000  87.910000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.650000  87.910000 41.510000  88.060000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.800000  88.060000 41.660000  88.210000 ;
      RECT 40.950000  88.210000 41.810000  88.360000 ;
      RECT 41.100000  88.360000 41.960000  88.510000 ;
      RECT 41.250000  88.510000 42.110000  88.660000 ;
      RECT 41.400000  88.660000 42.260000  88.810000 ;
      RECT 41.550000  88.810000 42.410000  88.960000 ;
      RECT 41.700000  88.960000 42.560000  89.110000 ;
      RECT 41.850000  89.110000 42.710000  89.260000 ;
      RECT 42.000000  89.260000 42.860000  89.410000 ;
      RECT 42.150000  89.410000 43.010000  89.560000 ;
      RECT 42.300000  89.560000 43.160000  89.710000 ;
      RECT 42.450000  89.710000 43.310000  89.860000 ;
      RECT 42.600000  89.860000 43.460000  90.010000 ;
      RECT 42.750000  90.010000 43.610000  90.160000 ;
      RECT 42.900000  90.160000 43.760000  90.310000 ;
      RECT 43.050000  90.310000 43.910000  90.460000 ;
      RECT 43.200000  90.460000 44.060000  90.610000 ;
      RECT 43.350000  90.610000 44.210000  90.760000 ;
      RECT 43.500000  90.760000 44.360000  90.910000 ;
      RECT 43.650000  90.910000 44.510000  91.060000 ;
      RECT 43.800000  91.060000 44.660000  91.210000 ;
      RECT 43.950000  91.210000 44.810000  91.360000 ;
      RECT 44.100000  91.360000 44.960000  91.510000 ;
      RECT 44.250000  91.510000 45.110000  91.660000 ;
      RECT 44.400000  91.660000 45.260000  91.810000 ;
      RECT 44.550000  91.810000 45.410000  91.960000 ;
      RECT 44.700000  91.960000 45.560000  92.110000 ;
      RECT 44.850000  92.110000 45.710000  92.260000 ;
      RECT 45.000000  92.260000 45.860000  92.410000 ;
      RECT 45.150000  92.410000 46.010000  92.560000 ;
      RECT 45.300000  92.560000 46.160000  92.710000 ;
      RECT 45.450000  92.710000 46.310000  92.860000 ;
      RECT 45.600000  92.860000 46.460000  93.010000 ;
      RECT 45.750000  93.010000 46.610000  93.160000 ;
      RECT 45.900000  93.160000 46.760000  93.310000 ;
      RECT 46.050000  93.310000 46.910000  93.460000 ;
      RECT 46.200000  93.460000 47.060000  93.610000 ;
      RECT 46.350000  93.610000 47.210000  93.760000 ;
      RECT 46.500000  93.760000 47.360000  93.910000 ;
      RECT 46.650000  93.910000 47.510000  94.060000 ;
      RECT 46.800000  94.060000 47.660000  94.210000 ;
      RECT 46.950000  94.210000 47.810000  94.360000 ;
      RECT 46.960000  74.340000 50.455000  76.650000 ;
      RECT 47.100000  94.360000 47.960000  94.510000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.250000  94.510000 48.110000  94.660000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.400000  94.660000 48.260000  94.810000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.550000  94.810000 48.410000  94.960000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.700000  94.960000 48.560000  95.110000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.850000  95.110000 48.710000  95.260000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 48.000000  95.260000 48.860000  95.410000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.150000  95.410000 49.010000  95.560000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.300000  95.560000 49.160000  95.710000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.450000  95.710000 49.310000  95.860000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.600000  95.860000 49.460000  96.010000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.750000  96.010000 49.610000  96.160000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.900000  96.160000 49.760000  96.310000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 49.050000  96.310000 49.910000  96.460000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.200000  96.460000 50.060000  96.610000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.610000 50.210000  96.645000 ;
      RECT 49.235000  96.645000 50.245000  96.795000 ;
      RECT 49.235000  96.645000 53.930000 100.330000 ;
      RECT 49.235000  96.795000 50.395000  96.945000 ;
      RECT 49.235000  96.945000 50.545000  97.095000 ;
      RECT 49.235000  97.095000 50.695000  97.245000 ;
      RECT 49.235000  97.245000 50.845000  97.395000 ;
      RECT 49.235000  97.395000 50.995000  97.545000 ;
      RECT 49.235000  97.545000 51.145000  97.695000 ;
      RECT 49.235000  97.695000 51.295000  97.845000 ;
      RECT 49.235000  97.845000 51.445000  97.995000 ;
      RECT 49.235000  97.995000 51.595000  98.145000 ;
      RECT 49.235000  98.145000 51.745000  98.295000 ;
      RECT 49.235000  98.295000 51.895000  98.445000 ;
      RECT 49.235000  98.445000 52.045000  98.595000 ;
      RECT 49.235000  98.595000 52.195000  98.745000 ;
      RECT 49.235000  98.745000 52.345000  98.895000 ;
      RECT 49.235000  98.895000 52.495000  99.045000 ;
      RECT 49.235000  99.045000 52.645000  99.195000 ;
      RECT 49.235000  99.195000 52.795000  99.345000 ;
      RECT 49.235000  99.345000 52.945000  99.495000 ;
      RECT 49.235000  99.495000 53.095000  99.645000 ;
      RECT 49.235000  99.645000 53.245000  99.795000 ;
      RECT 49.235000  99.795000 53.395000  99.945000 ;
      RECT 49.235000  99.945000 53.545000 100.095000 ;
      RECT 49.235000 100.095000 53.695000 100.245000 ;
      RECT 49.235000 100.245000 53.845000 100.330000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 164.295000 49.470000 168.755000 ;
      RECT 49.235000 164.295000 53.780000 164.445000 ;
      RECT 49.235000 164.445000 53.630000 164.595000 ;
      RECT 49.235000 164.595000 53.480000 164.745000 ;
      RECT 49.235000 164.745000 53.330000 164.895000 ;
      RECT 49.235000 164.895000 53.180000 165.045000 ;
      RECT 49.235000 165.045000 53.030000 165.195000 ;
      RECT 49.235000 165.195000 52.880000 165.345000 ;
      RECT 49.235000 165.345000 52.730000 165.495000 ;
      RECT 49.235000 165.495000 52.580000 165.645000 ;
      RECT 49.235000 165.645000 52.430000 165.795000 ;
      RECT 49.235000 165.795000 52.280000 165.945000 ;
      RECT 49.235000 165.945000 52.130000 166.095000 ;
      RECT 49.235000 166.095000 51.980000 166.245000 ;
      RECT 49.235000 166.245000 51.830000 166.395000 ;
      RECT 49.235000 166.395000 51.680000 166.545000 ;
      RECT 49.235000 166.545000 51.530000 166.695000 ;
      RECT 49.235000 166.695000 51.380000 166.845000 ;
      RECT 49.235000 166.845000 51.230000 166.995000 ;
      RECT 49.235000 166.995000 51.080000 167.145000 ;
      RECT 49.235000 167.145000 50.930000 167.295000 ;
      RECT 49.235000 167.295000 50.780000 167.445000 ;
      RECT 49.235000 167.445000 50.630000 167.595000 ;
      RECT 49.235000 167.595000 50.480000 167.745000 ;
      RECT 49.235000 167.745000 50.330000 167.895000 ;
      RECT 49.235000 167.895000 50.180000 168.045000 ;
      RECT 49.235000 168.045000 50.030000 168.195000 ;
      RECT 49.235000 168.195000 49.880000 168.345000 ;
      RECT 49.235000 168.345000 49.730000 168.495000 ;
      RECT 49.235000 168.495000 49.580000 168.645000 ;
      RECT 49.235000 168.645000 49.430000 168.795000 ;
      RECT 49.235000 168.755000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.280000 168.945000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.650000 50.455000  84.590000 ;
      RECT 49.270000  77.735000 50.355000  84.630000 ;
      RECT 49.270000  84.590000 50.510000  84.645000 ;
      RECT 49.270000  84.630000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.360000  84.640000 ;
      RECT 49.270000  84.640000 50.365000  84.645000 ;
      RECT 49.270000  84.645000 52.660000  86.795000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  84.645000 50.370000  84.795000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  84.795000 50.520000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  84.945000 50.670000  85.095000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  85.095000 50.820000  85.245000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  85.245000 50.970000  85.395000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  85.395000 51.120000  85.545000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  85.545000 51.270000  85.695000 ;
      RECT 50.470000  85.695000 51.420000  85.845000 ;
      RECT 50.620000  85.845000 51.570000  85.995000 ;
      RECT 50.770000  85.995000 51.720000  86.145000 ;
      RECT 50.920000  86.145000 51.870000  86.295000 ;
      RECT 51.070000  86.295000 52.020000  86.445000 ;
      RECT 51.220000  86.445000 52.170000  86.595000 ;
      RECT 51.370000  86.595000 52.320000  86.745000 ;
      RECT 51.420000  86.745000 52.470000  86.795000 ;
      RECT 51.420000  86.795000 52.520000  86.945000 ;
      RECT 51.420000  86.795000 54.075000  88.210000 ;
      RECT 51.420000  86.945000 52.670000  87.095000 ;
      RECT 51.420000  87.095000 52.820000  87.245000 ;
      RECT 51.420000  87.245000 52.970000  87.395000 ;
      RECT 51.420000  87.395000 53.120000  87.545000 ;
      RECT 51.420000  87.545000 53.270000  87.695000 ;
      RECT 51.420000  87.695000 53.420000  87.845000 ;
      RECT 51.420000  87.845000 53.570000  87.995000 ;
      RECT 51.420000  87.995000 53.720000  88.145000 ;
      RECT 51.420000  88.145000 53.870000  88.210000 ;
      RECT 51.420000  88.210000 61.745000  95.880000 ;
      RECT 51.570000  88.210000 53.935000  88.360000 ;
      RECT 51.720000  88.360000 54.085000  88.510000 ;
      RECT 51.870000  88.510000 54.235000  88.660000 ;
      RECT 52.020000  88.660000 54.385000  88.810000 ;
      RECT 52.170000  88.810000 54.535000  88.960000 ;
      RECT 52.320000  88.960000 54.685000  89.110000 ;
      RECT 52.470000  89.110000 54.835000  89.260000 ;
      RECT 52.620000  89.260000 54.985000  89.410000 ;
      RECT 52.770000  89.410000 55.135000  89.560000 ;
      RECT 52.920000  89.560000 55.285000  89.710000 ;
      RECT 53.070000  89.710000 55.435000  89.860000 ;
      RECT 53.220000  89.860000 55.585000  90.010000 ;
      RECT 53.370000  90.010000 55.735000  90.160000 ;
      RECT 53.520000  90.160000 55.885000  90.310000 ;
      RECT 53.670000  90.310000 56.035000  90.460000 ;
      RECT 53.820000  90.460000 56.185000  90.610000 ;
      RECT 53.970000  90.610000 56.335000  90.760000 ;
      RECT 54.120000  90.760000 56.485000  90.910000 ;
      RECT 54.270000  90.910000 56.635000  91.060000 ;
      RECT 54.420000  91.060000 56.785000  91.210000 ;
      RECT 54.570000  91.210000 56.935000  91.360000 ;
      RECT 54.720000  91.360000 57.085000  91.510000 ;
      RECT 54.870000  91.510000 57.235000  91.660000 ;
      RECT 55.020000  91.660000 57.385000  91.810000 ;
      RECT 55.170000  91.810000 57.535000  91.960000 ;
      RECT 55.320000  91.960000 57.685000  92.110000 ;
      RECT 55.470000  92.110000 57.835000  92.260000 ;
      RECT 55.620000  92.260000 57.985000  92.410000 ;
      RECT 55.770000  92.410000 58.135000  92.560000 ;
      RECT 55.920000  92.560000 58.285000  92.710000 ;
      RECT 56.070000  92.710000 58.435000  92.860000 ;
      RECT 56.220000  92.860000 58.585000  93.010000 ;
      RECT 56.370000  93.010000 58.735000  93.160000 ;
      RECT 56.520000  93.160000 58.885000  93.310000 ;
      RECT 56.670000  93.310000 59.035000  93.460000 ;
      RECT 56.820000  93.460000 59.185000  93.610000 ;
      RECT 56.970000  93.610000 59.335000  93.760000 ;
      RECT 57.120000  93.760000 59.485000  93.910000 ;
      RECT 57.270000  93.910000 59.635000  94.060000 ;
      RECT 57.420000  94.060000 59.785000  94.210000 ;
      RECT 57.570000  94.210000 59.935000  94.360000 ;
      RECT 57.720000  94.360000 60.085000  94.510000 ;
      RECT 57.870000  94.510000 60.235000  94.660000 ;
      RECT 58.020000  94.660000 60.385000  94.810000 ;
      RECT 58.170000  94.810000 60.535000  94.960000 ;
      RECT 58.320000  94.960000 60.685000  95.110000 ;
      RECT 58.470000  95.110000 60.835000  95.260000 ;
      RECT 58.620000  95.260000 60.985000  95.410000 ;
      RECT 58.770000  95.410000 61.135000  95.560000 ;
      RECT 58.920000  95.560000 61.285000  95.710000 ;
      RECT 59.070000  95.710000 61.435000  95.860000 ;
      RECT 59.090000  95.880000 61.745000  97.520000 ;
      RECT 59.130000  95.860000 61.585000  95.920000 ;
      RECT 59.280000  95.920000 61.645000  96.070000 ;
      RECT 59.430000  96.070000 61.645000  96.220000 ;
      RECT 59.580000  96.220000 61.645000  96.370000 ;
      RECT 59.730000  96.370000 61.645000  96.520000 ;
      RECT 59.880000  96.520000 61.645000  96.670000 ;
      RECT 60.030000  96.670000 61.645000  96.820000 ;
      RECT 60.180000  96.820000 61.645000  96.970000 ;
      RECT 60.330000  96.970000 61.645000  97.120000 ;
      RECT 60.480000  97.120000 61.645000  97.270000 ;
      RECT 60.630000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.420000 61.645000  97.520000 ;
      RECT 60.730000  97.520000 61.645000 172.635000 ;
      RECT 60.730000  97.520000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 198.000000 ;
    LAYER met4 ;
      RECT  4.820000 102.300000  7.470000 164.545000 ;
      RECT  5.440000 101.650000  5.945000 102.180000 ;
      RECT  5.440000 164.605000  5.945000 165.135000 ;
      RECT  6.070000 101.090000  8.445000 102.160000 ;
      RECT  6.070000 164.625000  8.445000 165.695000 ;
      RECT  6.555000 100.535000  7.060000 101.065000 ;
      RECT  6.555000 165.720000  7.060000 166.250000 ;
      RECT  7.350000  99.950000  9.725000 101.020000 ;
      RECT  7.350000 165.765000  9.725000 166.835000 ;
      RECT  7.535000 102.245000  8.040000 102.775000 ;
      RECT  7.535000 164.010000  8.040000 164.540000 ;
      RECT  7.750000  99.340000  8.255000  99.870000 ;
      RECT  7.750000 166.915000  8.255000 167.445000 ;
      RECT  8.340000  98.810000 10.715000  99.880000 ;
      RECT  8.415000 166.915000 10.700000 167.865000 ;
      RECT  8.650000 101.130000  9.155000 101.660000 ;
      RECT  8.650000 165.125000  9.155000 165.655000 ;
      RECT  8.825000  98.265000  9.330000  98.795000 ;
      RECT  8.825000 167.990000  9.330000 168.520000 ;
      RECT  9.460000  97.645000 11.835000  98.715000 ;
      RECT  9.460000 168.025000 11.835000 169.095000 ;
      RECT  9.845000  99.935000 10.350000 100.465000 ;
      RECT  9.845000 166.320000 10.350000 166.850000 ;
      RECT  9.985000  97.070000 10.490000  97.600000 ;
      RECT  9.985000 169.150000 10.490000 169.680000 ;
      RECT 10.595000  96.475000 11.850000  96.480000 ;
      RECT 10.595000  96.480000 11.835000  97.545000 ;
      RECT 10.610000 169.340000 11.745000 170.260000 ;
      RECT 10.920000  98.860000 11.425000  99.390000 ;
      RECT 10.920000 167.395000 11.425000 167.925000 ;
      RECT 11.095000  95.950000 11.850000  96.475000 ;
      RECT 11.095000 170.260000 11.850000 170.790000 ;
      RECT 11.965000  95.795000 12.835000  98.295000 ;
      RECT 11.965000 168.490000 12.835000 170.990000 ;
      RECT 25.035000  17.815000 25.465000  22.250000 ;
      RECT 25.035000  39.785000 25.365000  41.435000 ;
      RECT 62.225000  95.795000 63.095000  98.295000 ;
      RECT 62.225000 168.490000 63.095000 170.990000 ;
      RECT 63.225000  96.475000 64.465000  97.545000 ;
      RECT 63.225000  97.645000 65.600000  98.715000 ;
      RECT 63.225000 169.160000 64.465000 170.230000 ;
      RECT 63.235000 168.165000 65.495000 169.005000 ;
      RECT 63.635000  98.860000 64.140000  99.390000 ;
      RECT 63.635000 167.395000 64.140000 167.925000 ;
      RECT 64.345000  98.810000 66.720000  99.880000 ;
      RECT 64.345000 166.905000 66.720000 167.975000 ;
      RECT 64.570000  97.070000 65.075000  97.600000 ;
      RECT 64.570000 169.150000 65.075000 169.680000 ;
      RECT 64.710000  99.935000 65.215000 100.465000 ;
      RECT 64.710000 166.320000 65.215000 166.850000 ;
      RECT 65.335000  99.950000 67.710000 101.020000 ;
      RECT 65.335000 165.765000 67.710000 166.835000 ;
      RECT 65.730000  98.265000 66.235000  98.795000 ;
      RECT 65.730000 167.990000 66.235000 168.520000 ;
      RECT 65.905000 101.130000 66.410000 101.660000 ;
      RECT 65.905000 165.125000 66.410000 165.655000 ;
      RECT 66.615000 101.090000 68.990000 102.160000 ;
      RECT 66.615000 164.625000 68.990000 165.695000 ;
      RECT 66.805000  99.340000 67.310000  99.870000 ;
      RECT 66.805000 166.915000 67.310000 167.445000 ;
      RECT 67.020000 102.245000 70.110000 102.775000 ;
      RECT 67.020000 164.010000 70.165000 164.350000 ;
      RECT 67.020000 164.350000 67.525000 164.540000 ;
      RECT 67.515000 103.000000 70.165000 164.010000 ;
      RECT 68.000000 100.535000 68.505000 101.065000 ;
      RECT 68.000000 165.720000 68.505000 166.250000 ;
      RECT 69.115000 101.650000 69.620000 102.180000 ;
      RECT 69.115000 164.605000 69.620000 165.135000 ;
  END
END sky130_fd_io__top_ground_lvc_wpad
MACRO avsdpll_1v8
  CLASS CORE ;
  FOREIGN avsdpll_1v8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.180 BY 13.710 ;
  SITE unithddb1 ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 10.030 10.380 10.250 10.970 ;
        RECT 11.590 10.380 11.760 11.170 ;
        RECT 14.250 10.380 14.420 11.160 ;
        RECT 16.980 10.380 17.150 11.170 ;
        RECT 18.090 10.380 18.260 11.170 ;
        RECT 9.320 10.210 18.670 10.380 ;
        RECT 0.990 9.740 10.340 9.910 ;
        RECT 11.400 9.740 20.750 9.910 ;
        RECT 1.700 9.150 1.920 9.740 ;
        RECT 3.260 8.950 3.430 9.740 ;
        RECT 5.920 8.960 6.090 9.740 ;
        RECT 8.650 8.950 8.820 9.740 ;
        RECT 9.760 8.950 9.930 9.740 ;
        RECT 12.110 9.150 12.330 9.740 ;
        RECT 13.670 8.950 13.840 9.740 ;
        RECT 16.330 8.960 16.500 9.740 ;
        RECT 19.060 8.950 19.230 9.740 ;
        RECT 20.170 8.950 20.340 9.740 ;
      LAYER mcon ;
        RECT 9.670 10.210 9.840 10.380 ;
        RECT 10.510 10.210 10.680 10.380 ;
        RECT 11.350 10.210 11.520 10.380 ;
        RECT 12.530 10.210 12.700 10.380 ;
        RECT 13.370 10.210 13.540 10.380 ;
        RECT 14.430 10.210 14.600 10.380 ;
        RECT 15.350 10.210 15.520 10.380 ;
        RECT 16.700 10.210 16.870 10.380 ;
        RECT 17.500 10.210 17.670 10.380 ;
        RECT 18.340 10.210 18.510 10.380 ;
        RECT 1.340 9.740 1.510 9.910 ;
        RECT 2.180 9.740 2.350 9.910 ;
        RECT 3.020 9.740 3.190 9.910 ;
        RECT 4.200 9.740 4.370 9.910 ;
        RECT 5.040 9.740 5.210 9.910 ;
        RECT 6.100 9.740 6.270 9.910 ;
        RECT 7.020 9.740 7.190 9.910 ;
        RECT 8.370 9.740 8.540 9.910 ;
        RECT 9.170 9.740 9.340 9.910 ;
        RECT 10.010 9.740 10.180 9.910 ;
        RECT 11.750 9.740 11.920 9.910 ;
        RECT 12.590 9.740 12.760 9.910 ;
        RECT 13.430 9.740 13.600 9.910 ;
        RECT 14.610 9.740 14.780 9.910 ;
        RECT 15.450 9.740 15.620 9.910 ;
        RECT 16.510 9.740 16.680 9.910 ;
        RECT 17.430 9.740 17.600 9.910 ;
        RECT 18.780 9.740 18.950 9.910 ;
        RECT 19.580 9.740 19.750 9.910 ;
        RECT 20.420 9.740 20.590 9.910 ;
      LAYER met1 ;
        RECT 9.320 10.060 18.670 10.540 ;
        RECT 0.000 9.750 0.310 9.890 ;
        RECT 0.590 9.750 10.340 10.060 ;
        RECT 0.000 9.580 10.340 9.750 ;
        RECT 11.400 9.580 20.750 10.060 ;
        RECT 0.000 9.120 0.900 9.580 ;
        RECT 0.000 8.980 0.310 9.120 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 21.140 9.820 34.410 10.910 ;
        RECT 2.480 8.510 3.550 8.580 ;
        RECT 2.480 8.460 3.670 8.510 ;
        RECT 1.020 8.220 3.670 8.460 ;
        RECT 5.240 8.220 6.380 8.570 ;
        RECT 1.020 8.210 6.380 8.220 ;
        RECT 7.970 8.560 11.450 8.570 ;
        RECT 12.890 8.560 13.960 8.580 ;
        RECT 21.140 8.570 26.420 9.820 ;
        RECT 29.420 9.810 34.410 9.820 ;
        RECT 30.710 8.760 34.410 9.810 ;
        RECT 31.070 8.750 34.410 8.760 ;
        RECT 7.970 8.510 13.960 8.560 ;
        RECT 7.970 8.220 14.080 8.510 ;
        RECT 15.650 8.220 16.790 8.570 ;
        RECT 7.970 8.210 16.790 8.220 ;
        RECT 18.380 8.210 26.420 8.570 ;
        RECT 1.020 6.860 26.420 8.210 ;
        RECT 1.900 6.720 26.420 6.860 ;
        RECT 1.900 5.810 29.330 6.720 ;
        RECT 2.380 5.250 29.330 5.810 ;
        RECT 6.060 5.130 29.330 5.250 ;
        RECT 6.060 5.060 16.830 5.130 ;
        RECT 8.790 4.820 16.830 5.060 ;
        RECT 10.630 4.690 16.830 4.820 ;
        RECT 10.970 4.540 16.830 4.690 ;
        RECT 11.080 4.490 16.830 4.540 ;
        RECT 20.250 4.390 29.330 5.130 ;
        RECT 20.250 4.350 28.090 4.390 ;
        RECT 20.250 4.340 21.550 4.350 ;
        RECT 20.250 4.040 21.180 4.340 ;
      LAYER li1 ;
        RECT 33.940 8.930 34.110 10.240 ;
        RECT 1.700 7.230 1.930 7.840 ;
        RECT 3.260 7.230 3.430 8.330 ;
        RECT 5.920 7.230 6.090 8.340 ;
        RECT 8.650 7.230 8.820 8.330 ;
        RECT 9.760 7.230 9.930 8.330 ;
        RECT 12.110 7.230 12.340 7.840 ;
        RECT 13.670 7.230 13.840 8.330 ;
        RECT 16.330 7.230 16.500 8.340 ;
        RECT 19.060 7.230 19.230 8.330 ;
        RECT 20.170 7.230 20.340 8.330 ;
        RECT 1.020 7.040 10.340 7.230 ;
        RECT 11.430 7.040 20.750 7.230 ;
        RECT 23.360 7.210 23.700 7.990 ;
        RECT 21.140 7.040 30.160 7.210 ;
        RECT 8.470 6.680 29.330 6.700 ;
        RECT 1.010 6.530 29.330 6.680 ;
        RECT 1.010 6.510 8.680 6.530 ;
        RECT 2.660 6.180 3.080 6.510 ;
        RECT 2.520 5.970 3.230 6.180 ;
        RECT 6.780 5.540 7.010 6.510 ;
        RECT 11.150 6.310 29.150 6.530 ;
        RECT 22.050 4.660 28.820 4.870 ;
      LAYER mcon ;
        RECT 1.610 7.040 1.800 7.230 ;
        RECT 2.470 7.040 2.660 7.230 ;
        RECT 3.330 7.040 3.520 7.230 ;
        RECT 4.530 7.040 4.720 7.230 ;
        RECT 5.610 7.040 5.800 7.230 ;
        RECT 6.550 7.040 6.740 7.230 ;
        RECT 7.330 7.040 7.520 7.230 ;
        RECT 8.780 7.040 8.970 7.230 ;
        RECT 9.600 7.040 9.790 7.230 ;
        RECT 12.020 7.040 12.210 7.230 ;
        RECT 12.880 7.040 13.070 7.230 ;
        RECT 13.740 7.040 13.930 7.230 ;
        RECT 14.940 7.040 15.130 7.230 ;
        RECT 16.020 7.040 16.210 7.230 ;
        RECT 16.960 7.040 17.150 7.230 ;
        RECT 17.740 7.040 17.930 7.230 ;
        RECT 19.190 7.040 19.380 7.230 ;
        RECT 20.010 7.040 20.200 7.230 ;
        RECT 21.370 7.040 21.540 7.210 ;
        RECT 21.710 7.040 21.880 7.210 ;
        RECT 22.050 7.040 22.220 7.210 ;
        RECT 22.390 7.040 22.560 7.210 ;
        RECT 22.730 7.040 22.900 7.210 ;
        RECT 23.070 7.040 23.240 7.210 ;
        RECT 23.410 7.040 23.580 7.210 ;
        RECT 23.750 7.040 23.920 7.210 ;
        RECT 24.090 7.040 24.260 7.210 ;
        RECT 24.430 7.040 24.600 7.210 ;
        RECT 24.770 7.040 24.940 7.210 ;
        RECT 25.110 7.040 25.280 7.210 ;
        RECT 25.450 7.040 25.620 7.210 ;
        RECT 25.790 7.040 25.960 7.210 ;
        RECT 26.130 7.040 26.300 7.210 ;
        RECT 26.470 7.040 26.640 7.210 ;
        RECT 26.810 7.040 26.980 7.210 ;
        RECT 27.150 7.040 27.320 7.210 ;
        RECT 27.490 7.040 27.660 7.210 ;
        RECT 27.830 7.040 28.000 7.210 ;
        RECT 28.170 7.040 28.340 7.210 ;
        RECT 28.510 7.040 28.680 7.210 ;
        RECT 28.850 7.040 29.020 7.210 ;
        RECT 29.190 7.040 29.360 7.210 ;
        RECT 29.530 7.040 29.700 7.210 ;
        RECT 29.870 7.040 30.040 7.210 ;
        RECT 1.810 6.510 1.980 6.680 ;
        RECT 2.150 6.510 2.320 6.680 ;
        RECT 2.490 6.510 2.660 6.680 ;
        RECT 2.830 6.510 3.000 6.680 ;
        RECT 3.170 6.510 3.340 6.680 ;
        RECT 3.510 6.510 3.680 6.680 ;
        RECT 3.850 6.510 4.020 6.680 ;
        RECT 4.190 6.510 4.360 6.680 ;
        RECT 4.530 6.510 4.700 6.680 ;
        RECT 4.870 6.510 5.040 6.680 ;
        RECT 5.210 6.510 5.380 6.680 ;
        RECT 5.550 6.510 5.720 6.680 ;
        RECT 5.890 6.510 6.060 6.680 ;
        RECT 6.230 6.510 6.400 6.680 ;
        RECT 6.570 6.510 6.740 6.680 ;
        RECT 6.910 6.510 7.080 6.680 ;
        RECT 7.250 6.510 7.420 6.680 ;
        RECT 7.590 6.510 7.760 6.680 ;
        RECT 8.880 6.530 9.050 6.700 ;
        RECT 9.220 6.530 9.390 6.700 ;
        RECT 9.560 6.530 9.730 6.700 ;
        RECT 9.900 6.530 10.070 6.700 ;
        RECT 10.240 6.530 10.410 6.700 ;
        RECT 10.580 6.530 10.750 6.700 ;
        RECT 10.920 6.530 11.090 6.700 ;
        RECT 11.260 6.530 11.430 6.700 ;
        RECT 11.600 6.530 11.770 6.700 ;
        RECT 11.940 6.530 12.110 6.700 ;
        RECT 12.280 6.530 12.450 6.700 ;
        RECT 12.620 6.530 12.790 6.700 ;
        RECT 12.960 6.530 13.130 6.700 ;
        RECT 13.300 6.530 13.470 6.700 ;
        RECT 13.640 6.530 13.810 6.700 ;
        RECT 13.980 6.530 14.150 6.700 ;
        RECT 14.320 6.530 14.490 6.700 ;
        RECT 14.660 6.530 14.830 6.700 ;
        RECT 15.000 6.530 15.170 6.700 ;
        RECT 15.340 6.530 15.510 6.700 ;
        RECT 15.680 6.530 15.850 6.700 ;
        RECT 16.020 6.530 16.190 6.700 ;
        RECT 16.360 6.530 16.530 6.700 ;
        RECT 16.700 6.530 16.870 6.700 ;
        RECT 17.040 6.530 17.210 6.700 ;
        RECT 17.380 6.530 17.550 6.700 ;
        RECT 17.720 6.530 17.890 6.700 ;
        RECT 18.060 6.530 18.230 6.700 ;
        RECT 18.400 6.530 18.570 6.700 ;
        RECT 18.740 6.530 18.910 6.700 ;
        RECT 19.080 6.530 19.250 6.700 ;
        RECT 19.420 6.530 19.590 6.700 ;
        RECT 19.760 6.530 19.930 6.700 ;
        RECT 20.100 6.530 20.270 6.700 ;
        RECT 20.440 6.530 20.610 6.700 ;
        RECT 20.780 6.530 20.950 6.700 ;
        RECT 21.120 6.530 21.290 6.700 ;
        RECT 21.460 6.530 21.630 6.700 ;
        RECT 21.800 6.530 21.970 6.700 ;
        RECT 22.140 6.530 22.310 6.700 ;
        RECT 22.480 6.530 22.650 6.700 ;
        RECT 22.820 6.530 22.990 6.700 ;
        RECT 23.160 6.530 23.330 6.700 ;
        RECT 23.500 6.530 23.670 6.700 ;
        RECT 23.840 6.530 24.010 6.700 ;
        RECT 24.180 6.530 24.350 6.700 ;
        RECT 24.520 6.530 24.690 6.700 ;
        RECT 24.860 6.530 25.030 6.700 ;
        RECT 25.200 6.530 25.370 6.700 ;
        RECT 25.540 6.530 25.710 6.700 ;
        RECT 25.880 6.530 26.050 6.700 ;
        RECT 26.220 6.530 26.390 6.700 ;
        RECT 26.560 6.530 26.730 6.700 ;
        RECT 26.900 6.530 27.070 6.700 ;
        RECT 27.240 6.530 27.410 6.700 ;
        RECT 27.580 6.530 27.750 6.700 ;
        RECT 27.920 6.530 28.090 6.700 ;
        RECT 28.260 6.530 28.430 6.700 ;
        RECT 28.600 6.530 28.770 6.700 ;
        RECT 28.940 6.530 29.110 6.700 ;
        RECT 27.490 4.680 27.660 4.850 ;
        RECT 27.920 4.680 28.090 4.850 ;
      LAYER met1 ;
        RECT 0.000 7.340 0.310 7.410 ;
        RECT 0.000 6.860 10.340 7.340 ;
        RECT 11.430 7.030 20.750 7.340 ;
        RECT 21.140 7.030 30.160 7.340 ;
        RECT 11.430 6.860 30.160 7.030 ;
        RECT 0.000 6.670 29.330 6.860 ;
        RECT 0.000 6.500 0.320 6.670 ;
        RECT 1.010 6.380 29.330 6.670 ;
        RECT 27.430 4.920 28.130 6.380 ;
        RECT 27.430 4.620 28.150 4.920 ;
    END
  END VDD
  PIN ENb_CP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.024000 ;
    PORT
      LAYER li1 ;
        RECT 31.440 9.940 31.770 10.110 ;
        RECT 32.570 7.660 32.900 7.870 ;
        RECT 33.440 7.680 33.770 7.850 ;
        RECT 8.740 5.520 9.100 5.610 ;
        RECT 8.740 5.510 9.610 5.520 ;
        RECT 8.740 5.270 9.630 5.510 ;
        RECT 8.740 5.260 9.610 5.270 ;
        RECT 8.740 5.250 9.100 5.260 ;
      LAYER mcon ;
        RECT 31.520 9.940 31.690 10.110 ;
        RECT 32.650 7.680 32.820 7.850 ;
        RECT 33.520 7.680 33.690 7.850 ;
        RECT 8.770 5.340 8.940 5.510 ;
      LAYER met1 ;
        RECT 31.450 9.860 31.770 10.180 ;
        RECT 32.580 7.910 32.900 7.920 ;
        RECT 32.580 7.610 34.530 7.910 ;
        RECT 32.580 7.600 32.900 7.610 ;
        RECT 8.690 5.250 9.040 5.610 ;
      LAYER via ;
        RECT 31.480 9.890 31.740 10.150 ;
        RECT 32.610 7.630 32.870 7.890 ;
        RECT 8.720 5.280 9.010 5.570 ;
      LAYER met2 ;
        RECT 31.450 10.140 31.770 10.180 ;
        RECT 31.450 9.890 32.300 10.140 ;
        RECT 31.450 9.860 31.770 9.890 ;
        RECT 32.050 8.940 32.300 9.890 ;
        RECT 31.820 8.700 32.300 8.940 ;
        RECT 32.050 7.910 32.300 8.700 ;
        RECT 32.580 7.910 32.900 7.920 ;
        RECT 32.050 7.610 32.900 7.910 ;
        RECT 32.580 7.600 32.900 7.610 ;
        RECT 32.590 7.450 32.870 7.600 ;
        RECT 28.720 7.150 32.890 7.450 ;
        RECT 28.720 7.030 29.250 7.150 ;
        RECT 3.020 6.710 29.250 7.030 ;
        RECT 0.000 5.840 0.280 6.060 ;
        RECT 3.020 5.840 3.350 6.710 ;
        RECT 0.000 5.520 3.350 5.840 ;
        RECT 0.000 5.290 0.280 5.520 ;
        RECT 8.690 5.250 9.040 6.710 ;
    END
  END ENb_CP
  PIN CLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.351000 ;
    ANTENNADIFFAREA 0.469800 ;
    PORT
      LAYER li1 ;
        RECT 12.010 12.220 12.180 12.560 ;
        RECT 20.300 11.770 20.680 11.850 ;
        RECT 20.300 11.540 20.690 11.770 ;
        RECT 18.010 11.370 20.760 11.540 ;
        RECT 20.210 11.180 20.760 11.370 ;
        RECT 21.380 11.180 21.550 11.930 ;
        RECT 15.970 10.800 16.300 10.980 ;
        RECT 20.210 10.950 21.550 11.180 ;
        RECT 20.210 10.940 21.210 10.950 ;
        RECT 21.380 9.650 21.550 10.950 ;
      LAYER mcon ;
        RECT 12.010 12.300 12.180 12.470 ;
        RECT 20.420 11.570 20.590 11.740 ;
        RECT 18.090 11.370 18.260 11.540 ;
        RECT 16.050 10.810 16.220 10.980 ;
      LAYER met1 ;
        RECT 11.950 12.550 12.230 12.560 ;
        RECT 11.950 12.130 12.240 12.550 ;
        RECT 17.100 12.240 18.320 12.560 ;
        RECT 17.100 12.130 17.350 12.240 ;
        RECT 11.950 11.880 17.350 12.130 ;
        RECT 18.030 11.330 18.320 12.240 ;
        RECT 20.340 11.500 20.660 11.820 ;
        RECT 18.030 11.040 18.310 11.330 ;
        RECT 15.960 10.750 18.310 11.040 ;
      LAYER via ;
        RECT 20.370 11.530 20.630 11.790 ;
      LAYER met2 ;
        RECT 20.310 11.470 20.690 11.850 ;
        RECT 29.190 1.570 29.920 1.920 ;
        RECT 29.190 1.140 30.340 1.570 ;
        RECT 29.810 0.280 30.340 1.140 ;
        RECT 29.690 0.000 30.460 0.280 ;
      LAYER via2 ;
        RECT 20.360 11.520 20.640 11.800 ;
        RECT 29.250 1.200 29.850 1.860 ;
      LAYER met3 ;
        RECT 20.310 11.570 20.930 11.850 ;
        RECT 20.310 11.470 20.940 11.570 ;
        RECT 20.550 5.550 20.940 11.470 ;
        RECT 20.550 5.540 22.930 5.550 ;
        RECT 20.550 5.140 23.300 5.540 ;
        RECT 22.680 4.370 23.300 5.140 ;
        RECT 22.680 2.300 23.310 4.370 ;
        RECT 22.690 1.610 23.310 2.300 ;
        RECT 29.190 1.610 29.920 1.920 ;
        RECT 22.690 1.130 29.920 1.610 ;
    END
  END CLK
  PIN ENb_VCO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 23.350 8.360 23.700 8.700 ;
      LAYER mcon ;
        RECT 23.440 8.460 23.610 8.630 ;
      LAYER met1 ;
        RECT 21.260 8.380 23.670 8.690 ;
        RECT 21.360 8.100 21.800 8.380 ;
      LAYER via ;
        RECT 21.410 8.150 21.670 8.410 ;
      LAYER met2 ;
        RECT 2.890 10.200 19.740 10.210 ;
        RECT 2.890 9.920 21.720 10.200 ;
        RECT 0.000 8.280 0.280 8.540 ;
        RECT 2.890 8.280 3.200 9.920 ;
        RECT 18.040 9.910 21.720 9.920 ;
        RECT 21.380 8.460 21.720 9.910 ;
        RECT 0.000 7.990 3.200 8.280 ;
        RECT 21.360 8.090 21.720 8.460 ;
        RECT 0.000 7.770 0.280 7.990 ;
    END
  END ENb_VCO
  PIN GND#2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 5.350 3.750 6.020 4.560 ;
        RECT 6.790 3.820 7.010 4.340 ;
        RECT 6.570 3.750 7.240 3.820 ;
        RECT 5.350 3.730 8.850 3.750 ;
        RECT 9.970 3.730 15.040 4.010 ;
        RECT 17.270 3.730 17.690 3.980 ;
        RECT 5.350 3.580 19.080 3.730 ;
        RECT 8.680 3.560 19.080 3.580 ;
        RECT 19.810 3.560 29.330 3.730 ;
        RECT 1.790 3.220 2.000 3.240 ;
        RECT 1.710 3.050 2.070 3.220 ;
        RECT 1.790 2.970 2.000 3.050 ;
        RECT 9.600 2.500 9.790 3.560 ;
        RECT 10.840 2.500 11.030 3.560 ;
        RECT 12.680 3.190 17.920 3.560 ;
        RECT 20.750 3.280 28.240 3.560 ;
        RECT 12.680 3.180 18.090 3.190 ;
        RECT 12.550 3.010 18.090 3.180 ;
        RECT 13.290 3.000 18.090 3.010 ;
        RECT 2.740 1.380 2.920 1.740 ;
        RECT 7.040 1.160 7.260 1.490 ;
      LAYER mcon ;
        RECT 5.950 3.580 6.120 3.750 ;
        RECT 6.290 3.580 6.460 3.750 ;
        RECT 6.630 3.580 6.800 3.750 ;
        RECT 6.970 3.580 7.140 3.750 ;
        RECT 7.310 3.580 7.480 3.750 ;
        RECT 7.650 3.580 7.820 3.750 ;
        RECT 8.880 3.560 9.050 3.730 ;
        RECT 9.220 3.560 9.390 3.730 ;
        RECT 9.560 3.560 9.730 3.730 ;
        RECT 9.900 3.560 10.070 3.730 ;
        RECT 10.240 3.560 10.410 3.730 ;
        RECT 10.580 3.560 10.750 3.730 ;
        RECT 10.920 3.560 11.090 3.730 ;
        RECT 11.260 3.560 11.430 3.730 ;
        RECT 11.600 3.560 11.770 3.730 ;
        RECT 11.940 3.560 12.110 3.730 ;
        RECT 12.280 3.560 12.450 3.730 ;
        RECT 12.620 3.560 12.790 3.730 ;
        RECT 12.960 3.560 13.130 3.730 ;
        RECT 13.300 3.560 13.470 3.730 ;
        RECT 13.640 3.560 13.810 3.730 ;
        RECT 13.980 3.560 14.150 3.730 ;
        RECT 14.320 3.560 14.490 3.730 ;
        RECT 14.660 3.560 14.830 3.730 ;
        RECT 15.000 3.560 15.170 3.730 ;
        RECT 15.340 3.560 15.510 3.730 ;
        RECT 15.680 3.560 15.850 3.730 ;
        RECT 16.020 3.560 16.190 3.730 ;
        RECT 16.360 3.560 16.530 3.730 ;
        RECT 16.700 3.560 16.870 3.730 ;
        RECT 17.040 3.560 17.210 3.730 ;
        RECT 17.380 3.560 17.550 3.730 ;
        RECT 17.720 3.560 17.890 3.730 ;
        RECT 18.060 3.560 18.230 3.730 ;
        RECT 18.400 3.560 18.570 3.730 ;
        RECT 18.740 3.560 18.910 3.730 ;
        RECT 20.100 3.560 20.270 3.730 ;
        RECT 20.440 3.560 20.610 3.730 ;
        RECT 20.780 3.560 20.950 3.730 ;
        RECT 21.120 3.560 21.290 3.730 ;
        RECT 21.460 3.560 21.630 3.730 ;
        RECT 21.800 3.560 21.970 3.730 ;
        RECT 22.140 3.560 22.310 3.730 ;
        RECT 22.480 3.560 22.650 3.730 ;
        RECT 22.820 3.560 22.990 3.730 ;
        RECT 23.160 3.560 23.330 3.730 ;
        RECT 23.500 3.560 23.670 3.730 ;
        RECT 23.840 3.560 24.010 3.730 ;
        RECT 24.180 3.560 24.350 3.730 ;
        RECT 24.520 3.560 24.690 3.730 ;
        RECT 24.860 3.560 25.030 3.730 ;
        RECT 25.200 3.560 25.370 3.730 ;
        RECT 25.540 3.560 25.710 3.730 ;
        RECT 25.880 3.560 26.050 3.730 ;
        RECT 26.220 3.560 26.390 3.730 ;
        RECT 26.560 3.560 26.730 3.730 ;
        RECT 26.900 3.560 27.070 3.730 ;
        RECT 27.240 3.560 27.410 3.730 ;
        RECT 27.580 3.560 27.750 3.730 ;
        RECT 27.920 3.560 28.090 3.730 ;
        RECT 28.260 3.560 28.430 3.730 ;
        RECT 28.600 3.560 28.770 3.730 ;
        RECT 1.810 3.050 1.980 3.220 ;
        RECT 2.750 1.470 2.920 1.640 ;
        RECT 7.080 1.240 7.250 1.410 ;
      LAYER met1 ;
        RECT 0.000 4.660 0.310 4.830 ;
        RECT 0.000 4.230 1.020 4.660 ;
        RECT 0.000 3.920 0.310 4.230 ;
        RECT 0.650 3.900 1.020 4.230 ;
        RECT 0.650 3.420 29.330 3.900 ;
        RECT 1.750 2.990 2.050 3.420 ;
        RECT 3.290 1.700 3.530 3.420 ;
        RECT 2.690 1.410 3.530 1.700 ;
        RECT 6.610 1.470 6.880 3.420 ;
        RECT 6.610 1.180 7.280 1.470 ;
    END
  END GND#2
  PIN VDD#2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.780 3.530 8.930 3.540 ;
        RECT 5.440 3.410 8.930 3.530 ;
        RECT 4.980 2.140 8.930 3.410 ;
        RECT 4.980 2.030 11.820 2.140 ;
        RECT 4.980 0.770 6.150 2.030 ;
        RECT 8.090 1.630 11.820 2.030 ;
        RECT 8.090 0.780 12.570 1.630 ;
        RECT 19.220 1.610 20.060 2.060 ;
        RECT 19.220 0.770 21.080 1.610 ;
      LAYER li1 ;
        RECT 7.030 3.000 7.260 3.390 ;
        RECT 8.050 3.120 8.460 3.290 ;
        RECT 7.030 2.710 7.340 3.000 ;
        RECT 8.110 2.830 8.410 3.120 ;
        RECT 7.030 2.690 7.260 2.710 ;
        RECT 8.050 2.660 8.460 2.830 ;
        RECT 8.110 2.390 8.410 2.660 ;
        RECT 8.050 2.220 8.460 2.390 ;
        RECT 5.700 0.770 5.910 1.880 ;
        RECT 11.890 0.780 12.570 1.190 ;
        RECT 20.270 0.780 21.080 1.280 ;
        RECT 8.470 0.770 29.340 0.780 ;
        RECT 1.010 0.610 29.340 0.770 ;
        RECT 1.010 0.600 8.680 0.610 ;
      LAYER mcon ;
        RECT 7.170 2.770 7.340 2.940 ;
        RECT 8.150 2.640 8.360 2.850 ;
        RECT 1.810 0.600 1.980 0.770 ;
        RECT 2.150 0.600 2.320 0.770 ;
        RECT 2.490 0.600 2.660 0.770 ;
        RECT 2.830 0.600 3.000 0.770 ;
        RECT 3.170 0.600 3.340 0.770 ;
        RECT 3.510 0.600 3.680 0.770 ;
        RECT 3.850 0.600 4.020 0.770 ;
        RECT 4.190 0.600 4.360 0.770 ;
        RECT 4.530 0.600 4.700 0.770 ;
        RECT 4.870 0.600 5.040 0.770 ;
        RECT 5.210 0.600 5.380 0.770 ;
        RECT 5.550 0.600 5.720 0.770 ;
        RECT 5.890 0.600 6.060 0.770 ;
        RECT 6.230 0.600 6.400 0.770 ;
        RECT 6.570 0.600 6.740 0.770 ;
        RECT 6.910 0.600 7.080 0.770 ;
        RECT 7.250 0.600 7.420 0.770 ;
        RECT 7.590 0.600 7.760 0.770 ;
        RECT 8.880 0.610 9.050 0.780 ;
        RECT 9.220 0.610 9.390 0.780 ;
        RECT 9.560 0.610 9.730 0.780 ;
        RECT 9.900 0.610 10.070 0.780 ;
        RECT 10.240 0.610 10.410 0.780 ;
        RECT 10.580 0.610 10.750 0.780 ;
        RECT 10.920 0.610 11.090 0.780 ;
        RECT 11.260 0.610 11.430 0.780 ;
        RECT 11.600 0.610 11.770 0.780 ;
        RECT 11.940 0.610 12.110 0.780 ;
        RECT 12.280 0.610 12.450 0.780 ;
        RECT 12.620 0.610 12.790 0.780 ;
        RECT 12.960 0.610 13.130 0.780 ;
        RECT 13.300 0.610 13.470 0.780 ;
        RECT 13.640 0.610 13.810 0.780 ;
        RECT 13.980 0.610 14.150 0.780 ;
        RECT 14.320 0.610 14.490 0.780 ;
        RECT 14.660 0.610 14.830 0.780 ;
        RECT 15.000 0.610 15.170 0.780 ;
        RECT 15.340 0.610 15.510 0.780 ;
        RECT 15.680 0.610 15.850 0.780 ;
        RECT 16.020 0.610 16.190 0.780 ;
        RECT 16.360 0.610 16.530 0.780 ;
        RECT 16.700 0.610 16.870 0.780 ;
        RECT 17.040 0.610 17.210 0.780 ;
        RECT 17.380 0.610 17.550 0.780 ;
        RECT 17.720 0.610 17.890 0.780 ;
        RECT 18.060 0.610 18.230 0.780 ;
        RECT 18.400 0.610 18.570 0.780 ;
        RECT 18.740 0.610 18.910 0.780 ;
        RECT 19.080 0.610 19.250 0.780 ;
        RECT 19.420 0.610 19.590 0.780 ;
        RECT 19.760 0.610 19.930 0.780 ;
        RECT 20.100 0.610 20.270 0.780 ;
        RECT 20.440 0.610 20.610 0.780 ;
        RECT 20.780 0.610 20.950 0.780 ;
        RECT 21.120 0.610 21.290 0.780 ;
        RECT 21.460 0.610 21.630 0.780 ;
        RECT 21.800 0.610 21.970 0.780 ;
        RECT 22.140 0.610 22.310 0.780 ;
        RECT 22.480 0.610 22.650 0.780 ;
        RECT 22.820 0.610 22.990 0.780 ;
        RECT 23.160 0.610 23.330 0.780 ;
        RECT 23.500 0.610 23.670 0.780 ;
        RECT 23.840 0.610 24.010 0.780 ;
        RECT 24.180 0.610 24.350 0.780 ;
        RECT 24.520 0.610 24.690 0.780 ;
        RECT 24.860 0.610 25.030 0.780 ;
        RECT 25.200 0.610 25.370 0.780 ;
        RECT 25.540 0.610 25.710 0.780 ;
        RECT 25.880 0.610 26.050 0.780 ;
        RECT 26.220 0.610 26.390 0.780 ;
        RECT 26.560 0.610 26.730 0.780 ;
        RECT 26.900 0.610 27.070 0.780 ;
        RECT 27.240 0.610 27.410 0.780 ;
        RECT 27.580 0.610 27.750 0.780 ;
        RECT 27.920 0.610 28.090 0.780 ;
        RECT 28.260 0.610 28.430 0.780 ;
        RECT 28.600 0.610 28.770 0.780 ;
      LAYER met1 ;
        RECT 7.110 2.710 8.420 3.000 ;
        RECT 7.570 2.530 8.420 2.710 ;
        RECT 7.570 0.940 7.870 2.530 ;
        RECT 1.010 0.460 29.340 0.940 ;
        RECT 28.530 0.310 29.040 0.460 ;
        RECT 28.320 0.000 29.230 0.310 ;
    END
  END VDD#2
  PIN VCO_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.313200 ;
    PORT
      LAYER li1 ;
        RECT 32.880 8.800 33.050 9.650 ;
        RECT 32.880 8.530 33.200 8.800 ;
        RECT 32.880 8.050 33.050 8.530 ;
      LAYER mcon ;
        RECT 33.010 8.570 33.180 8.740 ;
      LAYER met1 ;
        RECT 35.210 8.810 35.530 8.820 ;
        RECT 32.950 8.510 35.530 8.810 ;
        RECT 35.210 8.500 35.530 8.510 ;
      LAYER via ;
        RECT 35.240 8.530 35.500 8.790 ;
      LAYER met2 ;
        RECT 35.900 8.820 36.180 9.040 ;
        RECT 35.210 8.500 36.180 8.820 ;
        RECT 35.900 8.270 36.180 8.500 ;
    END
  END VCO_IN
  PIN VDD#3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 9.350 11.910 18.670 13.260 ;
        RECT 9.350 11.900 14.710 11.910 ;
        RECT 9.350 11.660 12.000 11.900 ;
        RECT 10.810 11.610 12.000 11.660 ;
        RECT 10.810 11.540 11.880 11.610 ;
        RECT 13.570 11.550 14.710 11.900 ;
        RECT 16.300 11.550 18.670 11.910 ;
      LAYER li1 ;
        RECT 9.350 12.890 18.670 13.080 ;
        RECT 20.180 12.940 30.160 13.110 ;
        RECT 10.030 12.280 10.260 12.890 ;
        RECT 11.590 11.790 11.760 12.890 ;
        RECT 14.250 11.780 14.420 12.890 ;
        RECT 16.980 11.790 17.150 12.890 ;
        RECT 18.090 11.790 18.260 12.890 ;
      LAYER mcon ;
        RECT 9.940 12.890 10.130 13.080 ;
        RECT 10.800 12.890 10.990 13.080 ;
        RECT 11.660 12.890 11.850 13.080 ;
        RECT 12.860 12.890 13.050 13.080 ;
        RECT 13.940 12.890 14.130 13.080 ;
        RECT 14.880 12.890 15.070 13.080 ;
        RECT 15.660 12.890 15.850 13.080 ;
        RECT 17.110 12.890 17.300 13.080 ;
        RECT 17.930 12.890 18.120 13.080 ;
        RECT 20.350 12.940 20.520 13.110 ;
        RECT 20.690 12.940 20.860 13.110 ;
        RECT 21.030 12.940 21.200 13.110 ;
        RECT 21.370 12.940 21.540 13.110 ;
        RECT 21.710 12.940 21.880 13.110 ;
        RECT 22.050 12.940 22.220 13.110 ;
        RECT 22.390 12.940 22.560 13.110 ;
        RECT 22.730 12.940 22.900 13.110 ;
        RECT 23.070 12.940 23.240 13.110 ;
        RECT 23.410 12.940 23.580 13.110 ;
        RECT 23.750 12.940 23.920 13.110 ;
        RECT 24.090 12.940 24.260 13.110 ;
        RECT 24.430 12.940 24.600 13.110 ;
        RECT 24.770 12.940 24.940 13.110 ;
        RECT 25.110 12.940 25.280 13.110 ;
        RECT 25.450 12.940 25.620 13.110 ;
        RECT 25.790 12.940 25.960 13.110 ;
        RECT 26.130 12.940 26.300 13.110 ;
        RECT 26.470 12.940 26.640 13.110 ;
        RECT 26.810 12.940 26.980 13.110 ;
        RECT 27.150 12.940 27.320 13.110 ;
        RECT 27.490 12.940 27.660 13.110 ;
        RECT 27.830 12.940 28.000 13.110 ;
        RECT 28.170 12.940 28.340 13.110 ;
        RECT 28.510 12.940 28.680 13.110 ;
        RECT 28.850 12.940 29.020 13.110 ;
        RECT 29.190 12.940 29.360 13.110 ;
        RECT 29.530 12.940 29.700 13.110 ;
        RECT 29.870 12.940 30.040 13.110 ;
      LAYER met1 ;
        RECT 18.420 13.260 21.630 13.270 ;
        RECT 9.350 12.780 32.170 13.260 ;
        RECT 31.380 11.650 32.170 12.780 ;
        RECT 31.380 11.640 35.600 11.650 ;
        RECT 31.380 11.240 35.620 11.640 ;
        RECT 31.380 11.230 35.130 11.240 ;
        RECT 35.280 9.960 35.620 11.240 ;
        RECT 35.870 9.960 36.180 10.180 ;
        RECT 35.280 9.340 36.180 9.960 ;
        RECT 35.870 9.270 36.180 9.340 ;
    END
  END VDD#3
  PIN REF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 3.430 5.980 4.530 6.170 ;
        RECT 3.430 5.670 3.660 5.980 ;
        RECT 1.050 2.200 1.320 3.970 ;
        RECT 1.050 1.910 3.110 2.200 ;
        RECT 1.570 1.570 1.950 1.910 ;
      LAYER mcon ;
        RECT 1.680 1.670 1.850 1.840 ;
      LAYER met1 ;
        RECT 1.600 1.600 1.920 1.920 ;
      LAYER via ;
        RECT 1.630 1.630 1.890 1.890 ;
      LAYER met2 ;
        RECT 19.180 13.430 19.950 13.710 ;
        RECT 19.420 12.780 19.700 13.430 ;
        RECT 19.370 12.410 19.750 12.780 ;
        RECT 1.570 1.570 1.950 1.950 ;
      LAYER via2 ;
        RECT 19.420 12.450 19.700 12.730 ;
        RECT 1.620 1.620 1.900 1.900 ;
      LAYER met3 ;
        RECT 7.250 12.440 19.790 12.820 ;
        RECT 7.250 10.970 7.630 12.440 ;
        RECT 19.340 12.360 19.790 12.440 ;
        RECT 7.250 9.980 7.640 10.970 ;
        RECT 5.010 9.870 7.640 9.980 ;
        RECT 5.010 9.600 7.630 9.870 ;
        RECT 5.010 4.350 5.390 9.600 ;
        RECT 3.370 3.970 5.390 4.350 ;
        RECT 3.370 1.950 3.750 3.970 ;
        RECT 1.570 1.570 3.750 1.950 ;
    END
  END REF
  OBS
      LAYER li1 ;
        RECT 9.580 12.610 9.760 12.650 ;
        RECT 9.470 11.870 9.760 12.610 ;
        RECT 10.550 12.070 10.770 12.650 ;
        RECT 9.930 11.900 10.770 12.070 ;
        RECT 9.470 11.700 9.720 11.870 ;
        RECT 9.930 11.700 10.120 11.900 ;
        RECT 9.280 11.310 9.650 11.700 ;
        RECT 9.900 11.410 10.120 11.700 ;
        RECT 10.320 11.480 10.660 11.650 ;
        RECT 11.150 11.620 11.320 12.510 ;
        RECT 12.470 11.940 12.640 12.510 ;
        RECT 9.900 11.360 10.130 11.410 ;
        RECT 9.950 11.310 10.130 11.360 ;
        RECT 10.980 11.320 11.320 11.620 ;
        RECT 12.100 11.690 12.640 11.940 ;
        RECT 11.550 11.580 11.880 11.590 ;
        RECT 12.100 11.580 12.290 11.690 ;
        RECT 11.550 11.540 12.290 11.580 ;
        RECT 11.510 11.370 12.290 11.540 ;
        RECT 11.550 11.340 12.290 11.370 ;
        RECT 9.470 11.040 9.640 11.310 ;
        RECT 9.950 11.140 10.780 11.310 ;
        RECT 9.470 10.680 9.770 11.040 ;
        RECT 10.560 10.680 10.780 11.140 ;
        RECT 11.150 10.810 11.320 11.320 ;
        RECT 12.100 11.070 12.290 11.340 ;
        RECT 12.010 10.760 12.290 11.070 ;
        RECT 12.470 10.880 12.640 11.690 ;
        RECT 12.910 11.970 13.080 12.510 ;
        RECT 12.910 11.680 13.580 11.970 ;
        RECT 12.910 10.880 13.080 11.680 ;
        RECT 13.300 11.620 13.580 11.680 ;
        RECT 13.810 11.620 13.980 12.500 ;
        RECT 15.120 11.960 15.290 12.520 ;
        RECT 13.300 11.330 13.980 11.620 ;
        RECT 14.590 11.690 15.290 11.960 ;
        RECT 14.590 11.600 14.760 11.690 ;
        RECT 14.550 11.580 14.760 11.600 ;
        RECT 14.210 11.530 14.760 11.580 ;
        RECT 14.170 11.360 14.760 11.530 ;
        RECT 14.210 11.330 14.760 11.360 ;
        RECT 13.250 10.770 13.580 10.940 ;
        RECT 13.810 10.800 13.980 11.330 ;
        RECT 15.120 10.890 15.290 11.690 ;
        RECT 15.560 11.990 15.730 12.520 ;
        RECT 16.060 12.280 16.230 12.610 ;
        RECT 15.560 11.690 16.280 11.990 ;
        RECT 15.560 10.890 15.730 11.690 ;
        RECT 16.030 11.630 16.280 11.690 ;
        RECT 16.540 11.630 16.710 12.510 ;
        RECT 16.030 11.330 16.710 11.630 ;
        RECT 17.650 11.620 17.820 12.510 ;
        RECT 16.900 11.370 17.240 11.540 ;
        RECT 16.540 10.810 16.710 11.330 ;
        RECT 17.520 11.320 17.820 11.620 ;
        RECT 21.820 11.390 21.990 11.930 ;
        RECT 17.650 10.810 17.820 11.320 ;
        RECT 22.400 11.210 22.570 12.490 ;
        RECT 22.840 12.360 23.010 12.490 ;
        RECT 22.840 12.310 23.160 12.360 ;
        RECT 22.840 11.990 29.950 12.310 ;
        RECT 22.840 11.930 23.160 11.990 ;
        RECT 22.840 11.400 23.010 11.930 ;
        RECT 21.730 10.920 22.570 11.210 ;
        RECT 23.400 11.150 23.570 11.820 ;
        RECT 23.840 11.400 24.010 11.990 ;
        RECT 24.400 11.150 24.570 11.820 ;
        RECT 24.840 11.400 25.010 11.990 ;
        RECT 25.400 11.150 25.570 11.820 ;
        RECT 25.840 11.400 26.010 11.990 ;
        RECT 26.400 11.150 26.570 11.820 ;
        RECT 26.840 11.400 27.010 11.990 ;
        RECT 27.400 11.150 27.570 11.820 ;
        RECT 27.840 11.400 28.010 11.990 ;
        RECT 28.400 11.150 28.570 11.820 ;
        RECT 28.840 11.400 29.010 11.990 ;
        RECT 22.740 10.980 23.570 11.150 ;
        RECT 23.740 10.980 24.570 11.150 ;
        RECT 24.740 10.980 25.570 11.150 ;
        RECT 25.740 10.980 26.570 11.150 ;
        RECT 26.740 10.980 27.570 11.150 ;
        RECT 27.740 10.980 28.570 11.150 ;
        RECT 28.740 10.980 29.340 11.150 ;
        RECT 19.440 10.550 19.790 10.840 ;
        RECT 19.440 10.380 21.140 10.550 ;
        RECT 1.140 9.080 1.440 9.440 ;
        RECT 1.140 8.800 1.310 9.080 ;
        RECT 2.230 8.980 2.450 9.440 ;
        RECT 0.540 8.520 1.310 8.800 ;
        RECT 1.620 8.810 2.450 8.980 ;
        RECT 1.620 8.760 1.800 8.810 ;
        RECT 2.820 8.800 2.990 9.310 ;
        RECT 3.680 9.050 3.960 9.360 ;
        RECT 0.540 2.750 0.820 8.520 ;
        RECT 1.140 8.420 1.310 8.520 ;
        RECT 1.570 8.710 1.800 8.760 ;
        RECT 1.570 8.420 1.790 8.710 ;
        RECT 1.990 8.470 2.330 8.640 ;
        RECT 2.650 8.500 2.990 8.800 ;
        RECT 3.770 8.780 3.960 9.050 ;
        RECT 3.220 8.750 3.960 8.780 ;
        RECT 3.180 8.580 3.960 8.750 ;
        RECT 3.220 8.540 3.960 8.580 ;
        RECT 3.220 8.530 3.550 8.540 ;
        RECT 1.140 8.250 1.390 8.420 ;
        RECT 1.140 7.510 1.430 8.250 ;
        RECT 1.600 8.220 1.790 8.420 ;
        RECT 1.600 8.050 2.440 8.220 ;
        RECT 1.250 7.470 1.430 7.510 ;
        RECT 2.220 7.470 2.440 8.050 ;
        RECT 2.820 7.610 2.990 8.500 ;
        RECT 3.770 8.430 3.960 8.540 ;
        RECT 4.140 8.430 4.310 9.240 ;
        RECT 3.770 8.180 4.310 8.430 ;
        RECT 3.680 7.560 3.850 7.900 ;
        RECT 4.140 7.610 4.310 8.180 ;
        RECT 4.580 8.440 4.750 9.240 ;
        RECT 4.920 9.180 5.250 9.350 ;
        RECT 5.480 8.790 5.650 9.320 ;
        RECT 4.970 8.500 5.650 8.790 ;
        RECT 5.880 8.760 6.430 8.790 ;
        RECT 5.840 8.590 6.430 8.760 ;
        RECT 5.880 8.540 6.430 8.590 ;
        RECT 6.220 8.520 6.430 8.540 ;
        RECT 4.970 8.440 5.250 8.500 ;
        RECT 4.580 8.150 5.250 8.440 ;
        RECT 4.580 7.610 4.750 8.150 ;
        RECT 5.480 7.620 5.650 8.500 ;
        RECT 6.260 8.430 6.430 8.520 ;
        RECT 6.790 8.430 6.960 9.230 ;
        RECT 6.260 8.160 6.960 8.430 ;
        RECT 6.790 7.600 6.960 8.160 ;
        RECT 7.230 8.430 7.400 9.230 ;
        RECT 7.640 9.140 7.970 9.320 ;
        RECT 8.210 8.790 8.380 9.310 ;
        RECT 9.320 8.800 9.490 9.310 ;
        RECT 7.700 8.490 8.380 8.790 ;
        RECT 8.570 8.580 8.910 8.750 ;
        RECT 9.190 8.500 9.490 8.800 ;
        RECT 11.550 9.080 11.850 9.440 ;
        RECT 9.680 8.580 10.560 8.750 ;
        RECT 7.700 8.430 7.950 8.490 ;
        RECT 7.230 8.130 7.950 8.430 ;
        RECT 7.230 7.600 7.400 8.130 ;
        RECT 7.730 7.510 7.900 7.840 ;
        RECT 8.210 7.610 8.380 8.490 ;
        RECT 9.320 7.610 9.490 8.500 ;
        RECT 10.230 8.340 10.560 8.580 ;
        RECT 11.550 8.420 11.720 9.080 ;
        RECT 12.640 8.980 12.860 9.440 ;
        RECT 12.030 8.810 12.860 8.980 ;
        RECT 12.030 8.760 12.210 8.810 ;
        RECT 13.230 8.800 13.400 9.310 ;
        RECT 14.090 9.050 14.370 9.360 ;
        RECT 11.980 8.710 12.210 8.760 ;
        RECT 11.980 8.420 12.200 8.710 ;
        RECT 12.400 8.470 12.740 8.640 ;
        RECT 13.060 8.500 13.400 8.800 ;
        RECT 14.180 8.780 14.370 9.050 ;
        RECT 13.630 8.750 14.370 8.780 ;
        RECT 13.590 8.580 14.370 8.750 ;
        RECT 13.630 8.540 14.370 8.580 ;
        RECT 13.630 8.530 13.960 8.540 ;
        RECT 11.550 8.340 11.800 8.420 ;
        RECT 10.230 8.250 11.800 8.340 ;
        RECT 10.230 8.170 11.840 8.250 ;
        RECT 11.550 7.510 11.840 8.170 ;
        RECT 12.010 8.220 12.200 8.420 ;
        RECT 12.010 8.050 12.850 8.220 ;
        RECT 11.660 7.470 11.840 7.510 ;
        RECT 12.630 7.470 12.850 8.050 ;
        RECT 13.230 7.610 13.400 8.500 ;
        RECT 14.180 8.430 14.370 8.540 ;
        RECT 14.550 8.430 14.720 9.240 ;
        RECT 14.180 8.180 14.720 8.430 ;
        RECT 14.090 7.560 14.260 7.900 ;
        RECT 14.550 7.610 14.720 8.180 ;
        RECT 14.990 8.440 15.160 9.240 ;
        RECT 15.330 9.180 15.660 9.350 ;
        RECT 15.890 8.790 16.060 9.320 ;
        RECT 15.380 8.500 16.060 8.790 ;
        RECT 16.290 8.760 16.840 8.790 ;
        RECT 16.250 8.590 16.840 8.760 ;
        RECT 16.290 8.540 16.840 8.590 ;
        RECT 16.630 8.520 16.840 8.540 ;
        RECT 15.380 8.440 15.660 8.500 ;
        RECT 14.990 8.150 15.660 8.440 ;
        RECT 14.990 7.610 15.160 8.150 ;
        RECT 15.890 7.620 16.060 8.500 ;
        RECT 16.670 8.430 16.840 8.520 ;
        RECT 17.200 8.430 17.370 9.230 ;
        RECT 16.670 8.160 17.370 8.430 ;
        RECT 17.200 7.600 17.370 8.160 ;
        RECT 17.640 8.430 17.810 9.230 ;
        RECT 18.050 9.140 18.380 9.320 ;
        RECT 18.620 8.790 18.790 9.310 ;
        RECT 19.730 8.800 19.900 9.310 ;
        RECT 18.110 8.490 18.790 8.790 ;
        RECT 18.980 8.580 19.320 8.750 ;
        RECT 19.600 8.500 19.900 8.800 ;
        RECT 20.970 8.750 21.140 10.380 ;
        RECT 20.090 8.580 21.140 8.750 ;
        RECT 18.110 8.430 18.360 8.490 ;
        RECT 17.640 8.130 18.360 8.430 ;
        RECT 17.640 7.600 17.810 8.130 ;
        RECT 18.140 7.510 18.310 7.840 ;
        RECT 18.620 7.610 18.790 8.490 ;
        RECT 19.730 7.610 19.900 8.500 ;
        RECT 21.820 7.990 21.990 10.730 ;
        RECT 22.400 8.500 22.570 10.920 ;
        RECT 22.840 10.140 23.010 10.730 ;
        RECT 23.400 10.310 23.570 10.980 ;
        RECT 23.840 10.140 24.010 10.730 ;
        RECT 24.400 10.310 24.570 10.980 ;
        RECT 24.840 10.140 25.010 10.730 ;
        RECT 25.400 10.310 25.570 10.980 ;
        RECT 25.840 10.140 26.010 10.730 ;
        RECT 26.400 10.310 26.570 10.980 ;
        RECT 26.840 10.140 27.010 10.730 ;
        RECT 27.400 10.310 27.570 10.980 ;
        RECT 27.840 10.140 28.010 10.730 ;
        RECT 28.400 10.310 28.570 10.980 ;
        RECT 28.840 10.140 29.010 10.730 ;
        RECT 22.840 9.820 29.010 10.140 ;
        RECT 22.840 9.430 23.990 9.820 ;
        RECT 25.420 9.460 26.010 9.820 ;
        RECT 22.840 8.500 23.010 9.430 ;
        RECT 25.150 9.290 26.230 9.460 ;
        RECT 26.790 9.270 27.440 9.560 ;
        RECT 29.580 9.490 29.950 11.990 ;
        RECT 32.090 9.920 33.670 10.130 ;
        RECT 31.310 9.630 31.480 9.650 ;
        RECT 24.050 8.850 26.230 9.020 ;
        RECT 21.820 7.570 23.060 7.990 ;
        RECT 24.050 7.770 24.250 8.850 ;
        RECT 26.780 8.770 27.450 9.270 ;
        RECT 27.880 9.240 29.950 9.490 ;
        RECT 31.190 9.400 31.480 9.630 ;
        RECT 30.150 9.070 30.510 9.130 ;
        RECT 27.890 8.800 28.970 8.970 ;
        RECT 29.360 8.870 30.510 9.070 ;
        RECT 30.150 8.840 30.510 8.870 ;
        RECT 24.520 8.420 24.690 8.650 ;
        RECT 26.790 8.520 27.450 8.770 ;
        RECT 28.070 8.520 28.770 8.800 ;
        RECT 26.790 8.480 28.770 8.520 ;
        RECT 29.300 8.480 29.470 8.640 ;
        RECT 24.520 7.900 25.860 8.420 ;
        RECT 26.790 8.200 29.470 8.480 ;
        RECT 24.520 7.810 24.690 7.900 ;
        RECT 29.300 7.800 29.470 8.200 ;
        RECT 29.740 7.800 29.910 8.640 ;
        RECT 31.310 8.050 31.480 9.400 ;
        RECT 31.750 8.050 31.920 9.650 ;
        RECT 32.090 7.880 32.260 9.920 ;
        RECT 32.440 8.050 32.610 9.650 ;
        RECT 33.500 8.050 33.670 9.920 ;
        RECT 31.440 7.670 32.260 7.880 ;
        RECT 33.940 7.510 34.110 8.410 ;
        RECT 33.820 7.310 34.230 7.510 ;
        RECT 2.560 5.340 3.250 5.700 ;
        RECT 1.380 5.090 3.250 5.340 ;
        RECT 3.850 5.500 4.560 5.690 ;
        RECT 1.380 4.410 1.650 5.090 ;
        RECT 3.850 5.030 4.290 5.500 ;
        RECT 6.270 5.370 6.490 6.240 ;
        RECT 6.270 5.200 7.110 5.370 ;
        RECT 7.280 5.240 7.570 6.240 ;
        RECT 10.390 5.850 29.150 6.040 ;
        RECT 17.040 5.800 17.420 5.850 ;
        RECT 18.300 5.800 18.680 5.850 ;
        RECT 20.540 5.800 20.920 5.850 ;
        RECT 9.890 5.360 10.830 5.550 ;
        RECT 11.150 5.360 29.150 5.550 ;
        RECT 17.040 5.310 17.420 5.360 ;
        RECT 18.300 5.310 18.680 5.360 ;
        RECT 6.910 5.070 7.110 5.200 ;
        RECT 3.850 4.910 6.720 5.030 ;
        RECT 1.880 4.860 6.720 4.910 ;
        RECT 1.880 4.650 4.300 4.860 ;
        RECT 6.910 4.730 7.140 5.070 ;
        RECT 6.910 4.690 7.100 4.730 ;
        RECT 6.260 4.520 7.100 4.690 ;
        RECT 1.380 4.170 4.110 4.410 ;
        RECT 6.260 4.140 6.480 4.520 ;
        RECT 7.400 4.500 7.570 5.240 ;
        RECT 7.270 4.020 7.570 4.500 ;
        RECT 10.710 4.490 10.880 4.820 ;
        RECT 11.150 4.810 17.690 4.980 ;
        RECT 20.540 4.960 20.920 5.360 ;
        RECT 16.660 4.220 16.910 4.810 ;
        RECT 17.100 4.760 17.690 4.810 ;
        RECT 20.520 4.770 20.940 4.960 ;
        RECT 17.150 4.710 17.690 4.760 ;
        RECT 17.220 4.650 17.690 4.710 ;
        RECT 17.270 4.290 17.690 4.650 ;
        RECT 19.890 4.540 20.220 4.710 ;
        RECT 20.520 4.330 29.950 4.480 ;
        RECT 16.620 4.050 16.950 4.220 ;
        RECT 19.280 3.950 29.950 4.330 ;
        RECT 19.280 3.940 20.630 3.950 ;
        RECT 29.070 3.940 29.950 3.950 ;
        RECT 0.390 2.440 0.820 2.750 ;
        RECT 1.910 2.520 2.240 2.690 ;
        RECT 3.870 1.320 4.060 3.780 ;
        RECT 4.350 2.970 4.540 3.780 ;
        RECT 5.230 3.080 5.420 3.210 ;
        RECT 4.960 2.970 5.420 3.080 ;
        RECT 4.350 2.720 5.420 2.970 ;
        RECT 4.350 2.660 4.650 2.720 ;
        RECT 4.350 1.550 4.610 2.660 ;
        RECT 4.960 2.640 5.420 2.720 ;
        RECT 5.230 2.530 5.420 2.640 ;
        RECT 5.710 2.310 5.900 3.180 ;
        RECT 6.520 2.520 6.740 3.390 ;
        RECT 6.520 2.350 7.360 2.520 ;
        RECT 7.530 2.390 7.820 3.390 ;
        RECT 5.400 2.080 5.900 2.310 ;
        RECT 7.170 2.220 7.360 2.350 ;
        RECT 6.150 2.010 6.970 2.180 ;
        RECT 7.170 1.930 7.390 2.220 ;
        RECT 4.350 1.320 4.540 1.550 ;
        RECT 4.970 1.210 5.430 1.900 ;
        RECT 7.160 1.880 7.390 1.930 ;
        RECT 7.160 1.840 7.340 1.880 ;
        RECT 6.510 1.670 7.340 1.840 ;
        RECT 6.510 1.290 6.730 1.670 ;
        RECT 7.650 1.650 7.820 2.390 ;
        RECT 10.080 2.960 10.340 3.220 ;
        RECT 9.370 2.120 9.700 2.290 ;
        RECT 7.520 1.170 7.820 1.650 ;
        RECT 9.600 1.150 9.790 1.910 ;
        RECT 10.080 1.190 10.270 2.960 ;
        RECT 18.770 2.950 18.940 3.280 ;
        RECT 19.280 3.190 19.630 3.940 ;
        RECT 19.210 3.020 19.630 3.190 ;
        RECT 10.610 2.120 10.940 2.290 ;
        RECT 11.320 2.200 11.510 2.860 ;
        RECT 12.040 2.520 12.990 2.710 ;
        RECT 19.210 2.680 19.630 2.710 ;
        RECT 18.660 2.630 19.630 2.680 ;
        RECT 13.290 2.440 19.630 2.630 ;
        RECT 10.840 1.160 11.030 1.920 ;
        RECT 11.320 1.840 12.980 2.200 ;
        RECT 13.290 1.960 19.820 2.150 ;
        RECT 11.320 1.200 11.510 1.840 ;
        RECT 18.840 1.560 19.090 1.960 ;
        RECT 19.270 1.920 19.820 1.960 ;
        RECT 19.340 1.880 19.820 1.920 ;
        RECT 19.390 1.830 19.820 1.880 ;
        RECT 19.400 1.630 19.820 1.830 ;
        RECT 18.800 1.390 19.130 1.560 ;
        RECT 19.400 1.150 19.820 1.360 ;
      LAYER mcon ;
        RECT 9.320 11.400 9.490 11.570 ;
        RECT 10.400 11.480 10.570 11.650 ;
        RECT 11.060 11.380 11.230 11.550 ;
        RECT 12.040 10.830 12.210 11.000 ;
        RECT 13.330 10.770 13.500 10.940 ;
        RECT 16.060 12.350 16.230 12.530 ;
        RECT 16.980 11.370 17.150 11.540 ;
        RECT 17.590 11.380 17.760 11.550 ;
        RECT 21.820 11.590 21.990 11.760 ;
        RECT 22.070 10.980 22.240 11.150 ;
        RECT 29.170 10.980 29.340 11.150 ;
        RECT 19.480 10.640 19.650 10.810 ;
        RECT 3.710 9.120 3.880 9.290 ;
        RECT 2.070 8.470 2.240 8.640 ;
        RECT 2.730 8.570 2.900 8.740 ;
        RECT 3.680 7.650 3.850 7.820 ;
        RECT 5.000 9.180 5.170 9.350 ;
        RECT 7.720 9.140 7.890 9.310 ;
        RECT 8.650 8.580 8.820 8.750 ;
        RECT 9.260 8.570 9.430 8.740 ;
        RECT 9.760 8.580 9.930 8.750 ;
        RECT 7.730 7.590 7.900 7.770 ;
        RECT 14.120 9.120 14.290 9.290 ;
        RECT 12.480 8.470 12.650 8.640 ;
        RECT 13.140 8.570 13.310 8.740 ;
        RECT 14.090 7.650 14.260 7.820 ;
        RECT 15.410 9.180 15.580 9.350 ;
        RECT 18.130 9.140 18.300 9.310 ;
        RECT 19.060 8.580 19.230 8.750 ;
        RECT 19.670 8.570 19.840 8.740 ;
        RECT 20.170 8.580 20.340 8.750 ;
        RECT 18.140 7.590 18.310 7.770 ;
        RECT 27.040 9.310 27.210 9.480 ;
        RECT 31.220 9.430 31.390 9.600 ;
        RECT 27.040 8.840 27.210 9.010 ;
        RECT 30.190 8.860 30.480 9.110 ;
        RECT 22.880 7.700 23.050 7.870 ;
        RECT 24.080 7.970 24.250 8.140 ;
        RECT 25.580 7.960 25.800 8.160 ;
        RECT 29.740 8.030 29.910 8.200 ;
        RECT 31.750 9.430 31.920 9.600 ;
        RECT 32.440 8.590 32.610 8.760 ;
        RECT 21.480 5.860 21.650 6.030 ;
        RECT 21.820 5.860 21.990 6.030 ;
        RECT 10.710 4.570 10.880 4.740 ;
        RECT 19.970 4.540 20.140 4.710 ;
        RECT 29.580 4.170 29.750 4.340 ;
        RECT 0.450 2.480 0.760 2.700 ;
        RECT 1.990 2.520 2.160 2.690 ;
        RECT 3.880 1.700 4.050 1.870 ;
        RECT 4.440 2.690 4.610 2.860 ;
        RECT 6.210 2.010 6.380 2.180 ;
        RECT 5.100 1.460 5.270 1.630 ;
        RECT 10.130 3.000 10.300 3.170 ;
        RECT 18.770 3.030 18.940 3.200 ;
        RECT 9.450 2.120 9.620 2.290 ;
        RECT 9.610 1.570 9.780 1.740 ;
        RECT 9.610 1.230 9.780 1.400 ;
        RECT 10.690 2.120 10.860 2.290 ;
        RECT 10.850 1.580 11.020 1.750 ;
        RECT 10.850 1.240 11.020 1.410 ;
        RECT 19.530 1.180 19.700 1.350 ;
      LAYER met1 ;
        RECT 15.980 12.280 16.300 12.600 ;
        RECT 9.230 11.320 9.580 11.660 ;
        RECT 10.320 11.430 10.630 11.710 ;
        RECT 10.330 11.060 10.600 11.430 ;
        RECT 10.980 11.320 17.210 11.600 ;
        RECT 17.490 11.300 17.840 11.650 ;
        RECT 21.250 11.530 22.050 11.820 ;
        RECT 10.330 10.790 12.270 11.060 ;
        RECT 11.950 10.770 12.270 10.790 ;
        RECT 11.950 10.760 12.260 10.770 ;
        RECT 13.260 10.690 13.590 11.020 ;
        RECT 19.400 10.570 19.720 10.890 ;
        RECT 21.250 10.290 21.450 11.530 ;
        RECT 22.040 11.200 29.400 11.210 ;
        RECT 22.030 10.920 29.400 11.200 ;
        RECT 21.140 9.810 30.110 10.290 ;
        RECT 3.620 9.350 3.930 9.360 ;
        RECT 3.620 9.330 3.940 9.350 ;
        RECT 2.000 9.060 3.940 9.330 ;
        RECT 4.930 9.100 5.260 9.430 ;
        RECT 7.630 9.080 9.980 9.370 ;
        RECT 14.030 9.350 14.340 9.360 ;
        RECT 14.030 9.330 14.350 9.350 ;
        RECT 2.000 8.690 2.270 9.060 ;
        RECT 1.990 8.410 2.300 8.690 ;
        RECT 2.650 8.520 8.880 8.800 ;
        RECT 9.160 8.470 9.510 8.820 ;
        RECT 9.700 8.790 9.980 9.080 ;
        RECT 12.410 9.060 14.350 9.330 ;
        RECT 15.340 9.100 15.670 9.430 ;
        RECT 18.040 9.080 20.390 9.370 ;
        RECT 3.620 7.990 9.020 8.240 ;
        RECT 3.620 7.570 3.910 7.990 ;
        RECT 8.770 7.880 9.020 7.990 ;
        RECT 9.700 7.880 9.990 8.790 ;
        RECT 12.410 8.690 12.680 9.060 ;
        RECT 12.400 8.410 12.710 8.690 ;
        RECT 13.060 8.520 19.290 8.800 ;
        RECT 19.570 8.470 19.920 8.820 ;
        RECT 20.110 8.790 20.390 9.080 ;
        RECT 3.620 7.560 3.900 7.570 ;
        RECT 7.650 7.520 7.970 7.840 ;
        RECT 8.770 7.560 9.990 7.880 ;
        RECT 14.030 7.990 19.430 8.240 ;
        RECT 14.030 7.570 14.320 7.990 ;
        RECT 19.180 7.880 19.430 7.990 ;
        RECT 20.110 7.880 20.400 8.790 ;
        RECT 26.780 8.770 27.450 9.810 ;
        RECT 30.630 9.370 31.450 9.660 ;
        RECT 31.690 9.370 35.020 9.660 ;
        RECT 30.630 9.190 30.900 9.370 ;
        RECT 30.050 8.820 30.900 9.190 ;
        RECT 30.050 8.770 32.670 8.820 ;
        RECT 26.790 8.760 27.440 8.770 ;
        RECT 30.610 8.530 32.670 8.770 ;
        RECT 22.810 7.920 24.310 8.190 ;
        RECT 14.030 7.560 14.310 7.570 ;
        RECT 18.060 7.520 18.380 7.840 ;
        RECT 19.180 7.560 20.400 7.880 ;
        RECT 22.820 7.640 23.110 7.920 ;
        RECT 25.520 7.900 29.970 8.260 ;
        RECT 21.420 5.800 22.100 6.090 ;
        RECT 10.630 4.490 10.950 4.810 ;
        RECT 19.890 4.480 20.210 4.780 ;
        RECT 29.510 4.100 29.830 4.420 ;
        RECT 0.390 2.470 2.220 2.750 ;
        RECT 4.350 2.600 4.700 2.950 ;
        RECT 10.050 2.920 10.370 3.240 ;
        RECT 18.690 2.950 19.010 3.270 ;
        RECT 0.390 2.440 0.820 2.470 ;
        RECT 6.140 1.930 6.460 2.250 ;
        RECT 9.380 2.040 9.700 2.360 ;
        RECT 10.610 2.040 10.930 2.360 ;
        RECT 21.350 2.000 22.140 2.750 ;
        RECT 3.820 1.690 4.800 1.930 ;
        RECT 3.820 1.640 5.330 1.690 ;
        RECT 4.570 1.400 5.330 1.640 ;
        RECT 9.570 1.450 9.820 1.800 ;
        RECT 10.810 1.450 11.060 1.810 ;
        RECT 21.350 1.450 21.830 2.000 ;
        RECT 9.570 1.150 21.830 1.450 ;
      LAYER via ;
        RECT 16.010 12.310 16.270 12.570 ;
        RECT 9.260 11.350 9.540 11.630 ;
        RECT 17.530 11.350 17.790 11.610 ;
        RECT 13.290 10.720 13.560 10.990 ;
        RECT 19.430 10.600 19.690 10.860 ;
        RECT 4.960 9.130 5.230 9.400 ;
        RECT 9.200 8.510 9.460 8.770 ;
        RECT 15.370 9.130 15.640 9.400 ;
        RECT 19.610 8.510 19.870 8.770 ;
        RECT 7.680 7.550 7.940 7.810 ;
        RECT 34.730 9.390 34.990 9.650 ;
        RECT 18.090 7.550 18.350 7.810 ;
        RECT 21.600 5.800 21.860 6.060 ;
        RECT 10.660 4.520 10.920 4.780 ;
        RECT 19.920 4.490 20.180 4.750 ;
        RECT 29.540 4.130 29.800 4.390 ;
        RECT 10.080 2.950 10.340 3.210 ;
        RECT 18.720 2.980 18.980 3.240 ;
        RECT 4.380 2.630 4.670 2.920 ;
        RECT 6.170 1.960 6.430 2.220 ;
        RECT 9.410 2.070 9.670 2.330 ;
        RECT 10.640 2.070 10.900 2.330 ;
        RECT 21.480 2.200 22.020 2.560 ;
      LAYER met2 ;
        RECT 9.210 11.290 9.600 11.680 ;
        RECT 15.980 11.630 16.300 12.570 ;
        RECT 17.490 11.650 17.820 11.720 ;
        RECT 17.490 11.630 17.840 11.650 ;
        RECT 13.270 11.340 17.840 11.630 ;
        RECT 13.270 10.990 13.600 11.340 ;
        RECT 17.490 11.300 17.840 11.340 ;
        RECT 13.260 10.930 13.600 10.990 ;
        RECT 13.260 10.690 13.590 10.930 ;
        RECT 19.370 10.540 19.750 10.920 ;
        RECT 4.930 9.190 5.260 9.430 ;
        RECT 15.340 9.190 15.670 9.430 ;
        RECT 4.930 9.130 5.270 9.190 ;
        RECT 15.340 9.130 15.680 9.190 ;
        RECT 4.940 8.780 5.270 9.130 ;
        RECT 9.160 8.780 9.510 8.820 ;
        RECT 4.940 8.490 9.510 8.780 ;
        RECT 15.350 8.780 15.680 9.130 ;
        RECT 19.570 8.780 19.920 8.820 ;
        RECT 15.350 8.490 19.920 8.780 ;
        RECT 7.650 7.550 7.970 8.490 ;
        RECT 9.160 8.470 9.510 8.490 ;
        RECT 9.160 8.400 9.490 8.470 ;
        RECT 18.060 7.550 18.380 8.490 ;
        RECT 19.570 8.470 19.920 8.490 ;
        RECT 19.570 8.400 19.900 8.470 ;
        RECT 34.700 6.860 35.020 9.660 ;
        RECT 30.320 6.540 35.020 6.860 ;
        RECT 10.510 4.790 10.950 4.810 ;
        RECT 9.270 4.490 10.950 4.790 ;
        RECT 9.270 4.430 10.940 4.490 ;
        RECT 17.370 4.460 20.210 4.780 ;
        RECT 9.270 3.180 9.590 4.430 ;
        RECT 17.370 3.460 17.840 4.460 ;
        RECT 4.350 2.920 4.700 2.950 ;
        RECT 4.350 2.650 6.410 2.920 ;
        RECT 8.680 2.870 9.590 3.180 ;
        RECT 10.050 3.060 17.840 3.460 ;
        RECT 10.050 2.920 10.370 3.060 ;
        RECT 18.140 2.950 19.010 3.270 ;
        RECT 4.350 2.600 4.700 2.650 ;
        RECT 6.150 2.250 6.410 2.650 ;
        RECT 9.270 2.360 9.590 2.870 ;
        RECT 6.140 1.930 6.460 2.250 ;
        RECT 9.270 2.040 9.700 2.360 ;
        RECT 10.430 2.070 10.930 2.360 ;
        RECT 10.430 1.560 10.760 2.070 ;
        RECT 18.140 1.560 18.510 2.950 ;
        RECT 21.450 2.170 22.060 6.090 ;
        RECT 30.320 4.420 30.670 6.540 ;
        RECT 29.510 4.100 30.670 4.420 ;
        RECT 10.430 1.550 18.510 1.560 ;
        RECT 8.680 1.190 18.510 1.550 ;
      LAYER via2 ;
        RECT 9.260 11.340 9.540 11.620 ;
        RECT 19.420 10.590 19.700 10.870 ;
      LAYER met3 ;
        RECT 8.910 11.290 9.600 11.680 ;
        RECT 8.910 10.610 9.260 11.290 ;
        RECT 19.370 10.850 19.750 10.920 ;
        RECT 19.370 10.610 19.790 10.850 ;
        RECT 8.910 10.260 19.790 10.610 ;
  END
END avsdpll_1v8
MACRO sky130_fd_io__top_power_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN P_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END P_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END P_CORE
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.050000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 11.795000 144.635000 ;
      RECT 11.095000 144.635000 21.320000 145.145000 ;
      RECT 11.095000 145.145000 12.050000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.075000 ;
      RECT 11.275000  26.075000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.705000 ;
      RECT 11.275000  81.705000 23.280000  82.180000 ;
      RECT 11.275000  82.180000 68.140000  82.215000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.810000 100.865000 68.495000 101.035000 ;
      RECT 20.810000 101.035000 21.320000 109.275000 ;
      RECT 20.810000 109.275000 68.495000 109.445000 ;
      RECT 20.810000 109.445000 21.320000 117.770000 ;
      RECT 20.810000 117.770000 68.495000 117.940000 ;
      RECT 20.810000 117.940000 21.320000 144.635000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.215000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.600000  97.890000 23.110000  98.990000 ;
      RECT 22.600000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.075000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.605000 100.840000 68.495000 100.865000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.325000 72.000000 195.000000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.950000   3.000000 72.000000   6.330000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   9.705000 11.735000   9.715000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   9.705000 11.735000   9.710000 ;
      RECT 10.710000   9.710000 11.735000   9.715000 ;
      RECT 10.710000   9.715000 11.515000   9.935000 ;
      RECT 10.720000   8.145000 11.720000   8.160000 ;
      RECT 10.780000   9.715000 11.665000   9.785000 ;
      RECT 10.790000   8.075000 11.650000   8.145000 ;
      RECT 10.850000   9.785000 11.595000   9.855000 ;
      RECT 10.860000   8.005000 11.580000   8.075000 ;
      RECT 10.920000   9.855000 11.525000   9.925000 ;
      RECT 10.930000   7.935000 11.510000   8.005000 ;
      RECT 10.930000   7.935000 11.735000   8.160000 ;
      RECT 10.930000   9.925000 11.515000   9.935000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.860000  25.500000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.500000 65.860000  29.820000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.555000 65.720000  29.765000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.820000 64.810000  30.870000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.750000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.750000 65.860000  39.875000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.805000 65.720000  39.820000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.875000 64.885000  40.850000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.730000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.730000 65.860000  49.895000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.785000 65.720000  49.840000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.895000 64.885000  50.870000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.745000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.745000 65.855000  59.880000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.800000 65.715000  59.825000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.880000 64.885000  60.850000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.735000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.735000 65.855000  69.880000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.795000 65.715000  69.825000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.880000 64.885000  70.850000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.550000  74.180000 ;
      RECT 14.030000  73.910000 65.085000  73.980000 ;
      RECT 14.030000  73.980000 65.155000  74.050000 ;
      RECT 14.030000  74.050000 65.225000  74.120000 ;
      RECT 14.030000  74.120000 65.295000  74.180000 ;
      RECT 14.030000  74.180000 65.760000  74.390000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.100000  74.180000 65.350000  74.250000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.170000  74.250000 65.425000  74.320000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.860000  74.490000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.490000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.545000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.820000 ;
      RECT 14.240000  98.840000 75.000000 129.820000 ;
      RECT 14.240000 129.820000 75.000000 130.705000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 139.825000 75.000000 140.710000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 149.825000 75.000000 150.710000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 159.825000 75.000000 160.710000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 169.825000 75.000000 170.710000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 179.825000 75.000000 180.710000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 189.825000 75.000000 190.710000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 134.795000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 144.795000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 154.795000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 164.795000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 174.795000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 184.795000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.520000 130.705000 75.000000 130.845000 ;
      RECT 15.520000 140.710000 75.000000 140.850000 ;
      RECT 15.520000 150.710000 75.000000 150.850000 ;
      RECT 15.520000 160.710000 75.000000 160.850000 ;
      RECT 15.520000 170.710000 75.000000 170.850000 ;
      RECT 15.520000 180.710000 75.000000 180.850000 ;
      RECT 15.520000 190.710000 75.000000 190.850000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.660000 133.770000 75.000000 133.910000 ;
      RECT 15.660000 143.770000 75.000000 143.910000 ;
      RECT 15.660000 153.770000 75.000000 153.910000 ;
      RECT 15.660000 163.770000 75.000000 163.910000 ;
      RECT 15.660000 173.770000 75.000000 173.910000 ;
      RECT 15.660000 183.770000 75.000000 183.910000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.140000   5.235000 17.350000   9.250000 ;
      RECT 17.140000   5.235000 17.490000   9.250000 ;
      RECT 17.140000   9.250000 17.490000   9.600000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.210000   5.165000 17.350000   5.235000 ;
      RECT 17.210000   9.250000 17.350000   9.320000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.280000   5.095000 17.350000   5.165000 ;
      RECT 17.280000   9.320000 17.350000   9.390000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.320000   5.055000 17.490000   5.235000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 65.660000  25.300000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.570000   9.680000 55.880000   9.800000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.580000 193.770000 75.000000 193.910000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.400000  19.930000 53.955000  21.835000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.600000 ;
      RECT 20.775000   1.600000 20.785000   1.760000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.555000  17.775000 53.955000  19.930000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 56.110000  17.775000 ;
      RECT 53.675000   0.000000 53.955000   7.875000 ;
      RECT 53.675000   7.875000 55.760000   9.680000 ;
      RECT 53.815000   8.000000 53.885000   8.070000 ;
      RECT 53.815000   8.070000 53.955000   8.140000 ;
      RECT 53.815000   8.140000 54.025000   8.210000 ;
      RECT 53.815000   8.210000 54.095000   8.280000 ;
      RECT 53.815000   8.280000 54.165000   8.350000 ;
      RECT 53.815000   8.350000 54.235000   8.420000 ;
      RECT 53.815000   8.420000 54.305000   8.490000 ;
      RECT 53.815000   8.490000 54.375000   8.560000 ;
      RECT 53.815000   8.560000 54.445000   8.630000 ;
      RECT 53.815000   8.630000 54.515000   8.700000 ;
      RECT 53.815000   8.700000 54.585000   8.770000 ;
      RECT 53.815000   8.770000 54.655000   8.840000 ;
      RECT 53.815000   8.840000 54.725000   8.910000 ;
      RECT 53.815000   8.910000 54.795000   8.980000 ;
      RECT 53.815000   8.980000 54.865000   9.050000 ;
      RECT 53.815000   9.050000 54.935000   9.120000 ;
      RECT 53.815000   9.120000 55.005000   9.190000 ;
      RECT 53.815000   9.190000 55.075000   9.260000 ;
      RECT 53.815000   9.260000 55.145000   9.330000 ;
      RECT 53.815000   9.330000 55.215000   9.400000 ;
      RECT 53.815000   9.400000 55.285000   9.470000 ;
      RECT 53.815000   9.470000 55.355000   9.540000 ;
      RECT 53.815000   9.540000 55.425000   9.610000 ;
      RECT 53.815000   9.610000 55.495000   9.680000 ;
      RECT 53.815000   9.680000 55.565000   9.750000 ;
      RECT 53.815000   9.750000 55.635000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.030000 ;
      RECT 55.875000  10.030000 56.110000  17.360000 ;
      RECT 68.150000  74.490000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.545000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.865000  73.770000 75.000000  74.490000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.385000 15.205000 171.495000 ;
      RECT 13.300000  94.425000 15.205000 171.595000 ;
      RECT 13.440000  94.145000 15.205000  94.385000 ;
      RECT 13.440000  94.285000 15.205000  94.425000 ;
      RECT 13.580000  94.145000 15.205000  94.285000 ;
      RECT 13.725000  94.000000 15.205000  94.145000 ;
      RECT 13.875000  93.850000 15.350000  94.000000 ;
      RECT 14.025000  93.700000 15.500000  93.850000 ;
      RECT 14.175000  93.550000 15.650000  93.700000 ;
      RECT 14.325000  93.400000 15.800000  93.550000 ;
      RECT 14.475000  93.250000 15.950000  93.400000 ;
      RECT 14.625000  93.100000 16.100000  93.250000 ;
      RECT 14.775000  92.950000 16.250000  93.100000 ;
      RECT 14.925000  92.800000 16.400000  92.950000 ;
      RECT 15.075000  92.650000 16.550000  92.800000 ;
      RECT 15.225000  92.500000 16.700000  92.650000 ;
      RECT 15.375000  92.350000 16.850000  92.500000 ;
      RECT 15.525000  92.200000 17.000000  92.350000 ;
      RECT 15.675000  92.050000 17.150000  92.200000 ;
      RECT 15.825000  91.900000 17.300000  92.050000 ;
      RECT 15.975000  91.750000 17.450000  91.900000 ;
      RECT 16.125000  91.600000 17.600000  91.750000 ;
      RECT 16.275000  91.450000 17.750000  91.600000 ;
      RECT 16.425000  91.300000 17.900000  91.450000 ;
      RECT 16.575000  91.150000 18.050000  91.300000 ;
      RECT 16.725000  91.000000 18.200000  91.150000 ;
      RECT 16.875000  90.850000 18.350000  91.000000 ;
      RECT 17.025000  90.700000 18.500000  90.850000 ;
      RECT 17.175000  90.550000 18.650000  90.700000 ;
      RECT 17.325000  90.400000 18.800000  90.550000 ;
      RECT 17.475000  90.250000 18.950000  90.400000 ;
      RECT 17.625000  90.100000 19.100000  90.250000 ;
      RECT 17.775000  89.950000 19.250000  90.100000 ;
      RECT 17.925000  89.800000 19.400000  89.950000 ;
      RECT 18.075000  89.650000 19.550000  89.800000 ;
      RECT 18.225000  89.500000 19.700000  89.650000 ;
      RECT 18.375000  89.350000 19.850000  89.500000 ;
      RECT 18.525000  89.200000 20.000000  89.350000 ;
      RECT 18.675000  89.050000 20.150000  89.200000 ;
      RECT 18.825000  88.900000 20.300000  89.050000 ;
      RECT 18.975000  88.750000 20.450000  88.900000 ;
      RECT 19.125000  88.600000 20.600000  88.750000 ;
      RECT 19.275000  88.450000 20.750000  88.600000 ;
      RECT 19.425000  88.300000 20.900000  88.450000 ;
      RECT 19.575000  88.150000 21.050000  88.300000 ;
      RECT 19.725000  88.000000 21.200000  88.150000 ;
      RECT 19.875000  87.850000 21.350000  88.000000 ;
      RECT 20.025000  87.700000 21.500000  87.850000 ;
      RECT 20.175000  87.550000 21.650000  87.700000 ;
      RECT 20.325000  87.400000 21.800000  87.550000 ;
      RECT 20.475000  87.250000 21.950000  87.400000 ;
      RECT 20.625000  87.100000 22.100000  87.250000 ;
      RECT 20.775000  86.950000 22.250000  87.100000 ;
      RECT 20.925000  86.800000 22.400000  86.950000 ;
      RECT 21.075000  86.650000 22.550000  86.800000 ;
      RECT 21.225000  86.500000 22.700000  86.650000 ;
      RECT 21.375000  86.350000 22.850000  86.500000 ;
      RECT 21.525000  86.200000 23.000000  86.350000 ;
      RECT 21.675000  86.050000 23.150000  86.200000 ;
      RECT 21.825000  85.900000 23.300000  86.050000 ;
      RECT 21.950000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000 166.935000 25.635000 170.445000 ;
      RECT 22.075000  96.885000 25.635000  96.955000 ;
      RECT 22.100000  85.625000 23.450000  85.775000 ;
      RECT 22.155000 166.935000 25.635000 167.085000 ;
      RECT 22.225000  96.735000 25.635000  96.885000 ;
      RECT 22.250000  85.475000 23.450000  85.625000 ;
      RECT 22.305000 167.085000 25.635000 167.235000 ;
      RECT 22.375000  96.585000 25.635000  96.735000 ;
      RECT 22.400000  85.325000 23.450000  85.475000 ;
      RECT 22.455000 167.235000 25.635000 167.385000 ;
      RECT 22.525000  96.435000 25.635000  96.585000 ;
      RECT 22.550000  85.175000 23.450000  85.325000 ;
      RECT 22.605000 167.385000 25.635000 167.535000 ;
      RECT 22.675000  96.285000 25.635000  96.435000 ;
      RECT 22.700000  85.025000 23.450000  85.175000 ;
      RECT 22.755000 167.535000 25.635000 167.685000 ;
      RECT 22.825000  96.135000 25.635000  96.285000 ;
      RECT 22.850000  84.875000 23.450000  85.025000 ;
      RECT 22.905000 167.685000 25.635000 167.835000 ;
      RECT 22.975000  95.985000 25.635000  96.135000 ;
      RECT 23.000000  84.725000 23.450000  84.875000 ;
      RECT 23.055000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.485000 23.450000  85.900000 ;
      RECT 23.125000  95.835000 25.635000  95.985000 ;
      RECT 23.150000  84.575000 23.450000  84.725000 ;
      RECT 23.205000 167.985000 25.635000 168.135000 ;
      RECT 23.275000  95.685000 25.635000  95.835000 ;
      RECT 23.300000  84.425000 23.450000  84.575000 ;
      RECT 23.355000 168.135000 25.635000 168.285000 ;
      RECT 23.425000  95.535000 25.635000  95.685000 ;
      RECT 23.505000 168.285000 25.635000 168.435000 ;
      RECT 23.575000  95.385000 25.635000  95.535000 ;
      RECT 23.655000 168.435000 25.635000 168.585000 ;
      RECT 23.725000  95.235000 25.635000  95.385000 ;
      RECT 23.805000 168.585000 25.635000 168.735000 ;
      RECT 23.875000  95.085000 25.635000  95.235000 ;
      RECT 23.955000 168.735000 25.635000 168.885000 ;
      RECT 24.025000  94.935000 25.635000  95.085000 ;
      RECT 24.105000 168.885000 25.635000 169.035000 ;
      RECT 24.175000  94.785000 25.635000  94.935000 ;
      RECT 24.255000 169.035000 25.635000 169.185000 ;
      RECT 24.325000  94.635000 25.635000  94.785000 ;
      RECT 24.405000 169.185000 25.635000 169.335000 ;
      RECT 24.475000  94.485000 25.635000  94.635000 ;
      RECT 24.555000 169.335000 25.635000 169.485000 ;
      RECT 24.625000  94.335000 25.635000  94.485000 ;
      RECT 24.625000  94.335000 25.635000  96.955000 ;
      RECT 24.705000 169.485000 25.635000 169.635000 ;
      RECT 24.745000  94.215000 25.635000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.335000 ;
      RECT 24.800000  82.335000 25.150000  82.785000 ;
      RECT 24.855000 169.635000 25.635000 169.785000 ;
      RECT 24.895000  94.065000 25.755000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.335000 ;
      RECT 24.900000  82.335000 25.450000  82.485000 ;
      RECT 24.900000  82.485000 25.300000  82.635000 ;
      RECT 24.900000  82.635000 25.150000  82.785000 ;
      RECT 24.900000  82.785000 25.000000  82.935000 ;
      RECT 25.005000 169.785000 25.635000 169.935000 ;
      RECT 25.045000  93.915000 25.905000  94.065000 ;
      RECT 25.155000 169.935000 25.635000 170.085000 ;
      RECT 25.195000  93.765000 26.055000  93.915000 ;
      RECT 25.305000 170.085000 25.635000 170.235000 ;
      RECT 25.345000  93.615000 26.205000  93.765000 ;
      RECT 25.455000 170.235000 25.635000 170.385000 ;
      RECT 25.495000  93.465000 26.355000  93.615000 ;
      RECT 25.515000 170.445000 25.635000 189.915000 ;
      RECT 25.605000 170.385000 25.635000 170.535000 ;
      RECT 25.645000  93.315000 26.505000  93.465000 ;
      RECT 25.795000  93.165000 26.655000  93.315000 ;
      RECT 25.945000  93.015000 26.805000  93.165000 ;
      RECT 26.095000  92.865000 26.955000  93.015000 ;
      RECT 26.245000  92.715000 27.105000  92.865000 ;
      RECT 26.395000  92.565000 27.255000  92.715000 ;
      RECT 26.545000  92.415000 27.405000  92.565000 ;
      RECT 26.695000  92.265000 27.555000  92.415000 ;
      RECT 26.845000  92.115000 27.705000  92.265000 ;
      RECT 26.995000  91.965000 27.855000  92.115000 ;
      RECT 27.145000  91.815000 28.005000  91.965000 ;
      RECT 27.295000  91.665000 28.155000  91.815000 ;
      RECT 27.445000  91.515000 28.305000  91.665000 ;
      RECT 27.595000  91.365000 28.455000  91.515000 ;
      RECT 27.745000  91.215000 28.605000  91.365000 ;
      RECT 27.895000  91.065000 28.755000  91.215000 ;
      RECT 28.045000  90.915000 28.905000  91.065000 ;
      RECT 28.195000  90.765000 29.055000  90.915000 ;
      RECT 28.345000  90.615000 29.205000  90.765000 ;
      RECT 28.495000  90.465000 29.355000  90.615000 ;
      RECT 28.645000  90.315000 29.505000  90.465000 ;
      RECT 28.795000  90.165000 29.655000  90.315000 ;
      RECT 28.945000  90.015000 29.805000  90.165000 ;
      RECT 29.095000  89.865000 29.955000  90.015000 ;
      RECT 29.245000  89.715000 30.105000  89.865000 ;
      RECT 29.395000  89.565000 30.255000  89.715000 ;
      RECT 29.545000  89.415000 30.405000  89.565000 ;
      RECT 29.695000  89.265000 30.555000  89.415000 ;
      RECT 29.845000  89.115000 30.705000  89.265000 ;
      RECT 29.995000  88.965000 30.855000  89.115000 ;
      RECT 30.145000  88.815000 31.005000  88.965000 ;
      RECT 30.295000  88.665000 31.155000  88.815000 ;
      RECT 30.445000  88.515000 31.305000  88.665000 ;
      RECT 30.595000  88.365000 31.455000  88.515000 ;
      RECT 30.745000  88.215000 31.605000  88.365000 ;
      RECT 30.895000  88.065000 31.755000  88.215000 ;
      RECT 31.045000  87.915000 31.905000  88.065000 ;
      RECT 31.195000  87.765000 32.055000  87.915000 ;
      RECT 31.345000  87.615000 32.205000  87.765000 ;
      RECT 31.495000  87.465000 32.355000  87.615000 ;
      RECT 31.645000  87.315000 32.505000  87.465000 ;
      RECT 31.795000  87.165000 32.655000  87.315000 ;
      RECT 31.945000  87.015000 32.805000  87.165000 ;
      RECT 32.095000  86.865000 32.955000  87.015000 ;
      RECT 32.245000  86.715000 33.105000  86.865000 ;
      RECT 32.395000  86.565000 33.255000  86.715000 ;
      RECT 32.435000  93.555000 40.410000  93.705000 ;
      RECT 32.435000  93.555000 42.435000  95.580000 ;
      RECT 32.435000  93.705000 40.560000  93.855000 ;
      RECT 32.435000  93.855000 40.710000  94.005000 ;
      RECT 32.435000  94.005000 40.860000  94.155000 ;
      RECT 32.435000  94.155000 41.010000  94.305000 ;
      RECT 32.435000  94.305000 41.160000  94.455000 ;
      RECT 32.435000  94.455000 41.310000  94.605000 ;
      RECT 32.435000  94.605000 41.460000  94.755000 ;
      RECT 32.435000  94.755000 41.610000  94.905000 ;
      RECT 32.435000  94.905000 41.760000  95.055000 ;
      RECT 32.435000  95.055000 41.910000  95.205000 ;
      RECT 32.435000  95.205000 42.060000  95.355000 ;
      RECT 32.435000  95.355000 42.210000  95.505000 ;
      RECT 32.435000  95.505000 42.360000  95.580000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000 162.405000 42.435000 163.970000 ;
      RECT 32.515000  93.475000 40.330000  93.555000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  85.865000 33.555000  86.415000 ;
      RECT 32.545000  85.865000 33.955000  86.015000 ;
      RECT 32.545000  86.015000 33.805000  86.165000 ;
      RECT 32.545000  86.165000 33.655000  86.315000 ;
      RECT 32.545000  86.315000 33.555000  86.415000 ;
      RECT 32.545000  86.415000 33.405000  86.565000 ;
      RECT 32.570000  84.830000 34.080000  84.855000 ;
      RECT 32.585000 162.405000 42.435000 162.555000 ;
      RECT 32.665000  93.325000 40.180000  93.475000 ;
      RECT 32.720000  84.680000 33.930000  84.830000 ;
      RECT 32.735000 162.555000 42.435000 162.705000 ;
      RECT 32.815000  93.175000 40.030000  93.325000 ;
      RECT 32.870000  84.530000 33.780000  84.680000 ;
      RECT 32.885000 162.705000 42.435000 162.855000 ;
      RECT 32.965000  93.025000 39.880000  93.175000 ;
      RECT 33.020000  84.380000 33.630000  84.530000 ;
      RECT 33.020000  84.380000 34.105000  84.855000 ;
      RECT 33.035000 162.855000 42.435000 163.005000 ;
      RECT 33.115000  92.875000 39.730000  93.025000 ;
      RECT 33.185000 163.005000 42.435000 163.155000 ;
      RECT 33.265000  92.725000 39.580000  92.875000 ;
      RECT 33.335000 163.155000 42.435000 163.305000 ;
      RECT 33.415000  92.575000 39.430000  92.725000 ;
      RECT 33.485000 163.305000 42.435000 163.455000 ;
      RECT 33.565000  92.425000 39.280000  92.575000 ;
      RECT 33.635000 163.455000 42.435000 163.605000 ;
      RECT 33.715000  92.275000 39.130000  92.425000 ;
      RECT 33.785000 163.605000 42.435000 163.755000 ;
      RECT 33.865000  92.125000 38.980000  92.275000 ;
      RECT 33.935000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.905000 42.435000 163.970000 ;
      RECT 34.000000 163.970000 39.110000 167.295000 ;
      RECT 34.015000  91.975000 38.830000  92.125000 ;
      RECT 34.150000 163.970000 42.285000 164.120000 ;
      RECT 34.165000  91.825000 38.680000  91.975000 ;
      RECT 34.300000 164.120000 42.135000 164.270000 ;
      RECT 34.315000  91.675000 38.530000  91.825000 ;
      RECT 34.450000 164.270000 41.985000 164.420000 ;
      RECT 34.465000  91.525000 38.380000  91.675000 ;
      RECT 34.600000 164.420000 41.835000 164.570000 ;
      RECT 34.615000  91.375000 38.230000  91.525000 ;
      RECT 34.750000 164.570000 41.685000 164.720000 ;
      RECT 34.765000  91.225000 38.080000  91.375000 ;
      RECT 34.900000 164.720000 41.535000 164.870000 ;
      RECT 34.915000  91.075000 37.930000  91.225000 ;
      RECT 35.050000 164.870000 41.385000 165.020000 ;
      RECT 35.065000  90.925000 37.780000  91.075000 ;
      RECT 35.200000 165.020000 41.235000 165.170000 ;
      RECT 35.215000  90.775000 37.630000  90.925000 ;
      RECT 35.215000  90.775000 40.410000  93.555000 ;
      RECT 35.350000 165.170000 41.085000 165.320000 ;
      RECT 35.500000 165.320000 40.935000 165.470000 ;
      RECT 35.650000 165.470000 40.785000 165.620000 ;
      RECT 35.800000 165.620000 40.635000 165.770000 ;
      RECT 35.950000 165.770000 40.485000 165.920000 ;
      RECT 36.100000 165.920000 40.335000 166.070000 ;
      RECT 36.250000 166.070000 40.185000 166.220000 ;
      RECT 36.400000 166.220000 40.035000 166.370000 ;
      RECT 36.550000 166.370000 39.885000 166.520000 ;
      RECT 36.700000 166.520000 39.735000 166.670000 ;
      RECT 36.850000 166.670000 39.585000 166.820000 ;
      RECT 37.000000 166.820000 39.435000 166.970000 ;
      RECT 37.150000 166.970000 39.285000 167.120000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.940000 ;
      RECT 37.280000  69.890000 50.455000  70.940000 ;
      RECT 37.280000  70.940000 50.455000  74.340000 ;
      RECT 37.300000 167.120000 39.135000 167.270000 ;
      RECT 37.325000 167.270000 39.110000 167.295000 ;
      RECT 37.325000 167.295000 37.545000 168.860000 ;
      RECT 37.325000 167.295000 38.960000 167.445000 ;
      RECT 37.325000 167.445000 38.810000 167.595000 ;
      RECT 37.325000 167.595000 38.660000 167.745000 ;
      RECT 37.325000 167.745000 38.510000 167.895000 ;
      RECT 37.325000 167.895000 38.360000 168.045000 ;
      RECT 37.325000 168.045000 38.210000 168.195000 ;
      RECT 37.325000 168.195000 38.060000 168.345000 ;
      RECT 37.325000 168.345000 37.910000 168.495000 ;
      RECT 37.325000 168.495000 37.760000 168.645000 ;
      RECT 37.325000 168.645000 37.610000 168.795000 ;
      RECT 37.325000 168.795000 37.460000 168.945000 ;
      RECT 37.325000 168.860000 37.545000 189.915000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  87.195000 41.210000  87.610000 ;
      RECT 39.810000  84.830000 41.185000  84.855000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.935000  87.195000 41.210000  87.345000 ;
      RECT 39.960000  84.680000 41.035000  84.830000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 40.085000  87.345000 41.210000  87.495000 ;
      RECT 40.110000  84.530000 40.885000  84.680000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.200000  87.495000 41.210000  87.610000 ;
      RECT 40.200000  87.610000 50.245000  96.645000 ;
      RECT 40.260000  84.380000 40.735000  84.530000 ;
      RECT 40.260000  84.380000 41.210000  84.855000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.350000  87.610000 41.210000  87.760000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.500000  87.760000 41.360000  87.910000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.650000  87.910000 41.510000  88.060000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.800000  88.060000 41.660000  88.210000 ;
      RECT 40.950000  88.210000 41.810000  88.360000 ;
      RECT 41.100000  88.360000 41.960000  88.510000 ;
      RECT 41.250000  88.510000 42.110000  88.660000 ;
      RECT 41.400000  88.660000 42.260000  88.810000 ;
      RECT 41.550000  88.810000 42.410000  88.960000 ;
      RECT 41.700000  88.960000 42.560000  89.110000 ;
      RECT 41.850000  89.110000 42.710000  89.260000 ;
      RECT 42.000000  89.260000 42.860000  89.410000 ;
      RECT 42.150000  89.410000 43.010000  89.560000 ;
      RECT 42.300000  89.560000 43.160000  89.710000 ;
      RECT 42.450000  89.710000 43.310000  89.860000 ;
      RECT 42.600000  89.860000 43.460000  90.010000 ;
      RECT 42.750000  90.010000 43.610000  90.160000 ;
      RECT 42.900000  90.160000 43.760000  90.310000 ;
      RECT 43.050000  90.310000 43.910000  90.460000 ;
      RECT 43.200000  90.460000 44.060000  90.610000 ;
      RECT 43.350000  90.610000 44.210000  90.760000 ;
      RECT 43.500000  90.760000 44.360000  90.910000 ;
      RECT 43.650000  90.910000 44.510000  91.060000 ;
      RECT 43.800000  91.060000 44.660000  91.210000 ;
      RECT 43.950000  91.210000 44.810000  91.360000 ;
      RECT 44.100000  91.360000 44.960000  91.510000 ;
      RECT 44.250000  91.510000 45.110000  91.660000 ;
      RECT 44.400000  91.660000 45.260000  91.810000 ;
      RECT 44.550000  91.810000 45.410000  91.960000 ;
      RECT 44.700000  91.960000 45.560000  92.110000 ;
      RECT 44.850000  92.110000 45.710000  92.260000 ;
      RECT 45.000000  92.260000 45.860000  92.410000 ;
      RECT 45.150000  92.410000 46.010000  92.560000 ;
      RECT 45.300000  92.560000 46.160000  92.710000 ;
      RECT 45.450000  92.710000 46.310000  92.860000 ;
      RECT 45.600000  92.860000 46.460000  93.010000 ;
      RECT 45.750000  93.010000 46.610000  93.160000 ;
      RECT 45.900000  93.160000 46.760000  93.310000 ;
      RECT 46.050000  93.310000 46.910000  93.460000 ;
      RECT 46.200000  93.460000 47.060000  93.610000 ;
      RECT 46.350000  93.610000 47.210000  93.760000 ;
      RECT 46.500000  93.760000 47.360000  93.910000 ;
      RECT 46.650000  93.910000 47.510000  94.060000 ;
      RECT 46.800000  94.060000 47.660000  94.210000 ;
      RECT 46.950000  94.210000 47.810000  94.360000 ;
      RECT 46.960000  74.340000 50.455000  76.650000 ;
      RECT 47.100000  94.360000 47.960000  94.510000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.250000  94.510000 48.110000  94.660000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.400000  94.660000 48.260000  94.810000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.550000  94.810000 48.410000  94.960000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.700000  94.960000 48.560000  95.110000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.850000  95.110000 48.710000  95.260000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 48.000000  95.260000 48.860000  95.410000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.150000  95.410000 49.010000  95.560000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.300000  95.560000 49.160000  95.710000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.450000  95.710000 49.310000  95.860000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.600000  95.860000 49.460000  96.010000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.750000  96.010000 49.610000  96.160000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.900000  96.160000 49.760000  96.310000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 49.050000  96.310000 49.910000  96.460000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.200000  96.460000 50.060000  96.610000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.610000 50.210000  96.645000 ;
      RECT 49.235000  96.645000 50.245000  96.795000 ;
      RECT 49.235000  96.645000 53.930000 100.330000 ;
      RECT 49.235000  96.795000 50.395000  96.945000 ;
      RECT 49.235000  96.945000 50.545000  97.095000 ;
      RECT 49.235000  97.095000 50.695000  97.245000 ;
      RECT 49.235000  97.245000 50.845000  97.395000 ;
      RECT 49.235000  97.395000 50.995000  97.545000 ;
      RECT 49.235000  97.545000 51.145000  97.695000 ;
      RECT 49.235000  97.695000 51.295000  97.845000 ;
      RECT 49.235000  97.845000 51.445000  97.995000 ;
      RECT 49.235000  97.995000 51.595000  98.145000 ;
      RECT 49.235000  98.145000 51.745000  98.295000 ;
      RECT 49.235000  98.295000 51.895000  98.445000 ;
      RECT 49.235000  98.445000 52.045000  98.595000 ;
      RECT 49.235000  98.595000 52.195000  98.745000 ;
      RECT 49.235000  98.745000 52.345000  98.895000 ;
      RECT 49.235000  98.895000 52.495000  99.045000 ;
      RECT 49.235000  99.045000 52.645000  99.195000 ;
      RECT 49.235000  99.195000 52.795000  99.345000 ;
      RECT 49.235000  99.345000 52.945000  99.495000 ;
      RECT 49.235000  99.495000 53.095000  99.645000 ;
      RECT 49.235000  99.645000 53.245000  99.795000 ;
      RECT 49.235000  99.795000 53.395000  99.945000 ;
      RECT 49.235000  99.945000 53.545000 100.095000 ;
      RECT 49.235000 100.095000 53.695000 100.245000 ;
      RECT 49.235000 100.245000 53.845000 100.330000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 164.295000 49.470000 168.755000 ;
      RECT 49.235000 164.295000 53.780000 164.445000 ;
      RECT 49.235000 164.445000 53.630000 164.595000 ;
      RECT 49.235000 164.595000 53.480000 164.745000 ;
      RECT 49.235000 164.745000 53.330000 164.895000 ;
      RECT 49.235000 164.895000 53.180000 165.045000 ;
      RECT 49.235000 165.045000 53.030000 165.195000 ;
      RECT 49.235000 165.195000 52.880000 165.345000 ;
      RECT 49.235000 165.345000 52.730000 165.495000 ;
      RECT 49.235000 165.495000 52.580000 165.645000 ;
      RECT 49.235000 165.645000 52.430000 165.795000 ;
      RECT 49.235000 165.795000 52.280000 165.945000 ;
      RECT 49.235000 165.945000 52.130000 166.095000 ;
      RECT 49.235000 166.095000 51.980000 166.245000 ;
      RECT 49.235000 166.245000 51.830000 166.395000 ;
      RECT 49.235000 166.395000 51.680000 166.545000 ;
      RECT 49.235000 166.545000 51.530000 166.695000 ;
      RECT 49.235000 166.695000 51.380000 166.845000 ;
      RECT 49.235000 166.845000 51.230000 166.995000 ;
      RECT 49.235000 166.995000 51.080000 167.145000 ;
      RECT 49.235000 167.145000 50.930000 167.295000 ;
      RECT 49.235000 167.295000 50.780000 167.445000 ;
      RECT 49.235000 167.445000 50.630000 167.595000 ;
      RECT 49.235000 167.595000 50.480000 167.745000 ;
      RECT 49.235000 167.745000 50.330000 167.895000 ;
      RECT 49.235000 167.895000 50.180000 168.045000 ;
      RECT 49.235000 168.045000 50.030000 168.195000 ;
      RECT 49.235000 168.195000 49.880000 168.345000 ;
      RECT 49.235000 168.345000 49.730000 168.495000 ;
      RECT 49.235000 168.495000 49.580000 168.645000 ;
      RECT 49.235000 168.645000 49.430000 168.795000 ;
      RECT 49.235000 168.755000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.280000 168.945000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.650000 50.455000  84.590000 ;
      RECT 49.270000  77.735000 50.355000  84.630000 ;
      RECT 49.270000  84.590000 50.510000  84.645000 ;
      RECT 49.270000  84.630000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.360000  84.640000 ;
      RECT 49.270000  84.640000 50.365000  84.645000 ;
      RECT 49.270000  84.645000 52.660000  86.795000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  84.645000 50.370000  84.795000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  84.795000 50.520000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  84.945000 50.670000  85.095000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  85.095000 50.820000  85.245000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  85.245000 50.970000  85.395000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  85.395000 51.120000  85.545000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  85.545000 51.270000  85.695000 ;
      RECT 50.470000  85.695000 51.420000  85.845000 ;
      RECT 50.620000  85.845000 51.570000  85.995000 ;
      RECT 50.770000  85.995000 51.720000  86.145000 ;
      RECT 50.920000  86.145000 51.870000  86.295000 ;
      RECT 51.070000  86.295000 52.020000  86.445000 ;
      RECT 51.220000  86.445000 52.170000  86.595000 ;
      RECT 51.370000  86.595000 52.320000  86.745000 ;
      RECT 51.420000  86.745000 52.470000  86.795000 ;
      RECT 51.420000  86.795000 52.520000  86.945000 ;
      RECT 51.420000  86.795000 54.075000  88.210000 ;
      RECT 51.420000  86.945000 52.670000  87.095000 ;
      RECT 51.420000  87.095000 52.820000  87.245000 ;
      RECT 51.420000  87.245000 52.970000  87.395000 ;
      RECT 51.420000  87.395000 53.120000  87.545000 ;
      RECT 51.420000  87.545000 53.270000  87.695000 ;
      RECT 51.420000  87.695000 53.420000  87.845000 ;
      RECT 51.420000  87.845000 53.570000  87.995000 ;
      RECT 51.420000  87.995000 53.720000  88.145000 ;
      RECT 51.420000  88.145000 53.870000  88.210000 ;
      RECT 51.420000  88.210000 61.745000  95.880000 ;
      RECT 51.570000  88.210000 53.935000  88.360000 ;
      RECT 51.720000  88.360000 54.085000  88.510000 ;
      RECT 51.870000  88.510000 54.235000  88.660000 ;
      RECT 52.020000  88.660000 54.385000  88.810000 ;
      RECT 52.170000  88.810000 54.535000  88.960000 ;
      RECT 52.320000  88.960000 54.685000  89.110000 ;
      RECT 52.470000  89.110000 54.835000  89.260000 ;
      RECT 52.620000  89.260000 54.985000  89.410000 ;
      RECT 52.770000  89.410000 55.135000  89.560000 ;
      RECT 52.920000  89.560000 55.285000  89.710000 ;
      RECT 53.070000  89.710000 55.435000  89.860000 ;
      RECT 53.220000  89.860000 55.585000  90.010000 ;
      RECT 53.370000  90.010000 55.735000  90.160000 ;
      RECT 53.520000  90.160000 55.885000  90.310000 ;
      RECT 53.670000  90.310000 56.035000  90.460000 ;
      RECT 53.820000  90.460000 56.185000  90.610000 ;
      RECT 53.970000  90.610000 56.335000  90.760000 ;
      RECT 54.120000  90.760000 56.485000  90.910000 ;
      RECT 54.270000  90.910000 56.635000  91.060000 ;
      RECT 54.420000  91.060000 56.785000  91.210000 ;
      RECT 54.570000  91.210000 56.935000  91.360000 ;
      RECT 54.720000  91.360000 57.085000  91.510000 ;
      RECT 54.870000  91.510000 57.235000  91.660000 ;
      RECT 55.020000  91.660000 57.385000  91.810000 ;
      RECT 55.170000  91.810000 57.535000  91.960000 ;
      RECT 55.320000  91.960000 57.685000  92.110000 ;
      RECT 55.470000  92.110000 57.835000  92.260000 ;
      RECT 55.620000  92.260000 57.985000  92.410000 ;
      RECT 55.770000  92.410000 58.135000  92.560000 ;
      RECT 55.920000  92.560000 58.285000  92.710000 ;
      RECT 56.070000  92.710000 58.435000  92.860000 ;
      RECT 56.220000  92.860000 58.585000  93.010000 ;
      RECT 56.370000  93.010000 58.735000  93.160000 ;
      RECT 56.520000  93.160000 58.885000  93.310000 ;
      RECT 56.670000  93.310000 59.035000  93.460000 ;
      RECT 56.820000  93.460000 59.185000  93.610000 ;
      RECT 56.970000  93.610000 59.335000  93.760000 ;
      RECT 57.120000  93.760000 59.485000  93.910000 ;
      RECT 57.270000  93.910000 59.635000  94.060000 ;
      RECT 57.420000  94.060000 59.785000  94.210000 ;
      RECT 57.570000  94.210000 59.935000  94.360000 ;
      RECT 57.720000  94.360000 60.085000  94.510000 ;
      RECT 57.870000  94.510000 60.235000  94.660000 ;
      RECT 58.020000  94.660000 60.385000  94.810000 ;
      RECT 58.170000  94.810000 60.535000  94.960000 ;
      RECT 58.320000  94.960000 60.685000  95.110000 ;
      RECT 58.470000  95.110000 60.835000  95.260000 ;
      RECT 58.620000  95.260000 60.985000  95.410000 ;
      RECT 58.770000  95.410000 61.135000  95.560000 ;
      RECT 58.920000  95.560000 61.285000  95.710000 ;
      RECT 59.070000  95.710000 61.435000  95.860000 ;
      RECT 59.090000  95.880000 61.745000  97.520000 ;
      RECT 59.130000  95.860000 61.585000  95.920000 ;
      RECT 59.280000  95.920000 61.645000  96.070000 ;
      RECT 59.430000  96.070000 61.645000  96.220000 ;
      RECT 59.580000  96.220000 61.645000  96.370000 ;
      RECT 59.730000  96.370000 61.645000  96.520000 ;
      RECT 59.880000  96.520000 61.645000  96.670000 ;
      RECT 60.030000  96.670000 61.645000  96.820000 ;
      RECT 60.180000  96.820000 61.645000  96.970000 ;
      RECT 60.330000  96.970000 61.645000  97.120000 ;
      RECT 60.480000  97.120000 61.645000  97.270000 ;
      RECT 60.630000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.420000 61.645000  97.520000 ;
      RECT 60.730000  97.520000 61.645000 172.635000 ;
      RECT 60.730000  97.520000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000   5.885000 75.000000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  11.935000 75.000000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  16.785000 75.000000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  22.835000 75.000000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  28.885000 75.000000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  33.735000 75.000000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  38.585000 75.000000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  44.635000 75.000000  45.435000 ;
      RECT  0.000000  55.035000 75.000000  55.835000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  61.085000 75.000000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  66.935000 75.000000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.570000  45.435000 73.430000  55.035000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000  17.385000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT  0.000000  94.585000 75.000000 161.165000 ;
      RECT  0.000000 161.165000 30.095000 168.720000 ;
      RECT  0.000000 168.720000 75.000000 172.185000 ;
      RECT  2.565000  13.035000 72.435000  16.285000 ;
      RECT  2.870000   0.000000 72.130000  13.035000 ;
      RECT  2.870000  16.285000 72.130000  94.585000 ;
      RECT  2.870000 172.185000 72.130000 198.000000 ;
      RECT 53.940000 161.165000 75.000000 168.720000 ;
  END
END sky130_fd_io__top_power_lvc_wpad
MACRO simple_por
  CLASS BLOCK ;
  FOREIGN simple_por ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.800 BY 45.820 ;
  PIN porb_h
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.840 41.820 4.120 45.820 ;
    END
  END porb_h
  PIN vdd3v3
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.000 0.280 4.000 ;
    END
  END vdd3v3
  PIN vss
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 17.800 19.310 21.800 19.910 ;
    END
  END vss
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2.780 17.260 15.740 18.860 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2.780 19.295 15.740 20.895 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 2.780 16.195 15.740 28.575 ;
      LAYER met1 ;
        RECT 2.780 16.025 15.740 28.745 ;
      LAYER met2 ;
        RECT 4.400 41.540 14.320 41.820 ;
        RECT 3.850 16.025 14.320 41.540 ;
      LAYER met3 ;
        RECT 4.140 16.115 14.380 28.655 ;
      LAYER met4 ;
        RECT 4.140 16.025 14.380 28.745 ;
      LAYER met5 ;
        RECT 2.780 22.495 15.740 27.000 ;
  END
END simple_por
MACRO sky130_fd_io__top_ground_hvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  284.1730 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 36.645000 139.325000 37.970000 145.935000 ;
    END
  END G_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.620000 185.295000 74.290000 190.015000 ;
        RECT 16.805000  47.455000 74.290000  54.765000 ;
        RECT 16.805000 139.455000 74.290000 146.710000 ;
        RECT 16.805000 162.455000 74.290000 171.155000 ;
        RECT 16.875000 146.710000 74.290000 146.780000 ;
        RECT 16.945000 146.780000 74.290000 146.850000 ;
        RECT 17.015000 146.850000 74.290000 146.920000 ;
        RECT 17.085000 146.920000 74.290000 146.990000 ;
        RECT 17.155000 146.990000 74.290000 147.060000 ;
        RECT 17.225000 147.060000 74.290000 147.130000 ;
        RECT 17.295000 147.130000 74.290000 147.200000 ;
        RECT 17.365000 147.200000 74.290000 147.270000 ;
        RECT 17.435000 147.270000 74.290000 147.340000 ;
        RECT 17.505000 147.340000 74.290000 147.410000 ;
        RECT 17.530000  54.765000 74.290000  54.835000 ;
        RECT 17.575000 147.410000 74.290000 147.480000 ;
        RECT 17.600000  54.835000 74.290000  54.905000 ;
        RECT 17.645000 147.480000 74.290000 147.550000 ;
        RECT 17.670000  54.905000 74.290000  54.975000 ;
        RECT 17.715000 147.550000 74.290000 147.620000 ;
        RECT 17.740000  54.975000 74.290000  55.045000 ;
        RECT 17.785000 147.620000 74.290000 147.690000 ;
        RECT 17.810000  55.045000 74.290000  55.115000 ;
        RECT 17.855000 147.690000 74.290000 147.760000 ;
        RECT 17.880000  55.115000 74.290000  55.185000 ;
        RECT 17.925000 147.760000 74.290000 147.830000 ;
        RECT 17.950000  55.185000 74.290000  55.255000 ;
        RECT 17.995000 147.830000 74.290000 147.900000 ;
        RECT 18.020000  55.255000 74.290000  55.325000 ;
        RECT 18.065000 147.900000 74.290000 147.970000 ;
        RECT 18.090000  55.325000 74.290000  55.395000 ;
        RECT 18.135000 147.970000 74.290000 148.040000 ;
        RECT 18.160000  55.395000 74.290000  55.465000 ;
        RECT 18.205000 148.040000 74.290000 148.110000 ;
        RECT 18.230000  55.465000 74.290000  55.535000 ;
        RECT 18.250000 148.110000 74.290000 148.155000 ;
        RECT 18.300000  55.535000 74.290000  55.605000 ;
        RECT 18.370000  55.605000 74.290000  55.675000 ;
        RECT 18.410000  74.155000 74.290000  74.415000 ;
        RECT 18.440000  55.675000 74.290000  55.745000 ;
        RECT 18.510000  55.745000 74.290000  55.815000 ;
        RECT 18.580000  55.815000 74.290000  55.885000 ;
        RECT 18.650000  55.885000 74.290000  55.955000 ;
        RECT 18.720000  55.955000 74.290000  56.025000 ;
        RECT 18.790000  56.025000 74.290000  56.095000 ;
        RECT 18.850000  56.095000 74.290000  56.155000 ;
        RECT 23.690000  74.415000 74.290000  74.485000 ;
        RECT 23.700000  74.105000 74.290000  74.155000 ;
        RECT 23.760000  74.485000 74.290000  74.555000 ;
        RECT 23.770000  74.035000 74.290000  74.105000 ;
        RECT 23.830000  74.555000 74.290000  74.625000 ;
        RECT 23.840000  73.965000 74.290000  74.035000 ;
        RECT 23.900000  74.625000 74.290000  74.695000 ;
        RECT 23.910000  73.895000 74.290000  73.965000 ;
        RECT 23.970000  74.695000 74.290000  74.765000 ;
        RECT 23.980000  73.825000 74.290000  73.895000 ;
        RECT 24.040000  74.765000 74.290000  74.835000 ;
        RECT 24.050000  73.755000 74.290000  73.825000 ;
        RECT 24.110000  74.835000 74.290000  74.905000 ;
        RECT 24.120000  73.685000 74.290000  73.755000 ;
        RECT 24.180000  74.905000 74.290000  74.975000 ;
        RECT 24.190000  73.615000 74.290000  73.685000 ;
        RECT 24.250000  74.975000 74.290000  75.045000 ;
        RECT 24.260000  73.545000 74.290000  73.615000 ;
        RECT 24.320000  75.045000 74.290000  75.115000 ;
        RECT 24.330000  73.475000 74.290000  73.545000 ;
        RECT 24.390000  75.115000 74.290000  75.185000 ;
        RECT 24.400000  73.405000 74.290000  73.475000 ;
        RECT 24.460000  75.185000 74.290000  75.255000 ;
        RECT 24.470000  73.335000 74.290000  73.405000 ;
        RECT 24.530000  75.255000 74.290000  75.325000 ;
        RECT 24.540000  73.265000 74.290000  73.335000 ;
        RECT 24.600000  75.325000 74.290000  75.395000 ;
        RECT 24.610000  73.195000 74.290000  73.265000 ;
        RECT 24.670000  75.395000 74.290000  75.465000 ;
        RECT 24.680000  73.125000 74.290000  73.195000 ;
        RECT 24.740000  75.465000 74.290000  75.535000 ;
        RECT 24.750000  73.055000 74.290000  73.125000 ;
        RECT 24.810000  75.535000 74.290000  75.605000 ;
        RECT 24.820000  70.455000 74.290000  72.985000 ;
        RECT 24.820000  72.985000 74.290000  73.055000 ;
        RECT 24.820000  75.605000 74.290000  75.615000 ;
        RECT 24.820000  75.615000 74.290000  79.155000 ;
        RECT 24.820000  93.455000 74.290000 102.155000 ;
        RECT 24.820000 116.455000 74.290000 125.155000 ;
        RECT 37.890000  12.295000 74.290000  25.660000 ;
        RECT 46.750000  12.265000 74.290000  12.295000 ;
        RECT 46.820000  12.195000 74.290000  12.265000 ;
        RECT 46.890000  12.125000 74.290000  12.195000 ;
        RECT 46.960000  12.055000 74.290000  12.125000 ;
        RECT 47.030000  11.985000 74.290000  12.055000 ;
        RECT 47.100000  11.915000 74.290000  11.985000 ;
        RECT 47.170000  11.845000 74.290000  11.915000 ;
        RECT 47.240000  11.775000 74.290000  11.845000 ;
        RECT 47.310000  11.705000 74.290000  11.775000 ;
        RECT 47.380000  11.635000 74.290000  11.705000 ;
        RECT 47.450000  11.565000 74.290000  11.635000 ;
        RECT 47.520000  11.495000 74.290000  11.565000 ;
        RECT 47.590000  11.425000 74.290000  11.495000 ;
        RECT 47.660000  11.355000 74.290000  11.425000 ;
        RECT 47.730000  11.285000 74.290000  11.355000 ;
        RECT 47.800000  11.215000 74.290000  11.285000 ;
        RECT 47.870000  11.145000 74.290000  11.215000 ;
        RECT 47.940000  11.075000 74.290000  11.145000 ;
        RECT 48.010000  11.005000 74.290000  11.075000 ;
        RECT 48.080000  10.935000 74.290000  11.005000 ;
        RECT 48.150000  10.865000 74.290000  10.935000 ;
        RECT 48.220000  10.795000 74.290000  10.865000 ;
        RECT 48.290000  10.725000 74.290000  10.795000 ;
        RECT 48.360000  10.655000 74.290000  10.725000 ;
        RECT 48.430000  10.585000 74.290000  10.655000 ;
        RECT 48.500000  10.515000 74.290000  10.585000 ;
        RECT 48.570000  10.445000 74.290000  10.515000 ;
        RECT 48.640000  10.375000 74.290000  10.445000 ;
        RECT 48.710000  10.305000 74.290000  10.375000 ;
        RECT 48.780000  10.235000 74.290000  10.305000 ;
        RECT 48.850000  10.165000 74.290000  10.235000 ;
        RECT 48.920000  10.095000 74.290000  10.165000 ;
        RECT 48.990000  10.025000 74.290000  10.095000 ;
        RECT 49.060000   9.955000 74.290000  10.025000 ;
        RECT 49.130000   9.885000 74.290000   9.955000 ;
        RECT 49.200000   9.815000 74.290000   9.885000 ;
        RECT 49.270000   9.745000 74.290000   9.815000 ;
        RECT 49.340000   9.675000 74.290000   9.745000 ;
        RECT 49.410000   9.605000 74.290000   9.675000 ;
        RECT 49.480000   9.535000 74.290000   9.605000 ;
        RECT 49.550000   9.465000 74.290000   9.535000 ;
        RECT 49.620000   9.395000 74.290000   9.465000 ;
        RECT 49.690000   9.325000 74.290000   9.395000 ;
        RECT 49.760000   9.255000 74.290000   9.325000 ;
        RECT 49.830000   9.185000 74.290000   9.255000 ;
        RECT 49.900000   9.115000 74.290000   9.185000 ;
        RECT 49.970000   9.045000 74.290000   9.115000 ;
        RECT 50.040000   8.975000 74.290000   9.045000 ;
        RECT 50.110000   8.905000 74.290000   8.975000 ;
        RECT 50.180000   8.835000 74.290000   8.905000 ;
        RECT 50.250000   8.765000 74.290000   8.835000 ;
        RECT 50.320000   8.695000 74.290000   8.765000 ;
        RECT 50.390000   0.000000 74.290000   8.625000 ;
        RECT 50.390000   8.625000 74.290000   8.695000 ;
        RECT 55.885000  25.660000 74.290000  25.730000 ;
        RECT 55.955000  25.730000 74.290000  25.800000 ;
        RECT 56.025000  25.800000 74.290000  25.870000 ;
        RECT 56.095000  25.870000 74.290000  25.940000 ;
        RECT 56.165000  25.940000 74.290000  26.010000 ;
        RECT 56.235000  26.010000 74.290000  26.080000 ;
        RECT 56.305000  26.080000 74.290000  26.150000 ;
        RECT 56.375000  26.150000 74.290000  26.220000 ;
        RECT 56.445000  26.220000 74.290000  26.290000 ;
        RECT 56.515000  26.290000 74.290000  26.360000 ;
        RECT 56.585000  26.360000 74.290000  26.430000 ;
        RECT 56.655000  26.430000 74.290000  26.500000 ;
        RECT 56.725000  26.500000 74.290000  26.570000 ;
        RECT 56.795000  26.570000 74.290000  26.640000 ;
        RECT 56.865000  26.640000 74.290000  26.710000 ;
        RECT 56.935000  26.710000 74.290000  26.780000 ;
        RECT 57.005000  26.780000 74.290000  26.850000 ;
        RECT 57.075000  26.850000 74.290000  26.920000 ;
        RECT 57.145000  26.920000 74.290000  26.990000 ;
        RECT 57.215000  26.990000 74.290000  27.060000 ;
        RECT 57.285000  27.060000 74.290000  27.130000 ;
        RECT 57.355000  27.130000 74.290000  27.200000 ;
        RECT 57.425000  27.200000 74.290000  27.270000 ;
        RECT 57.495000  27.270000 74.290000  27.340000 ;
        RECT 57.540000  47.390000 74.290000  47.455000 ;
        RECT 57.540000  70.420000 74.290000  70.455000 ;
        RECT 57.540000 116.390000 74.290000 116.455000 ;
        RECT 57.540000 139.425000 74.290000 139.455000 ;
        RECT 57.540000 162.440000 74.290000 162.455000 ;
        RECT 57.555000 148.155000 74.290000 148.225000 ;
        RECT 57.565000  27.340000 74.290000  27.410000 ;
        RECT 57.595000  56.155000 74.290000  56.225000 ;
        RECT 57.610000  47.320000 74.290000  47.390000 ;
        RECT 57.610000  70.350000 74.290000  70.420000 ;
        RECT 57.610000  93.410000 74.290000  93.455000 ;
        RECT 57.610000 116.320000 74.290000 116.390000 ;
        RECT 57.610000 139.355000 74.290000 139.425000 ;
        RECT 57.610000 162.370000 74.290000 162.440000 ;
        RECT 57.625000  79.155000 74.290000  79.225000 ;
        RECT 57.625000 102.155000 74.290000 102.225000 ;
        RECT 57.625000 125.155000 74.290000 125.225000 ;
        RECT 57.625000 148.225000 74.290000 148.295000 ;
        RECT 57.635000  27.410000 74.290000  27.480000 ;
        RECT 57.635000 171.155000 74.290000 171.225000 ;
        RECT 57.665000  56.225000 74.290000  56.295000 ;
        RECT 57.680000  47.250000 74.290000  47.320000 ;
        RECT 57.680000  70.280000 74.290000  70.350000 ;
        RECT 57.680000  93.340000 74.290000  93.410000 ;
        RECT 57.680000 116.250000 74.290000 116.320000 ;
        RECT 57.680000 139.285000 74.290000 139.355000 ;
        RECT 57.680000 162.300000 74.290000 162.370000 ;
        RECT 57.695000  79.225000 74.290000  79.295000 ;
        RECT 57.695000 102.225000 74.290000 102.295000 ;
        RECT 57.695000 125.225000 74.290000 125.295000 ;
        RECT 57.695000 148.295000 74.290000 148.365000 ;
        RECT 57.705000  27.480000 74.290000  27.550000 ;
        RECT 57.705000 171.225000 74.290000 171.295000 ;
        RECT 57.735000  56.295000 74.290000  56.365000 ;
        RECT 57.750000  47.180000 74.290000  47.250000 ;
        RECT 57.750000  70.210000 74.290000  70.280000 ;
        RECT 57.750000  93.270000 74.290000  93.340000 ;
        RECT 57.750000 116.180000 74.290000 116.250000 ;
        RECT 57.750000 139.215000 74.290000 139.285000 ;
        RECT 57.750000 162.230000 74.290000 162.300000 ;
        RECT 57.765000  79.295000 74.290000  79.365000 ;
        RECT 57.765000 102.295000 74.290000 102.365000 ;
        RECT 57.765000 125.295000 74.290000 125.365000 ;
        RECT 57.765000 148.365000 74.290000 148.435000 ;
        RECT 57.775000  27.550000 74.290000  27.620000 ;
        RECT 57.775000 171.295000 74.290000 171.365000 ;
        RECT 57.805000  56.365000 74.290000  56.435000 ;
        RECT 57.820000  47.110000 74.290000  47.180000 ;
        RECT 57.820000  70.140000 74.290000  70.210000 ;
        RECT 57.820000  93.200000 74.290000  93.270000 ;
        RECT 57.820000 116.110000 74.290000 116.180000 ;
        RECT 57.820000 139.145000 74.290000 139.215000 ;
        RECT 57.820000 162.160000 74.290000 162.230000 ;
        RECT 57.835000  79.365000 74.290000  79.435000 ;
        RECT 57.835000 102.365000 74.290000 102.435000 ;
        RECT 57.835000 125.365000 74.290000 125.435000 ;
        RECT 57.835000 148.435000 74.290000 148.505000 ;
        RECT 57.845000  27.620000 74.290000  27.690000 ;
        RECT 57.845000 171.365000 74.290000 171.435000 ;
        RECT 57.875000  56.435000 74.290000  56.505000 ;
        RECT 57.890000  47.040000 74.290000  47.110000 ;
        RECT 57.890000  70.070000 74.290000  70.140000 ;
        RECT 57.890000  93.130000 74.290000  93.200000 ;
        RECT 57.890000 116.040000 74.290000 116.110000 ;
        RECT 57.890000 139.075000 74.290000 139.145000 ;
        RECT 57.890000 162.090000 74.290000 162.160000 ;
        RECT 57.905000  79.435000 74.290000  79.505000 ;
        RECT 57.905000 102.435000 74.290000 102.505000 ;
        RECT 57.905000 125.435000 74.290000 125.505000 ;
        RECT 57.905000 148.505000 74.290000 148.575000 ;
        RECT 57.915000  27.690000 74.290000  27.760000 ;
        RECT 57.915000 171.435000 74.290000 171.505000 ;
        RECT 57.945000  56.505000 74.290000  56.575000 ;
        RECT 57.960000  46.970000 74.290000  47.040000 ;
        RECT 57.960000  70.000000 74.290000  70.070000 ;
        RECT 57.960000  93.060000 74.290000  93.130000 ;
        RECT 57.960000 115.970000 74.290000 116.040000 ;
        RECT 57.960000 139.005000 74.290000 139.075000 ;
        RECT 57.960000 162.020000 74.290000 162.090000 ;
        RECT 57.975000  79.505000 74.290000  79.575000 ;
        RECT 57.975000 102.505000 74.290000 102.575000 ;
        RECT 57.975000 125.505000 74.290000 125.575000 ;
        RECT 57.975000 148.575000 74.290000 148.645000 ;
        RECT 57.985000  27.760000 74.290000  27.830000 ;
        RECT 57.985000 171.505000 74.290000 171.575000 ;
        RECT 58.015000  56.575000 74.290000  56.645000 ;
        RECT 58.030000  46.900000 74.290000  46.970000 ;
        RECT 58.030000  69.930000 74.290000  70.000000 ;
        RECT 58.030000  92.990000 74.290000  93.060000 ;
        RECT 58.030000 115.900000 74.290000 115.970000 ;
        RECT 58.030000 138.935000 74.290000 139.005000 ;
        RECT 58.030000 161.950000 74.290000 162.020000 ;
        RECT 58.045000  79.575000 74.290000  79.645000 ;
        RECT 58.045000 102.575000 74.290000 102.645000 ;
        RECT 58.045000 125.575000 74.290000 125.645000 ;
        RECT 58.045000 148.645000 74.290000 148.715000 ;
        RECT 58.055000  27.830000 74.290000  27.900000 ;
        RECT 58.055000 171.575000 74.290000 171.645000 ;
        RECT 58.085000  56.645000 74.290000  56.715000 ;
        RECT 58.100000  46.830000 74.290000  46.900000 ;
        RECT 58.100000  69.860000 74.290000  69.930000 ;
        RECT 58.100000  92.920000 74.290000  92.990000 ;
        RECT 58.100000 115.830000 74.290000 115.900000 ;
        RECT 58.100000 138.865000 74.290000 138.935000 ;
        RECT 58.100000 161.880000 74.290000 161.950000 ;
        RECT 58.115000  79.645000 74.290000  79.715000 ;
        RECT 58.115000 102.645000 74.290000 102.715000 ;
        RECT 58.115000 125.645000 74.290000 125.715000 ;
        RECT 58.115000 148.715000 74.290000 148.785000 ;
        RECT 58.125000  27.900000 74.290000  27.970000 ;
        RECT 58.125000 171.645000 74.290000 171.715000 ;
        RECT 58.155000  56.715000 74.290000  56.785000 ;
        RECT 58.170000  46.760000 74.290000  46.830000 ;
        RECT 58.170000  69.790000 74.290000  69.860000 ;
        RECT 58.170000  92.850000 74.290000  92.920000 ;
        RECT 58.170000 115.760000 74.290000 115.830000 ;
        RECT 58.170000 138.795000 74.290000 138.865000 ;
        RECT 58.170000 161.810000 74.290000 161.880000 ;
        RECT 58.185000  79.715000 74.290000  79.785000 ;
        RECT 58.185000 102.715000 74.290000 102.785000 ;
        RECT 58.185000 125.715000 74.290000 125.785000 ;
        RECT 58.185000 148.785000 74.290000 148.855000 ;
        RECT 58.195000  27.970000 74.290000  28.040000 ;
        RECT 58.195000 171.715000 74.290000 171.785000 ;
        RECT 58.225000  56.785000 74.290000  56.855000 ;
        RECT 58.240000  46.690000 74.290000  46.760000 ;
        RECT 58.240000  69.720000 74.290000  69.790000 ;
        RECT 58.240000  92.780000 74.290000  92.850000 ;
        RECT 58.240000 115.690000 74.290000 115.760000 ;
        RECT 58.240000 138.725000 74.290000 138.795000 ;
        RECT 58.240000 161.740000 74.290000 161.810000 ;
        RECT 58.255000  79.785000 74.290000  79.855000 ;
        RECT 58.255000 102.785000 74.290000 102.855000 ;
        RECT 58.255000 125.785000 74.290000 125.855000 ;
        RECT 58.255000 148.855000 74.290000 148.925000 ;
        RECT 58.265000  28.040000 74.290000  28.110000 ;
        RECT 58.265000 171.785000 74.290000 171.855000 ;
        RECT 58.295000  56.855000 74.290000  56.925000 ;
        RECT 58.310000  46.620000 74.290000  46.690000 ;
        RECT 58.310000  69.650000 74.290000  69.720000 ;
        RECT 58.310000  92.710000 74.290000  92.780000 ;
        RECT 58.310000 115.620000 74.290000 115.690000 ;
        RECT 58.310000 138.655000 74.290000 138.725000 ;
        RECT 58.310000 161.670000 74.290000 161.740000 ;
        RECT 58.325000  79.855000 74.290000  79.925000 ;
        RECT 58.325000 102.855000 74.290000 102.925000 ;
        RECT 58.325000 125.855000 74.290000 125.925000 ;
        RECT 58.325000 148.925000 74.290000 148.995000 ;
        RECT 58.335000  28.110000 74.290000  28.180000 ;
        RECT 58.335000 171.855000 74.290000 171.925000 ;
        RECT 58.365000  56.925000 74.290000  56.995000 ;
        RECT 58.380000  46.550000 74.290000  46.620000 ;
        RECT 58.380000  69.580000 74.290000  69.650000 ;
        RECT 58.380000  92.640000 74.290000  92.710000 ;
        RECT 58.380000 115.550000 74.290000 115.620000 ;
        RECT 58.380000 138.585000 74.290000 138.655000 ;
        RECT 58.380000 161.600000 74.290000 161.670000 ;
        RECT 58.395000  79.925000 74.290000  79.995000 ;
        RECT 58.395000 102.925000 74.290000 102.995000 ;
        RECT 58.395000 125.925000 74.290000 125.995000 ;
        RECT 58.395000 148.995000 74.290000 149.065000 ;
        RECT 58.405000  28.180000 74.290000  28.250000 ;
        RECT 58.405000 171.925000 74.290000 171.995000 ;
        RECT 58.435000  56.995000 74.290000  57.065000 ;
        RECT 58.450000  46.480000 74.290000  46.550000 ;
        RECT 58.450000  69.510000 74.290000  69.580000 ;
        RECT 58.450000  92.570000 74.290000  92.640000 ;
        RECT 58.450000 115.480000 74.290000 115.550000 ;
        RECT 58.450000 138.515000 74.290000 138.585000 ;
        RECT 58.450000 161.530000 74.290000 161.600000 ;
        RECT 58.465000  79.995000 74.290000  80.065000 ;
        RECT 58.465000 102.995000 74.290000 103.065000 ;
        RECT 58.465000 125.995000 74.290000 126.065000 ;
        RECT 58.465000 149.065000 74.290000 149.135000 ;
        RECT 58.475000  28.250000 74.290000  28.320000 ;
        RECT 58.475000 171.995000 74.290000 172.065000 ;
        RECT 58.505000  57.065000 74.290000  57.135000 ;
        RECT 58.520000  46.410000 74.290000  46.480000 ;
        RECT 58.520000  69.440000 74.290000  69.510000 ;
        RECT 58.520000  92.500000 74.290000  92.570000 ;
        RECT 58.520000 115.410000 74.290000 115.480000 ;
        RECT 58.520000 138.445000 74.290000 138.515000 ;
        RECT 58.520000 161.460000 74.290000 161.530000 ;
        RECT 58.535000  80.065000 74.290000  80.135000 ;
        RECT 58.535000 103.065000 74.290000 103.135000 ;
        RECT 58.535000 126.065000 74.290000 126.135000 ;
        RECT 58.535000 149.135000 74.290000 149.205000 ;
        RECT 58.545000  28.320000 74.290000  28.390000 ;
        RECT 58.545000 172.065000 74.290000 172.135000 ;
        RECT 58.575000  57.135000 74.290000  57.205000 ;
        RECT 58.590000  46.340000 74.290000  46.410000 ;
        RECT 58.590000  69.370000 74.290000  69.440000 ;
        RECT 58.590000  92.430000 74.290000  92.500000 ;
        RECT 58.590000 115.340000 74.290000 115.410000 ;
        RECT 58.590000 138.375000 74.290000 138.445000 ;
        RECT 58.590000 161.390000 74.290000 161.460000 ;
        RECT 58.605000  80.135000 74.290000  80.205000 ;
        RECT 58.605000 103.135000 74.290000 103.205000 ;
        RECT 58.605000 126.135000 74.290000 126.205000 ;
        RECT 58.605000 149.205000 74.290000 149.275000 ;
        RECT 58.615000  28.390000 74.290000  28.460000 ;
        RECT 58.615000 172.135000 74.290000 172.205000 ;
        RECT 58.645000  57.205000 74.290000  57.275000 ;
        RECT 58.660000  46.270000 74.290000  46.340000 ;
        RECT 58.660000  69.300000 74.290000  69.370000 ;
        RECT 58.660000  92.360000 74.290000  92.430000 ;
        RECT 58.660000 115.270000 74.290000 115.340000 ;
        RECT 58.660000 138.305000 74.290000 138.375000 ;
        RECT 58.660000 161.320000 74.290000 161.390000 ;
        RECT 58.675000  80.205000 74.290000  80.275000 ;
        RECT 58.675000 103.205000 74.290000 103.275000 ;
        RECT 58.675000 126.205000 74.290000 126.275000 ;
        RECT 58.675000 149.275000 74.290000 149.345000 ;
        RECT 58.685000  28.460000 74.290000  28.530000 ;
        RECT 58.685000 172.205000 74.290000 172.275000 ;
        RECT 58.715000  57.275000 74.290000  57.345000 ;
        RECT 58.730000  46.200000 74.290000  46.270000 ;
        RECT 58.730000  69.230000 74.290000  69.300000 ;
        RECT 58.730000  92.290000 74.290000  92.360000 ;
        RECT 58.730000 115.200000 74.290000 115.270000 ;
        RECT 58.730000 138.235000 74.290000 138.305000 ;
        RECT 58.730000 161.250000 74.290000 161.320000 ;
        RECT 58.730000 185.260000 74.290000 185.295000 ;
        RECT 58.745000  80.275000 74.290000  80.345000 ;
        RECT 58.745000 103.275000 74.290000 103.345000 ;
        RECT 58.745000 126.275000 74.290000 126.345000 ;
        RECT 58.745000 149.345000 74.290000 149.415000 ;
        RECT 58.755000  28.530000 74.290000  28.600000 ;
        RECT 58.755000 172.275000 74.290000 172.345000 ;
        RECT 58.785000  57.345000 74.290000  57.415000 ;
        RECT 58.800000  46.130000 74.290000  46.200000 ;
        RECT 58.800000  69.160000 74.290000  69.230000 ;
        RECT 58.800000  92.220000 74.290000  92.290000 ;
        RECT 58.800000 115.130000 74.290000 115.200000 ;
        RECT 58.800000 138.165000 74.290000 138.235000 ;
        RECT 58.800000 161.180000 74.290000 161.250000 ;
        RECT 58.800000 185.190000 74.290000 185.260000 ;
        RECT 58.815000  80.345000 74.290000  80.415000 ;
        RECT 58.815000 103.345000 74.290000 103.415000 ;
        RECT 58.815000 126.345000 74.290000 126.415000 ;
        RECT 58.815000 149.415000 74.290000 149.485000 ;
        RECT 58.825000  28.600000 74.290000  28.670000 ;
        RECT 58.825000 172.345000 74.290000 172.415000 ;
        RECT 58.855000  57.415000 74.290000  57.485000 ;
        RECT 58.870000  46.060000 74.290000  46.130000 ;
        RECT 58.870000  69.090000 74.290000  69.160000 ;
        RECT 58.870000  92.150000 74.290000  92.220000 ;
        RECT 58.870000 115.060000 74.290000 115.130000 ;
        RECT 58.870000 138.095000 74.290000 138.165000 ;
        RECT 58.870000 161.110000 74.290000 161.180000 ;
        RECT 58.870000 185.120000 74.290000 185.190000 ;
        RECT 58.885000  80.415000 74.290000  80.485000 ;
        RECT 58.885000 103.415000 74.290000 103.485000 ;
        RECT 58.885000 126.415000 74.290000 126.485000 ;
        RECT 58.885000 149.485000 74.290000 149.555000 ;
        RECT 58.895000  28.670000 74.290000  28.740000 ;
        RECT 58.895000 172.415000 74.290000 172.485000 ;
        RECT 58.925000  57.485000 74.290000  57.555000 ;
        RECT 58.940000  45.990000 74.290000  46.060000 ;
        RECT 58.940000  69.020000 74.290000  69.090000 ;
        RECT 58.940000  92.080000 74.290000  92.150000 ;
        RECT 58.940000 114.990000 74.290000 115.060000 ;
        RECT 58.940000 138.025000 74.290000 138.095000 ;
        RECT 58.940000 161.040000 74.290000 161.110000 ;
        RECT 58.940000 185.050000 74.290000 185.120000 ;
        RECT 58.955000  80.485000 74.290000  80.555000 ;
        RECT 58.955000 103.485000 74.290000 103.555000 ;
        RECT 58.955000 126.485000 74.290000 126.555000 ;
        RECT 58.955000 149.555000 74.290000 149.625000 ;
        RECT 58.965000  28.740000 74.290000  28.810000 ;
        RECT 58.965000 172.485000 74.290000 172.555000 ;
        RECT 58.995000  57.555000 74.290000  57.625000 ;
        RECT 59.010000  45.920000 74.290000  45.990000 ;
        RECT 59.010000  68.950000 74.290000  69.020000 ;
        RECT 59.010000  92.010000 74.290000  92.080000 ;
        RECT 59.010000 114.920000 74.290000 114.990000 ;
        RECT 59.010000 137.955000 74.290000 138.025000 ;
        RECT 59.010000 160.970000 74.290000 161.040000 ;
        RECT 59.010000 184.980000 74.290000 185.050000 ;
        RECT 59.025000  80.555000 74.290000  80.625000 ;
        RECT 59.025000 103.555000 74.290000 103.625000 ;
        RECT 59.025000 126.555000 74.290000 126.625000 ;
        RECT 59.025000 149.625000 74.290000 149.695000 ;
        RECT 59.035000  28.810000 74.290000  28.880000 ;
        RECT 59.035000 172.555000 74.290000 172.625000 ;
        RECT 59.065000  57.625000 74.290000  57.695000 ;
        RECT 59.080000  45.850000 74.290000  45.920000 ;
        RECT 59.080000  68.880000 74.290000  68.950000 ;
        RECT 59.080000  91.940000 74.290000  92.010000 ;
        RECT 59.080000 114.850000 74.290000 114.920000 ;
        RECT 59.080000 137.885000 74.290000 137.955000 ;
        RECT 59.080000 160.900000 74.290000 160.970000 ;
        RECT 59.080000 184.910000 74.290000 184.980000 ;
        RECT 59.095000  80.625000 74.290000  80.695000 ;
        RECT 59.095000 103.625000 74.290000 103.695000 ;
        RECT 59.095000 126.625000 74.290000 126.695000 ;
        RECT 59.095000 149.695000 74.290000 149.765000 ;
        RECT 59.105000  28.880000 74.290000  28.950000 ;
        RECT 59.105000 172.625000 74.290000 172.695000 ;
        RECT 59.135000  57.695000 74.290000  57.765000 ;
        RECT 59.150000  45.780000 74.290000  45.850000 ;
        RECT 59.150000  68.810000 74.290000  68.880000 ;
        RECT 59.150000  91.870000 74.290000  91.940000 ;
        RECT 59.150000 114.780000 74.290000 114.850000 ;
        RECT 59.150000 137.815000 74.290000 137.885000 ;
        RECT 59.150000 160.830000 74.290000 160.900000 ;
        RECT 59.150000 184.840000 74.290000 184.910000 ;
        RECT 59.165000  80.695000 74.290000  80.765000 ;
        RECT 59.165000 103.695000 74.290000 103.765000 ;
        RECT 59.165000 126.695000 74.290000 126.765000 ;
        RECT 59.165000 149.765000 74.290000 149.835000 ;
        RECT 59.175000  28.950000 74.290000  29.020000 ;
        RECT 59.175000 172.695000 74.290000 172.765000 ;
        RECT 59.205000  57.765000 74.290000  57.835000 ;
        RECT 59.220000  45.710000 74.290000  45.780000 ;
        RECT 59.220000  68.740000 74.290000  68.810000 ;
        RECT 59.220000  91.800000 74.290000  91.870000 ;
        RECT 59.220000 114.710000 74.290000 114.780000 ;
        RECT 59.220000 137.745000 74.290000 137.815000 ;
        RECT 59.220000 160.760000 74.290000 160.830000 ;
        RECT 59.220000 184.770000 74.290000 184.840000 ;
        RECT 59.235000  80.765000 74.290000  80.835000 ;
        RECT 59.235000 103.765000 74.290000 103.835000 ;
        RECT 59.235000 126.765000 74.290000 126.835000 ;
        RECT 59.235000 149.835000 74.290000 149.905000 ;
        RECT 59.245000  29.020000 74.290000  29.090000 ;
        RECT 59.245000 172.765000 74.290000 172.835000 ;
        RECT 59.275000  57.835000 74.290000  57.905000 ;
        RECT 59.290000  45.640000 74.290000  45.710000 ;
        RECT 59.290000  68.670000 74.290000  68.740000 ;
        RECT 59.290000  91.730000 74.290000  91.800000 ;
        RECT 59.290000 114.640000 74.290000 114.710000 ;
        RECT 59.290000 137.675000 74.290000 137.745000 ;
        RECT 59.290000 160.690000 74.290000 160.760000 ;
        RECT 59.290000 184.700000 74.290000 184.770000 ;
        RECT 59.305000  80.835000 74.290000  80.905000 ;
        RECT 59.305000 103.835000 74.290000 103.905000 ;
        RECT 59.305000 126.835000 74.290000 126.905000 ;
        RECT 59.305000 149.905000 74.290000 149.975000 ;
        RECT 59.315000  29.090000 74.290000  29.160000 ;
        RECT 59.315000 172.835000 74.290000 172.905000 ;
        RECT 59.345000  57.905000 74.290000  57.975000 ;
        RECT 59.360000  45.570000 74.290000  45.640000 ;
        RECT 59.360000  68.600000 74.290000  68.670000 ;
        RECT 59.360000  91.660000 74.290000  91.730000 ;
        RECT 59.360000 114.570000 74.290000 114.640000 ;
        RECT 59.360000 137.605000 74.290000 137.675000 ;
        RECT 59.360000 160.620000 74.290000 160.690000 ;
        RECT 59.360000 184.630000 74.290000 184.700000 ;
        RECT 59.375000  80.905000 74.290000  80.975000 ;
        RECT 59.375000 103.905000 74.290000 103.975000 ;
        RECT 59.375000 126.905000 74.290000 126.975000 ;
        RECT 59.375000 149.975000 74.290000 150.045000 ;
        RECT 59.385000  29.160000 74.290000  29.230000 ;
        RECT 59.385000 172.905000 74.290000 172.975000 ;
        RECT 59.415000  57.975000 74.290000  58.045000 ;
        RECT 59.430000  45.500000 74.290000  45.570000 ;
        RECT 59.430000  68.530000 74.290000  68.600000 ;
        RECT 59.430000  91.590000 74.290000  91.660000 ;
        RECT 59.430000 114.500000 74.290000 114.570000 ;
        RECT 59.430000 137.535000 74.290000 137.605000 ;
        RECT 59.430000 160.550000 74.290000 160.620000 ;
        RECT 59.430000 184.560000 74.290000 184.630000 ;
        RECT 59.445000  80.975000 74.290000  81.045000 ;
        RECT 59.445000 103.975000 74.290000 104.045000 ;
        RECT 59.445000 126.975000 74.290000 127.045000 ;
        RECT 59.445000 150.045000 74.290000 150.115000 ;
        RECT 59.455000  29.230000 74.290000  29.300000 ;
        RECT 59.455000 172.975000 74.290000 173.045000 ;
        RECT 59.485000  58.045000 74.290000  58.115000 ;
        RECT 59.500000  45.430000 74.290000  45.500000 ;
        RECT 59.500000  68.460000 74.290000  68.530000 ;
        RECT 59.500000  91.520000 74.290000  91.590000 ;
        RECT 59.500000 114.430000 74.290000 114.500000 ;
        RECT 59.500000 137.465000 74.290000 137.535000 ;
        RECT 59.500000 160.480000 74.290000 160.550000 ;
        RECT 59.500000 184.490000 74.290000 184.560000 ;
        RECT 59.515000  81.045000 74.290000  81.115000 ;
        RECT 59.515000 104.045000 74.290000 104.115000 ;
        RECT 59.515000 127.045000 74.290000 127.115000 ;
        RECT 59.515000 150.115000 74.290000 150.185000 ;
        RECT 59.525000  29.300000 74.290000  29.370000 ;
        RECT 59.525000 173.045000 74.290000 173.115000 ;
        RECT 59.555000  58.115000 74.290000  58.185000 ;
        RECT 59.570000  45.360000 74.290000  45.430000 ;
        RECT 59.570000  68.390000 74.290000  68.460000 ;
        RECT 59.570000  91.450000 74.290000  91.520000 ;
        RECT 59.570000 114.360000 74.290000 114.430000 ;
        RECT 59.570000 137.395000 74.290000 137.465000 ;
        RECT 59.570000 160.410000 74.290000 160.480000 ;
        RECT 59.570000 184.420000 74.290000 184.490000 ;
        RECT 59.585000  81.115000 74.290000  81.185000 ;
        RECT 59.585000 104.115000 74.290000 104.185000 ;
        RECT 59.585000 127.115000 74.290000 127.185000 ;
        RECT 59.585000 150.185000 74.290000 150.255000 ;
        RECT 59.595000  29.370000 74.290000  29.440000 ;
        RECT 59.595000 173.115000 74.290000 173.185000 ;
        RECT 59.625000  58.185000 74.290000  58.255000 ;
        RECT 59.640000  45.290000 74.290000  45.360000 ;
        RECT 59.640000  68.320000 74.290000  68.390000 ;
        RECT 59.640000  91.380000 74.290000  91.450000 ;
        RECT 59.640000 114.290000 74.290000 114.360000 ;
        RECT 59.640000 137.325000 74.290000 137.395000 ;
        RECT 59.640000 160.340000 74.290000 160.410000 ;
        RECT 59.640000 184.350000 74.290000 184.420000 ;
        RECT 59.655000  81.185000 74.290000  81.255000 ;
        RECT 59.655000 104.185000 74.290000 104.255000 ;
        RECT 59.655000 127.185000 74.290000 127.255000 ;
        RECT 59.655000 150.255000 74.290000 150.325000 ;
        RECT 59.665000  29.440000 74.290000  29.510000 ;
        RECT 59.665000 173.185000 74.290000 173.255000 ;
        RECT 59.695000  58.255000 74.290000  58.325000 ;
        RECT 59.710000  45.220000 74.290000  45.290000 ;
        RECT 59.710000  68.250000 74.290000  68.320000 ;
        RECT 59.710000  91.310000 74.290000  91.380000 ;
        RECT 59.710000 114.220000 74.290000 114.290000 ;
        RECT 59.710000 137.255000 74.290000 137.325000 ;
        RECT 59.710000 160.270000 74.290000 160.340000 ;
        RECT 59.710000 184.280000 74.290000 184.350000 ;
        RECT 59.725000  81.255000 74.290000  81.325000 ;
        RECT 59.725000 104.255000 74.290000 104.325000 ;
        RECT 59.725000 127.255000 74.290000 127.325000 ;
        RECT 59.725000 150.325000 74.290000 150.395000 ;
        RECT 59.735000  29.510000 74.290000  29.580000 ;
        RECT 59.735000 173.255000 74.290000 173.325000 ;
        RECT 59.765000  58.325000 74.290000  58.395000 ;
        RECT 59.780000  45.150000 74.290000  45.220000 ;
        RECT 59.780000  68.180000 74.290000  68.250000 ;
        RECT 59.780000  91.240000 74.290000  91.310000 ;
        RECT 59.780000 114.150000 74.290000 114.220000 ;
        RECT 59.780000 137.185000 74.290000 137.255000 ;
        RECT 59.780000 160.200000 74.290000 160.270000 ;
        RECT 59.780000 184.210000 74.290000 184.280000 ;
        RECT 59.795000  81.325000 74.290000  81.395000 ;
        RECT 59.795000 104.325000 74.290000 104.395000 ;
        RECT 59.795000 127.325000 74.290000 127.395000 ;
        RECT 59.795000 150.395000 74.290000 150.465000 ;
        RECT 59.805000  29.580000 74.290000  29.650000 ;
        RECT 59.805000 173.325000 74.290000 173.395000 ;
        RECT 59.835000  58.395000 74.290000  58.465000 ;
        RECT 59.850000  45.080000 74.290000  45.150000 ;
        RECT 59.850000  68.110000 74.290000  68.180000 ;
        RECT 59.850000  91.170000 74.290000  91.240000 ;
        RECT 59.850000 114.080000 74.290000 114.150000 ;
        RECT 59.850000 137.115000 74.290000 137.185000 ;
        RECT 59.850000 160.130000 74.290000 160.200000 ;
        RECT 59.850000 184.140000 74.290000 184.210000 ;
        RECT 59.865000  81.395000 74.290000  81.465000 ;
        RECT 59.865000 104.395000 74.290000 104.465000 ;
        RECT 59.865000 127.395000 74.290000 127.465000 ;
        RECT 59.865000 150.465000 74.290000 150.535000 ;
        RECT 59.875000  29.650000 74.290000  29.720000 ;
        RECT 59.875000 173.395000 74.290000 173.465000 ;
        RECT 59.905000  58.465000 74.290000  58.535000 ;
        RECT 59.920000  45.010000 74.290000  45.080000 ;
        RECT 59.920000  68.040000 74.290000  68.110000 ;
        RECT 59.920000  91.100000 74.290000  91.170000 ;
        RECT 59.920000 114.010000 74.290000 114.080000 ;
        RECT 59.920000 137.045000 74.290000 137.115000 ;
        RECT 59.920000 160.060000 74.290000 160.130000 ;
        RECT 59.920000 184.070000 74.290000 184.140000 ;
        RECT 59.935000  81.465000 74.290000  81.535000 ;
        RECT 59.935000 104.465000 74.290000 104.535000 ;
        RECT 59.935000 127.465000 74.290000 127.535000 ;
        RECT 59.935000 150.535000 74.290000 150.605000 ;
        RECT 59.945000  29.720000 74.290000  29.790000 ;
        RECT 59.945000 173.465000 74.290000 173.535000 ;
        RECT 59.975000  58.535000 74.290000  58.605000 ;
        RECT 59.990000  44.940000 74.290000  45.010000 ;
        RECT 59.990000  67.970000 74.290000  68.040000 ;
        RECT 59.990000  91.030000 74.290000  91.100000 ;
        RECT 59.990000 113.940000 74.290000 114.010000 ;
        RECT 59.990000 136.975000 74.290000 137.045000 ;
        RECT 59.990000 159.990000 74.290000 160.060000 ;
        RECT 59.990000 184.000000 74.290000 184.070000 ;
        RECT 60.005000  81.535000 74.290000  81.605000 ;
        RECT 60.005000 104.535000 74.290000 104.605000 ;
        RECT 60.005000 127.535000 74.290000 127.605000 ;
        RECT 60.005000 150.605000 74.290000 150.675000 ;
        RECT 60.015000  29.790000 74.290000  29.860000 ;
        RECT 60.015000 173.535000 74.290000 173.605000 ;
        RECT 60.045000  58.605000 74.290000  58.675000 ;
        RECT 60.060000  44.870000 74.290000  44.940000 ;
        RECT 60.060000  67.900000 74.290000  67.970000 ;
        RECT 60.060000  90.960000 74.290000  91.030000 ;
        RECT 60.060000 113.870000 74.290000 113.940000 ;
        RECT 60.060000 136.905000 74.290000 136.975000 ;
        RECT 60.060000 159.920000 74.290000 159.990000 ;
        RECT 60.060000 183.930000 74.290000 184.000000 ;
        RECT 60.075000  81.605000 74.290000  81.675000 ;
        RECT 60.075000 104.605000 74.290000 104.675000 ;
        RECT 60.075000 127.605000 74.290000 127.675000 ;
        RECT 60.075000 150.675000 74.290000 150.745000 ;
        RECT 60.085000  29.860000 74.290000  29.930000 ;
        RECT 60.085000 173.605000 74.290000 173.675000 ;
        RECT 60.115000  58.675000 74.290000  58.745000 ;
        RECT 60.130000  44.800000 74.290000  44.870000 ;
        RECT 60.130000  67.830000 74.290000  67.900000 ;
        RECT 60.130000  90.890000 74.290000  90.960000 ;
        RECT 60.130000 113.800000 74.290000 113.870000 ;
        RECT 60.130000 136.835000 74.290000 136.905000 ;
        RECT 60.130000 159.850000 74.290000 159.920000 ;
        RECT 60.130000 183.860000 74.290000 183.930000 ;
        RECT 60.145000  81.675000 74.290000  81.745000 ;
        RECT 60.145000 104.675000 74.290000 104.745000 ;
        RECT 60.145000 127.675000 74.290000 127.745000 ;
        RECT 60.145000 150.745000 74.290000 150.815000 ;
        RECT 60.155000  29.930000 74.290000  30.000000 ;
        RECT 60.155000 173.675000 74.290000 173.745000 ;
        RECT 60.185000  58.745000 74.290000  58.815000 ;
        RECT 60.200000  44.730000 74.290000  44.800000 ;
        RECT 60.200000  67.760000 74.290000  67.830000 ;
        RECT 60.200000  90.820000 74.290000  90.890000 ;
        RECT 60.200000 113.730000 74.290000 113.800000 ;
        RECT 60.200000 136.765000 74.290000 136.835000 ;
        RECT 60.200000 159.780000 74.290000 159.850000 ;
        RECT 60.200000 183.790000 74.290000 183.860000 ;
        RECT 60.215000  81.745000 74.290000  81.815000 ;
        RECT 60.215000 104.745000 74.290000 104.815000 ;
        RECT 60.215000 127.745000 74.290000 127.815000 ;
        RECT 60.215000 150.815000 74.290000 150.885000 ;
        RECT 60.225000  30.000000 74.290000  30.070000 ;
        RECT 60.225000 173.745000 74.290000 173.815000 ;
        RECT 60.255000  58.815000 74.290000  58.885000 ;
        RECT 60.270000  44.660000 74.290000  44.730000 ;
        RECT 60.270000  67.690000 74.290000  67.760000 ;
        RECT 60.270000  90.750000 74.290000  90.820000 ;
        RECT 60.270000 113.660000 74.290000 113.730000 ;
        RECT 60.270000 136.695000 74.290000 136.765000 ;
        RECT 60.270000 159.710000 74.290000 159.780000 ;
        RECT 60.270000 183.720000 74.290000 183.790000 ;
        RECT 60.285000  81.815000 74.290000  81.885000 ;
        RECT 60.285000 104.815000 74.290000 104.885000 ;
        RECT 60.285000 127.815000 74.290000 127.885000 ;
        RECT 60.285000 150.885000 74.290000 150.955000 ;
        RECT 60.295000  30.070000 74.290000  30.140000 ;
        RECT 60.295000 173.815000 74.290000 173.885000 ;
        RECT 60.325000  58.885000 74.290000  58.955000 ;
        RECT 60.340000  44.590000 74.290000  44.660000 ;
        RECT 60.340000  67.620000 74.290000  67.690000 ;
        RECT 60.340000  90.680000 74.290000  90.750000 ;
        RECT 60.340000 113.590000 74.290000 113.660000 ;
        RECT 60.340000 136.625000 74.290000 136.695000 ;
        RECT 60.340000 159.640000 74.290000 159.710000 ;
        RECT 60.340000 183.650000 74.290000 183.720000 ;
        RECT 60.355000  81.885000 74.290000  81.955000 ;
        RECT 60.355000 104.885000 74.290000 104.955000 ;
        RECT 60.355000 127.885000 74.290000 127.955000 ;
        RECT 60.355000 150.955000 74.290000 151.025000 ;
        RECT 60.365000  30.140000 74.290000  30.210000 ;
        RECT 60.365000 173.885000 74.290000 173.955000 ;
        RECT 60.395000  58.955000 74.290000  59.025000 ;
        RECT 60.410000  44.520000 74.290000  44.590000 ;
        RECT 60.410000  67.550000 74.290000  67.620000 ;
        RECT 60.410000  90.610000 74.290000  90.680000 ;
        RECT 60.410000 113.520000 74.290000 113.590000 ;
        RECT 60.410000 136.555000 74.290000 136.625000 ;
        RECT 60.410000 159.570000 74.290000 159.640000 ;
        RECT 60.410000 183.580000 74.290000 183.650000 ;
        RECT 60.425000  81.955000 74.290000  82.025000 ;
        RECT 60.425000 104.955000 74.290000 105.025000 ;
        RECT 60.425000 127.955000 74.290000 128.025000 ;
        RECT 60.425000 151.025000 74.290000 151.095000 ;
        RECT 60.435000  30.210000 74.290000  30.280000 ;
        RECT 60.435000 173.955000 74.290000 174.025000 ;
        RECT 60.465000  59.025000 74.290000  59.095000 ;
        RECT 60.480000  44.450000 74.290000  44.520000 ;
        RECT 60.480000  67.480000 74.290000  67.550000 ;
        RECT 60.480000  90.540000 74.290000  90.610000 ;
        RECT 60.480000 113.450000 74.290000 113.520000 ;
        RECT 60.480000 136.485000 74.290000 136.555000 ;
        RECT 60.480000 159.500000 74.290000 159.570000 ;
        RECT 60.480000 183.510000 74.290000 183.580000 ;
        RECT 60.495000  82.025000 74.290000  82.095000 ;
        RECT 60.495000 105.025000 74.290000 105.095000 ;
        RECT 60.495000 128.025000 74.290000 128.095000 ;
        RECT 60.495000 151.095000 74.290000 151.165000 ;
        RECT 60.505000  30.280000 74.290000  30.350000 ;
        RECT 60.505000 174.025000 74.290000 174.095000 ;
        RECT 60.535000  59.095000 74.290000  59.165000 ;
        RECT 60.550000  44.380000 74.290000  44.450000 ;
        RECT 60.550000  67.410000 74.290000  67.480000 ;
        RECT 60.550000  90.470000 74.290000  90.540000 ;
        RECT 60.550000 113.380000 74.290000 113.450000 ;
        RECT 60.550000 136.415000 74.290000 136.485000 ;
        RECT 60.550000 159.430000 74.290000 159.500000 ;
        RECT 60.550000 183.440000 74.290000 183.510000 ;
        RECT 60.565000  82.095000 74.290000  82.165000 ;
        RECT 60.565000 105.095000 74.290000 105.165000 ;
        RECT 60.565000 128.095000 74.290000 128.165000 ;
        RECT 60.565000 151.165000 74.290000 151.235000 ;
        RECT 60.575000  30.350000 74.290000  30.420000 ;
        RECT 60.575000 174.095000 74.290000 174.165000 ;
        RECT 60.605000  59.165000 74.290000  59.235000 ;
        RECT 60.620000  44.310000 74.290000  44.380000 ;
        RECT 60.620000  67.340000 74.290000  67.410000 ;
        RECT 60.620000  90.400000 74.290000  90.470000 ;
        RECT 60.620000 113.310000 74.290000 113.380000 ;
        RECT 60.620000 136.345000 74.290000 136.415000 ;
        RECT 60.620000 159.360000 74.290000 159.430000 ;
        RECT 60.620000 183.370000 74.290000 183.440000 ;
        RECT 60.635000  82.165000 74.290000  82.235000 ;
        RECT 60.635000 105.165000 74.290000 105.235000 ;
        RECT 60.635000 128.165000 74.290000 128.235000 ;
        RECT 60.635000 151.235000 74.290000 151.305000 ;
        RECT 60.645000  30.420000 74.290000  30.490000 ;
        RECT 60.645000 174.165000 74.290000 174.235000 ;
        RECT 60.675000  59.235000 74.290000  59.305000 ;
        RECT 60.690000  44.240000 74.290000  44.310000 ;
        RECT 60.690000  67.270000 74.290000  67.340000 ;
        RECT 60.690000  90.330000 74.290000  90.400000 ;
        RECT 60.690000 113.240000 74.290000 113.310000 ;
        RECT 60.690000 136.275000 74.290000 136.345000 ;
        RECT 60.690000 159.290000 74.290000 159.360000 ;
        RECT 60.690000 183.300000 74.290000 183.370000 ;
        RECT 60.705000  82.235000 74.290000  82.305000 ;
        RECT 60.705000 105.235000 74.290000 105.305000 ;
        RECT 60.705000 128.235000 74.290000 128.305000 ;
        RECT 60.705000 151.305000 74.290000 151.375000 ;
        RECT 60.715000  30.490000 74.290000  30.560000 ;
        RECT 60.715000 174.235000 74.290000 174.305000 ;
        RECT 60.745000  59.305000 74.290000  59.375000 ;
        RECT 60.760000  44.170000 74.290000  44.240000 ;
        RECT 60.760000  67.200000 74.290000  67.270000 ;
        RECT 60.760000  90.260000 74.290000  90.330000 ;
        RECT 60.760000 113.170000 74.290000 113.240000 ;
        RECT 60.760000 136.205000 74.290000 136.275000 ;
        RECT 60.760000 159.220000 74.290000 159.290000 ;
        RECT 60.760000 183.230000 74.290000 183.300000 ;
        RECT 60.775000  82.305000 74.290000  82.375000 ;
        RECT 60.775000 105.305000 74.290000 105.375000 ;
        RECT 60.775000 128.305000 74.290000 128.375000 ;
        RECT 60.775000 151.375000 74.290000 151.445000 ;
        RECT 60.785000  30.560000 74.290000  30.630000 ;
        RECT 60.785000 174.305000 74.290000 174.375000 ;
        RECT 60.815000  59.375000 74.290000  59.445000 ;
        RECT 60.830000  44.100000 74.290000  44.170000 ;
        RECT 60.830000  67.130000 74.290000  67.200000 ;
        RECT 60.830000  90.190000 74.290000  90.260000 ;
        RECT 60.830000 113.100000 74.290000 113.170000 ;
        RECT 60.830000 136.135000 74.290000 136.205000 ;
        RECT 60.830000 159.150000 74.290000 159.220000 ;
        RECT 60.830000 183.160000 74.290000 183.230000 ;
        RECT 60.845000  82.375000 74.290000  82.445000 ;
        RECT 60.845000 105.375000 74.290000 105.445000 ;
        RECT 60.845000 128.375000 74.290000 128.445000 ;
        RECT 60.845000 151.445000 74.290000 151.515000 ;
        RECT 60.855000  30.630000 74.290000  30.700000 ;
        RECT 60.855000 174.375000 74.290000 174.445000 ;
        RECT 60.885000  59.445000 74.290000  59.515000 ;
        RECT 60.900000  44.030000 74.290000  44.100000 ;
        RECT 60.900000  67.060000 74.290000  67.130000 ;
        RECT 60.900000  90.120000 74.290000  90.190000 ;
        RECT 60.900000 113.030000 74.290000 113.100000 ;
        RECT 60.900000 136.065000 74.290000 136.135000 ;
        RECT 60.900000 159.080000 74.290000 159.150000 ;
        RECT 60.900000 183.090000 74.290000 183.160000 ;
        RECT 60.915000  82.445000 74.290000  82.515000 ;
        RECT 60.915000 105.445000 74.290000 105.515000 ;
        RECT 60.915000 128.445000 74.290000 128.515000 ;
        RECT 60.915000 151.515000 74.290000 151.585000 ;
        RECT 60.925000  30.700000 74.290000  30.770000 ;
        RECT 60.925000 174.445000 74.290000 174.515000 ;
        RECT 60.955000  59.515000 74.290000  59.585000 ;
        RECT 60.970000  43.960000 74.290000  44.030000 ;
        RECT 60.970000  66.990000 74.290000  67.060000 ;
        RECT 60.970000  90.050000 74.290000  90.120000 ;
        RECT 60.970000 112.960000 74.290000 113.030000 ;
        RECT 60.970000 135.995000 74.290000 136.065000 ;
        RECT 60.970000 159.010000 74.290000 159.080000 ;
        RECT 60.970000 183.020000 74.290000 183.090000 ;
        RECT 60.985000  82.515000 74.290000  82.585000 ;
        RECT 60.985000 105.515000 74.290000 105.585000 ;
        RECT 60.985000 128.515000 74.290000 128.585000 ;
        RECT 60.985000 151.585000 74.290000 151.655000 ;
        RECT 60.995000  30.770000 74.290000  30.840000 ;
        RECT 60.995000 174.515000 74.290000 174.585000 ;
        RECT 61.025000  59.585000 74.290000  59.655000 ;
        RECT 61.040000  43.890000 74.290000  43.960000 ;
        RECT 61.040000  66.920000 74.290000  66.990000 ;
        RECT 61.040000  89.980000 74.290000  90.050000 ;
        RECT 61.040000 112.890000 74.290000 112.960000 ;
        RECT 61.040000 135.925000 74.290000 135.995000 ;
        RECT 61.040000 158.940000 74.290000 159.010000 ;
        RECT 61.040000 182.950000 74.290000 183.020000 ;
        RECT 61.055000  82.585000 74.290000  82.655000 ;
        RECT 61.055000 105.585000 74.290000 105.655000 ;
        RECT 61.055000 128.585000 74.290000 128.655000 ;
        RECT 61.055000 151.655000 74.290000 151.725000 ;
        RECT 61.065000  30.840000 74.290000  30.910000 ;
        RECT 61.065000 174.585000 74.290000 174.655000 ;
        RECT 61.095000  59.655000 74.290000  59.725000 ;
        RECT 61.110000  30.910000 74.290000  30.955000 ;
        RECT 61.110000  30.955000 74.290000  43.820000 ;
        RECT 61.110000  43.820000 74.290000  43.890000 ;
        RECT 61.110000  59.725000 74.290000  59.740000 ;
        RECT 61.110000  59.740000 74.290000  66.850000 ;
        RECT 61.110000  66.850000 74.290000  66.920000 ;
        RECT 61.110000  82.655000 74.290000  82.710000 ;
        RECT 61.110000  82.710000 74.290000  89.910000 ;
        RECT 61.110000  89.910000 74.290000  89.980000 ;
        RECT 61.110000 105.655000 74.290000 105.710000 ;
        RECT 61.110000 105.710000 74.290000 112.820000 ;
        RECT 61.110000 112.820000 74.290000 112.890000 ;
        RECT 61.110000 128.655000 74.290000 128.710000 ;
        RECT 61.110000 128.710000 74.290000 135.855000 ;
        RECT 61.110000 135.855000 74.290000 135.925000 ;
        RECT 61.110000 151.725000 74.290000 151.780000 ;
        RECT 61.110000 151.780000 74.290000 158.870000 ;
        RECT 61.110000 158.870000 74.290000 158.940000 ;
        RECT 61.110000 174.655000 74.290000 174.700000 ;
        RECT 61.110000 174.700000 74.290000 182.880000 ;
        RECT 61.110000 182.880000 74.290000 182.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000   0.000000 48.890000  96.150000 ;
        RECT 37.890000  96.150000 48.890000  96.300000 ;
        RECT 37.890000  96.300000 49.040000  96.450000 ;
        RECT 37.890000  96.450000 49.190000  96.600000 ;
        RECT 37.890000  96.600000 49.340000  96.750000 ;
        RECT 37.890000  96.750000 49.490000  96.900000 ;
        RECT 37.890000  96.900000 49.640000  97.050000 ;
        RECT 37.890000  97.050000 49.790000  97.200000 ;
        RECT 37.890000  97.200000 49.940000  97.350000 ;
        RECT 37.890000  97.350000 50.090000  97.500000 ;
        RECT 37.890000  97.500000 50.240000  97.650000 ;
        RECT 37.890000  97.650000 50.390000  97.800000 ;
        RECT 37.890000  97.800000 50.540000  97.950000 ;
        RECT 37.890000  97.950000 50.690000  98.100000 ;
        RECT 37.890000  98.100000 50.840000  98.250000 ;
        RECT 37.890000  98.250000 50.990000  98.300000 ;
        RECT 37.890000  98.300000 51.040000  99.505000 ;
        RECT 37.890000  99.505000 43.400000  99.655000 ;
        RECT 37.890000  99.655000 43.250000  99.805000 ;
        RECT 37.890000  99.805000 43.100000  99.955000 ;
        RECT 37.890000  99.955000 42.950000 100.105000 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
        RECT 37.890000 104.385000 45.090000 104.535000 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
        RECT 38.340000 105.955000 46.660000 106.105000 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
        RECT 40.385000 108.055000 48.760000 108.150000 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
        RECT 42.705000 170.610000 48.855000 170.760000 ;
        RECT 42.785000 110.400000 48.855000 110.550000 ;
        RECT 42.855000 110.550000 48.855000 110.620000 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
        RECT 44.655000  99.505000 51.040000  99.610000 ;
        RECT 44.760000  99.610000 51.040000  99.715000 ;
        RECT 44.910000  99.715000 51.040000  99.865000 ;
        RECT 45.060000  99.865000 51.190000 100.015000 ;
        RECT 45.210000 100.015000 51.340000 100.165000 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
        RECT 47.360000 104.365000 55.690000 104.515000 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
        RECT 48.710000 105.715000 57.040000 105.865000 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
        RECT 49.775000 173.020000 59.285000 173.170000 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
        RECT 49.775000 174.670000 60.935000 174.680000 ;
        RECT 49.775000 174.680000 60.945000 190.040000 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
        RECT 50.805000 107.815000 59.140000 107.960000 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
        RECT 50.955000 107.960000 59.285000 108.110000 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
        RECT 53.135000 169.285000 59.285000 169.435000 ;
        RECT 53.205000 110.210000 59.285000 110.360000 ;
        RECT 53.285000 110.360000 59.285000 110.440000 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
  END DRN_HVC
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000   0.000000 24.395000  36.510000 ;
        RECT 0.495000  46.960000 24.395000  90.500000 ;
        RECT 0.495000  90.500000 24.245000  90.650000 ;
        RECT 0.495000  90.650000 24.095000  90.800000 ;
        RECT 0.495000  90.800000 23.945000  90.950000 ;
        RECT 0.495000  90.950000 23.795000  91.100000 ;
        RECT 0.495000  91.100000 23.645000  91.250000 ;
        RECT 0.495000  91.250000 23.495000  91.400000 ;
        RECT 0.495000  91.400000 23.345000  91.550000 ;
        RECT 0.495000  91.550000 23.195000  91.700000 ;
        RECT 0.495000  91.700000 23.045000  91.850000 ;
        RECT 0.495000  91.850000 22.895000  92.000000 ;
        RECT 0.495000  92.000000 22.745000  92.150000 ;
        RECT 0.495000  92.150000 22.595000  92.300000 ;
        RECT 0.495000  92.300000 22.445000  92.450000 ;
        RECT 0.495000  92.450000 22.295000  92.600000 ;
        RECT 0.495000  92.600000 22.145000  92.750000 ;
        RECT 0.495000  92.750000 21.995000  92.900000 ;
        RECT 0.495000  92.900000 21.845000  93.050000 ;
        RECT 0.495000  93.050000 21.695000  93.200000 ;
        RECT 0.495000  93.200000 21.545000  93.350000 ;
        RECT 0.495000  93.350000 21.395000  93.500000 ;
        RECT 0.495000  93.500000 21.245000  93.650000 ;
        RECT 0.495000  93.650000 21.095000  93.800000 ;
        RECT 0.495000  93.800000 20.945000  93.950000 ;
        RECT 0.495000  93.950000 20.795000  94.100000 ;
        RECT 0.495000  94.100000 20.645000  94.250000 ;
        RECT 0.495000  94.250000 20.495000  94.400000 ;
        RECT 0.495000  94.400000 20.345000  94.550000 ;
        RECT 0.495000  94.550000 20.195000  94.700000 ;
        RECT 0.495000  94.700000 20.045000  94.850000 ;
        RECT 0.495000  94.850000 19.895000  95.000000 ;
        RECT 0.495000  95.000000 19.745000  95.150000 ;
        RECT 0.495000  95.150000 19.595000  95.300000 ;
        RECT 0.495000  95.300000 19.445000  95.450000 ;
        RECT 0.495000  95.450000 19.295000  95.600000 ;
        RECT 0.495000  95.600000 19.145000  95.750000 ;
        RECT 0.495000  95.750000 18.995000  95.900000 ;
        RECT 0.495000  95.900000 18.845000  96.050000 ;
        RECT 0.495000  96.050000 18.695000  96.200000 ;
        RECT 0.495000  96.200000 18.545000  96.350000 ;
        RECT 0.495000  96.350000 18.395000  96.500000 ;
        RECT 0.495000  96.500000 18.245000  96.650000 ;
        RECT 0.495000  96.650000 18.095000  96.800000 ;
        RECT 0.495000  96.800000 17.945000  96.950000 ;
        RECT 0.495000  96.950000 17.795000  97.100000 ;
        RECT 0.495000  97.100000 17.645000  97.250000 ;
        RECT 0.495000  97.250000 17.495000  97.400000 ;
        RECT 0.495000  97.400000 17.345000  97.550000 ;
        RECT 0.495000  97.550000 17.195000  97.700000 ;
        RECT 0.495000  97.700000 17.045000  97.850000 ;
        RECT 0.495000  97.850000 16.895000  98.000000 ;
        RECT 0.495000  98.000000 16.745000  98.150000 ;
        RECT 0.495000  98.150000 16.595000  98.300000 ;
        RECT 0.495000  98.300000 16.445000  98.450000 ;
        RECT 0.495000  98.450000 16.295000  98.600000 ;
        RECT 0.495000  98.600000 16.145000  98.750000 ;
        RECT 0.495000  98.750000 15.995000  98.900000 ;
        RECT 0.495000  98.900000 15.845000  99.050000 ;
        RECT 0.495000  99.050000 15.695000  99.200000 ;
        RECT 0.495000  99.200000 15.545000  99.350000 ;
        RECT 0.495000  99.350000 15.395000  99.500000 ;
        RECT 0.495000  99.500000 15.245000  99.650000 ;
        RECT 0.495000  99.650000 15.095000  99.800000 ;
        RECT 0.495000  99.800000 14.945000  99.950000 ;
        RECT 0.495000  99.950000 14.795000 100.100000 ;
        RECT 0.495000 100.100000 14.645000 100.250000 ;
        RECT 0.495000 100.250000 14.495000 100.400000 ;
        RECT 0.495000 100.400000 14.345000 100.550000 ;
        RECT 0.495000 100.550000 14.195000 100.700000 ;
        RECT 0.495000 100.700000 14.045000 100.850000 ;
        RECT 0.495000 100.850000 13.895000 101.000000 ;
        RECT 0.495000 101.000000 13.745000 101.150000 ;
        RECT 0.495000 101.150000 13.595000 101.300000 ;
        RECT 0.495000 101.300000 13.500000 101.395000 ;
        RECT 0.495000 101.395000 13.500000 173.155000 ;
        RECT 0.520000  46.935000 24.395000  46.960000 ;
        RECT 0.645000  36.510000 24.395000  36.660000 ;
        RECT 0.670000  46.785000 24.395000  46.935000 ;
        RECT 0.795000  36.660000 24.395000  36.810000 ;
        RECT 0.820000  46.635000 24.395000  46.785000 ;
        RECT 0.945000  36.810000 24.395000  36.960000 ;
        RECT 0.970000  36.960000 24.395000  36.985000 ;
        RECT 0.970000  36.985000 24.395000  46.485000 ;
        RECT 0.970000  46.485000 24.395000  46.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000   0.000000 74.290000  90.185000 ;
        RECT 50.540000  90.185000 74.290000  90.335000 ;
        RECT 50.690000  90.335000 74.290000  90.485000 ;
        RECT 50.840000  90.485000 74.290000  90.635000 ;
        RECT 50.990000  90.635000 74.290000  90.785000 ;
        RECT 51.140000  90.785000 74.290000  90.935000 ;
        RECT 51.290000  90.935000 74.290000  91.085000 ;
        RECT 51.440000  91.085000 74.290000  91.235000 ;
        RECT 51.590000  91.235000 74.290000  91.385000 ;
        RECT 51.740000  91.385000 74.290000  91.535000 ;
        RECT 51.890000  91.535000 74.290000  91.685000 ;
        RECT 52.040000  91.685000 74.290000  91.835000 ;
        RECT 52.190000  91.835000 74.290000  91.985000 ;
        RECT 52.340000  91.985000 74.290000  92.135000 ;
        RECT 52.490000  92.135000 74.290000  92.285000 ;
        RECT 52.640000  92.285000 74.290000  92.435000 ;
        RECT 52.790000  92.435000 74.290000  92.585000 ;
        RECT 52.940000  92.585000 74.290000  92.735000 ;
        RECT 53.090000  92.735000 74.290000  92.885000 ;
        RECT 53.240000  92.885000 74.290000  93.035000 ;
        RECT 53.390000  93.035000 74.290000  93.185000 ;
        RECT 53.540000  93.185000 74.290000  93.335000 ;
        RECT 53.690000  93.335000 74.290000  93.485000 ;
        RECT 53.840000  93.485000 74.290000  93.635000 ;
        RECT 53.990000  93.635000 74.290000  93.785000 ;
        RECT 54.140000  93.785000 74.290000  93.935000 ;
        RECT 54.290000  93.935000 74.290000  94.085000 ;
        RECT 54.440000  94.085000 74.290000  94.235000 ;
        RECT 54.590000  94.235000 74.290000  94.385000 ;
        RECT 54.740000  94.385000 74.290000  94.535000 ;
        RECT 54.890000  94.535000 74.290000  94.685000 ;
        RECT 55.040000  94.685000 74.290000  94.835000 ;
        RECT 55.190000  94.835000 74.290000  94.985000 ;
        RECT 55.340000  94.985000 74.290000  95.135000 ;
        RECT 55.490000  95.135000 74.290000  95.285000 ;
        RECT 55.640000  95.285000 74.290000  95.435000 ;
        RECT 55.790000  95.435000 74.290000  95.585000 ;
        RECT 55.940000  95.585000 74.290000  95.735000 ;
        RECT 56.090000  95.735000 74.290000  95.885000 ;
        RECT 56.240000  95.885000 74.290000  96.035000 ;
        RECT 56.390000  96.035000 74.290000  96.185000 ;
        RECT 56.540000  96.185000 74.290000  96.335000 ;
        RECT 56.690000  96.335000 74.290000  96.485000 ;
        RECT 56.840000  96.485000 74.290000  96.635000 ;
        RECT 56.990000  96.635000 74.290000  96.785000 ;
        RECT 57.140000  96.785000 74.290000  96.935000 ;
        RECT 57.290000  96.935000 74.290000  97.085000 ;
        RECT 57.440000  97.085000 74.290000  97.235000 ;
        RECT 57.590000  97.235000 74.290000  97.385000 ;
        RECT 57.740000  97.385000 74.290000  97.535000 ;
        RECT 57.890000  97.535000 74.290000  97.685000 ;
        RECT 58.040000  97.685000 74.290000  97.835000 ;
        RECT 58.190000  97.835000 74.290000  97.985000 ;
        RECT 58.340000  97.985000 74.290000  98.135000 ;
        RECT 58.490000  98.135000 74.290000  98.285000 ;
        RECT 58.640000  98.285000 74.290000  98.435000 ;
        RECT 58.790000  98.435000 74.290000  98.585000 ;
        RECT 58.940000  98.585000 74.290000  98.735000 ;
        RECT 59.090000  98.735000 74.290000  98.885000 ;
        RECT 59.240000  98.885000 74.290000  99.035000 ;
        RECT 59.390000  99.035000 74.290000  99.185000 ;
        RECT 59.540000  99.185000 74.290000  99.335000 ;
        RECT 59.690000  99.335000 74.290000  99.485000 ;
        RECT 59.840000  99.485000 74.290000  99.635000 ;
        RECT 59.990000  99.635000 74.290000  99.785000 ;
        RECT 60.140000  99.785000 74.290000  99.935000 ;
        RECT 60.290000  99.935000 74.290000 100.085000 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
        RECT 61.490000 101.135000 74.290000 101.285000 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END G_CORE
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.495000   0.000000 24.395000   2.055000 ;
        RECT  0.565000   2.055000 24.395000   2.125000 ;
        RECT  0.635000   2.125000 24.395000   2.195000 ;
        RECT  0.705000   2.195000 24.395000   2.265000 ;
        RECT  0.775000   2.265000 24.395000   2.335000 ;
        RECT  0.845000   2.335000 24.395000   2.405000 ;
        RECT  0.915000   2.405000 24.395000   2.475000 ;
        RECT  0.985000   2.475000 24.395000   2.545000 ;
        RECT  1.005000   2.545000 24.395000   2.565000 ;
        RECT  1.005000   2.565000 24.395000   8.595000 ;
        RECT  1.005000   8.595000 24.395000   8.665000 ;
        RECT  1.005000   8.665000 24.465000   8.735000 ;
        RECT  1.005000   8.735000 24.535000   8.805000 ;
        RECT  1.005000   8.805000 24.605000   8.875000 ;
        RECT  1.005000   8.875000 24.675000   8.945000 ;
        RECT  1.005000   8.945000 24.745000   9.015000 ;
        RECT  1.005000   9.015000 24.815000   9.085000 ;
        RECT  1.005000   9.085000 24.885000   9.155000 ;
        RECT  1.005000   9.155000 24.955000   9.225000 ;
        RECT  1.005000   9.225000 25.025000   9.295000 ;
        RECT  1.005000   9.295000 25.095000   9.365000 ;
        RECT  1.005000   9.365000 25.165000   9.435000 ;
        RECT  1.005000   9.435000 25.235000   9.505000 ;
        RECT  1.005000   9.505000 25.305000   9.575000 ;
        RECT  1.005000   9.575000 25.375000   9.645000 ;
        RECT  1.005000   9.645000 25.445000   9.715000 ;
        RECT  1.005000   9.715000 25.515000   9.785000 ;
        RECT  1.005000   9.785000 25.585000   9.855000 ;
        RECT  1.005000   9.855000 25.655000   9.925000 ;
        RECT  1.005000   9.925000 25.725000   9.995000 ;
        RECT  1.005000   9.995000 25.795000  10.065000 ;
        RECT  1.005000  10.065000 25.865000  10.135000 ;
        RECT  1.005000  10.135000 25.935000  10.205000 ;
        RECT  1.005000  10.205000 26.005000  10.275000 ;
        RECT  1.005000  10.275000 26.075000  10.345000 ;
        RECT  1.005000  10.345000 26.145000  10.415000 ;
        RECT  1.005000  10.415000 26.215000  10.485000 ;
        RECT  1.005000  10.485000 26.285000  10.555000 ;
        RECT  1.005000  10.555000 26.355000  10.625000 ;
        RECT  1.005000  10.625000 26.425000  10.695000 ;
        RECT  1.005000  10.695000 26.495000  10.765000 ;
        RECT  1.005000  10.765000 26.565000  10.835000 ;
        RECT  1.005000  10.835000 26.635000  10.905000 ;
        RECT  1.005000  10.905000 26.705000  10.975000 ;
        RECT  1.005000  10.975000 26.775000  11.045000 ;
        RECT  1.005000  11.045000 26.845000  11.115000 ;
        RECT  1.005000  11.115000 26.915000  11.185000 ;
        RECT  1.005000  11.185000 26.985000  11.255000 ;
        RECT  1.005000  11.255000 27.055000  11.325000 ;
        RECT  1.005000  11.325000 27.125000  11.395000 ;
        RECT  1.005000  11.395000 27.195000  11.465000 ;
        RECT  1.005000  11.465000 27.265000  11.535000 ;
        RECT  1.005000  11.535000 27.335000  11.605000 ;
        RECT  1.005000  11.605000 27.405000  11.675000 ;
        RECT  1.005000  11.675000 27.475000  11.745000 ;
        RECT  1.005000  11.745000 27.545000  11.815000 ;
        RECT  1.005000  11.815000 27.615000  11.885000 ;
        RECT  1.005000  11.885000 27.685000  11.955000 ;
        RECT  1.005000  11.955000 27.755000  12.025000 ;
        RECT  1.005000  12.025000 27.825000  12.095000 ;
        RECT  1.005000  12.095000 27.895000  12.165000 ;
        RECT  1.005000  12.165000 27.965000  12.235000 ;
        RECT  1.005000  12.235000 28.035000  12.305000 ;
        RECT  1.005000  12.305000 28.105000  12.375000 ;
        RECT  1.005000  12.375000 28.175000  12.400000 ;
        RECT  1.005000  12.400000 36.895000  25.700000 ;
        RECT  1.005000  25.700000 18.750000  25.770000 ;
        RECT  1.005000  25.770000 18.680000  25.840000 ;
        RECT  1.005000  25.840000 18.610000  25.910000 ;
        RECT  1.005000  25.910000 18.540000  25.980000 ;
        RECT  1.005000  25.980000 18.470000  26.050000 ;
        RECT  1.005000  26.050000 18.400000  26.120000 ;
        RECT  1.005000  26.120000 18.330000  26.190000 ;
        RECT  1.005000  26.190000 18.260000  26.260000 ;
        RECT  1.005000  26.260000 18.190000  26.330000 ;
        RECT  1.005000  26.330000 18.120000  26.400000 ;
        RECT  1.005000  26.400000 18.050000  26.470000 ;
        RECT  1.005000  26.470000 17.980000  26.540000 ;
        RECT  1.005000  26.540000 17.910000  26.610000 ;
        RECT  1.005000  26.610000 17.840000  26.680000 ;
        RECT  1.005000  26.680000 17.770000  26.750000 ;
        RECT  1.005000  26.750000 17.700000  26.820000 ;
        RECT  1.005000  26.820000 17.630000  26.890000 ;
        RECT  1.005000  26.890000 17.560000  26.960000 ;
        RECT  1.005000  26.960000 17.490000  27.030000 ;
        RECT  1.005000  27.030000 17.420000  27.100000 ;
        RECT  1.005000  27.100000 17.350000  27.170000 ;
        RECT  1.005000  27.170000 17.280000  27.240000 ;
        RECT  1.005000  27.240000 17.210000  27.310000 ;
        RECT  1.005000  27.310000 17.140000  27.380000 ;
        RECT  1.005000  27.380000 17.070000  27.450000 ;
        RECT  1.005000  27.450000 17.000000  27.520000 ;
        RECT  1.005000  27.520000 16.930000  27.590000 ;
        RECT  1.005000  27.590000 16.860000  27.660000 ;
        RECT  1.005000  27.660000 16.790000  27.730000 ;
        RECT  1.005000  27.730000 16.720000  27.800000 ;
        RECT  1.005000  27.800000 16.650000  27.870000 ;
        RECT  1.005000  27.870000 16.580000  27.940000 ;
        RECT  1.005000  27.940000 16.510000  28.010000 ;
        RECT  1.005000  28.010000 16.440000  28.080000 ;
        RECT  1.005000  28.080000 16.370000  28.150000 ;
        RECT  1.005000  28.150000 16.300000  28.220000 ;
        RECT  1.005000  28.220000 16.230000  28.290000 ;
        RECT  1.005000  28.290000 16.160000  28.360000 ;
        RECT  1.005000  28.360000 16.090000  28.430000 ;
        RECT  1.005000  28.430000 16.020000  28.500000 ;
        RECT  1.005000  28.500000 15.950000  28.570000 ;
        RECT  1.005000  28.570000 15.880000  28.640000 ;
        RECT  1.005000  28.640000 15.810000  28.710000 ;
        RECT  1.005000  28.710000 15.740000  28.780000 ;
        RECT  1.005000  28.780000 15.670000  28.850000 ;
        RECT  1.005000  28.850000 15.600000  28.920000 ;
        RECT  1.005000  28.920000 15.530000  28.990000 ;
        RECT  1.005000  28.990000 15.460000  29.060000 ;
        RECT  1.005000  29.060000 15.390000  29.130000 ;
        RECT  1.005000  29.130000 15.320000  29.200000 ;
        RECT  1.005000  29.200000 15.250000  29.270000 ;
        RECT  1.005000  29.270000 15.205000  29.315000 ;
        RECT  1.005000  29.315000 15.205000  35.665000 ;
        RECT  1.005000  35.665000 15.205000  35.735000 ;
        RECT  1.005000  35.735000 15.275000  35.805000 ;
        RECT  1.005000  35.805000 15.345000  35.875000 ;
        RECT  1.005000  35.875000 15.415000  35.945000 ;
        RECT  1.005000  35.945000 15.485000  36.015000 ;
        RECT  1.005000  36.015000 15.555000  36.085000 ;
        RECT  1.005000  36.085000 15.625000  36.155000 ;
        RECT  1.005000  36.155000 15.695000  36.225000 ;
        RECT  1.005000  36.225000 15.765000  36.295000 ;
        RECT  1.005000  36.295000 15.835000  36.365000 ;
        RECT  1.005000  36.365000 15.905000  36.435000 ;
        RECT  1.005000  36.435000 15.975000  36.505000 ;
        RECT  1.005000  36.505000 16.045000  36.575000 ;
        RECT  1.005000  36.575000 16.115000  36.640000 ;
        RECT  1.005000  47.130000 14.120000  54.215000 ;
        RECT  1.005000  54.215000 14.120000  54.285000 ;
        RECT  1.005000  54.285000 14.190000  54.355000 ;
        RECT  1.005000  54.355000 14.260000  54.425000 ;
        RECT  1.005000  54.425000 14.330000  54.495000 ;
        RECT  1.005000  54.495000 14.400000  54.565000 ;
        RECT  1.005000  54.565000 14.470000  54.635000 ;
        RECT  1.005000  54.635000 14.540000  54.705000 ;
        RECT  1.005000  54.705000 14.610000  54.775000 ;
        RECT  1.005000  54.775000 14.680000  54.845000 ;
        RECT  1.005000  54.845000 14.750000  54.915000 ;
        RECT  1.005000  54.915000 14.820000  54.985000 ;
        RECT  1.005000  54.985000 14.890000  55.055000 ;
        RECT  1.005000  55.055000 14.960000  55.125000 ;
        RECT  1.005000  55.125000 15.030000  55.195000 ;
        RECT  1.005000  55.195000 15.100000  55.265000 ;
        RECT  1.005000  55.265000 15.170000  55.335000 ;
        RECT  1.005000  55.335000 15.240000  55.405000 ;
        RECT  1.005000  55.405000 15.310000  55.475000 ;
        RECT  1.005000  55.475000 15.380000  55.545000 ;
        RECT  1.005000  55.545000 15.450000  55.615000 ;
        RECT  1.005000  55.615000 15.520000  55.685000 ;
        RECT  1.005000  55.685000 15.590000  55.755000 ;
        RECT  1.005000  55.755000 15.660000  55.825000 ;
        RECT  1.005000  55.825000 15.730000  55.895000 ;
        RECT  1.005000  55.895000 15.800000  55.965000 ;
        RECT  1.005000  55.965000 15.870000  56.035000 ;
        RECT  1.005000  56.035000 15.940000  56.105000 ;
        RECT  1.005000  56.105000 16.010000  56.175000 ;
        RECT  1.005000  56.175000 16.080000  56.245000 ;
        RECT  1.005000  56.245000 16.150000  56.315000 ;
        RECT  1.005000  56.315000 16.220000  56.385000 ;
        RECT  1.005000  56.385000 16.290000  56.455000 ;
        RECT  1.005000  56.455000 16.360000  56.525000 ;
        RECT  1.005000  56.525000 16.430000  56.595000 ;
        RECT  1.005000  56.595000 16.500000  56.665000 ;
        RECT  1.005000  56.665000 16.570000  56.735000 ;
        RECT  1.005000  56.735000 16.640000  56.805000 ;
        RECT  1.005000  56.805000 16.710000  56.875000 ;
        RECT  1.005000  56.875000 16.780000  56.945000 ;
        RECT  1.005000  56.945000 16.850000  57.015000 ;
        RECT  1.005000  57.015000 16.920000  57.085000 ;
        RECT  1.005000  57.085000 16.990000  57.155000 ;
        RECT  1.005000  57.155000 17.060000  57.225000 ;
        RECT  1.005000  57.225000 17.130000  57.295000 ;
        RECT  1.005000  57.295000 17.200000  57.365000 ;
        RECT  1.005000  57.365000 17.270000  57.435000 ;
        RECT  1.005000  57.435000 17.340000  57.505000 ;
        RECT  1.005000  57.505000 17.410000  57.575000 ;
        RECT  1.005000  57.575000 17.480000  57.645000 ;
        RECT  1.005000  57.645000 17.550000  57.715000 ;
        RECT  1.005000  57.715000 17.620000  57.780000 ;
        RECT  1.005000  57.780000 56.710000  66.480000 ;
        RECT  1.005000  66.480000 17.595000  66.550000 ;
        RECT  1.005000  66.550000 17.525000  66.620000 ;
        RECT  1.005000  66.620000 17.455000  66.690000 ;
        RECT  1.005000  66.690000 17.385000  66.760000 ;
        RECT  1.005000  66.760000 17.315000  66.830000 ;
        RECT  1.005000  66.830000 17.245000  66.900000 ;
        RECT  1.005000  66.900000 17.175000  66.970000 ;
        RECT  1.005000  66.970000 17.105000  67.040000 ;
        RECT  1.005000  67.040000 17.035000  67.110000 ;
        RECT  1.005000  67.110000 16.965000  67.180000 ;
        RECT  1.005000  67.180000 16.895000  67.250000 ;
        RECT  1.005000  67.250000 16.825000  67.320000 ;
        RECT  1.005000  67.320000 16.755000  67.390000 ;
        RECT  1.005000  67.390000 16.685000  67.460000 ;
        RECT  1.005000  67.460000 16.615000  67.530000 ;
        RECT  1.005000  67.530000 16.545000  67.600000 ;
        RECT  1.005000  67.600000 16.475000  67.670000 ;
        RECT  1.005000  67.670000 16.405000  67.740000 ;
        RECT  1.005000  67.740000 16.335000  67.810000 ;
        RECT  1.005000  67.810000 16.265000  67.880000 ;
        RECT  1.005000  67.880000 16.195000  67.950000 ;
        RECT  1.005000  67.950000 16.125000  68.020000 ;
        RECT  1.005000  68.020000 16.055000  68.090000 ;
        RECT  1.005000  68.090000 15.985000  68.160000 ;
        RECT  1.005000  68.160000 15.915000  68.230000 ;
        RECT  1.005000  68.230000 15.845000  68.300000 ;
        RECT  1.005000  68.300000 15.775000  68.370000 ;
        RECT  1.005000  68.370000 15.705000  68.440000 ;
        RECT  1.005000  68.440000 15.635000  68.510000 ;
        RECT  1.005000  68.510000 15.565000  68.580000 ;
        RECT  1.005000  68.580000 15.495000  68.650000 ;
        RECT  1.005000  68.650000 15.425000  68.720000 ;
        RECT  1.005000  68.720000 15.355000  68.790000 ;
        RECT  1.005000  68.790000 15.285000  68.860000 ;
        RECT  1.005000  68.860000 15.215000  68.930000 ;
        RECT  1.005000  68.930000 15.145000  69.000000 ;
        RECT  1.005000  69.000000 15.075000  69.070000 ;
        RECT  1.005000  69.070000 15.005000  69.140000 ;
        RECT  1.005000  69.140000 14.935000  69.210000 ;
        RECT  1.005000  69.210000 14.865000  69.280000 ;
        RECT  1.005000  69.280000 14.795000  69.350000 ;
        RECT  1.005000  69.350000 14.725000  69.420000 ;
        RECT  1.005000  69.420000 14.655000  69.490000 ;
        RECT  1.005000  69.490000 14.585000  69.560000 ;
        RECT  1.005000  69.560000 14.515000  69.630000 ;
        RECT  1.005000  69.630000 14.445000  69.700000 ;
        RECT  1.005000  69.700000 14.375000  69.770000 ;
        RECT  1.005000  69.770000 14.305000  69.840000 ;
        RECT  1.005000  69.840000 14.235000  69.910000 ;
        RECT  1.005000  69.910000 14.165000  69.980000 ;
        RECT  1.005000  69.980000 14.120000  70.025000 ;
        RECT  1.005000  70.025000 14.120000  77.240000 ;
        RECT  1.005000  77.240000 14.120000  77.310000 ;
        RECT  1.005000  77.310000 14.190000  77.380000 ;
        RECT  1.005000  77.380000 14.260000  77.450000 ;
        RECT  1.005000  77.450000 14.330000  77.520000 ;
        RECT  1.005000  77.520000 14.400000  77.590000 ;
        RECT  1.005000  77.590000 14.470000  77.660000 ;
        RECT  1.005000  77.660000 14.540000  77.730000 ;
        RECT  1.005000  77.730000 14.610000  77.800000 ;
        RECT  1.005000  77.800000 14.680000  77.870000 ;
        RECT  1.005000  77.870000 14.750000  77.940000 ;
        RECT  1.005000  77.940000 14.820000  78.010000 ;
        RECT  1.005000  78.010000 14.890000  78.080000 ;
        RECT  1.005000  78.080000 14.960000  78.150000 ;
        RECT  1.005000  78.150000 15.030000  78.220000 ;
        RECT  1.005000  78.220000 15.100000  78.290000 ;
        RECT  1.005000  78.290000 15.170000  78.360000 ;
        RECT  1.005000  78.360000 15.240000  78.430000 ;
        RECT  1.005000  78.430000 15.310000  78.500000 ;
        RECT  1.005000  78.500000 15.380000  78.570000 ;
        RECT  1.005000  78.570000 15.450000  78.640000 ;
        RECT  1.005000  78.640000 15.520000  78.710000 ;
        RECT  1.005000  78.710000 15.590000  78.780000 ;
        RECT  1.005000  78.780000 15.660000  78.850000 ;
        RECT  1.005000  78.850000 15.730000  78.920000 ;
        RECT  1.005000  78.920000 15.800000  78.990000 ;
        RECT  1.005000  78.990000 15.870000  79.060000 ;
        RECT  1.005000  79.060000 15.940000  79.130000 ;
        RECT  1.005000  79.130000 16.010000  79.200000 ;
        RECT  1.005000  79.200000 16.080000  79.270000 ;
        RECT  1.005000  79.270000 16.150000  79.340000 ;
        RECT  1.005000  79.340000 16.220000  79.410000 ;
        RECT  1.005000  79.410000 16.290000  79.480000 ;
        RECT  1.005000  79.480000 16.360000  79.550000 ;
        RECT  1.005000  79.550000 16.430000  79.620000 ;
        RECT  1.005000  79.620000 16.500000  79.690000 ;
        RECT  1.005000  79.690000 16.570000  79.760000 ;
        RECT  1.005000  79.760000 16.640000  79.830000 ;
        RECT  1.005000  79.830000 16.710000  79.900000 ;
        RECT  1.005000  79.900000 16.780000  79.970000 ;
        RECT  1.005000  79.970000 16.850000  80.040000 ;
        RECT  1.005000  80.040000 16.920000  80.110000 ;
        RECT  1.005000  80.110000 16.990000  80.180000 ;
        RECT  1.005000  80.180000 17.060000  80.250000 ;
        RECT  1.005000  80.250000 17.130000  80.320000 ;
        RECT  1.005000  80.320000 17.200000  80.390000 ;
        RECT  1.005000  80.390000 17.270000  80.460000 ;
        RECT  1.005000  80.460000 17.340000  80.530000 ;
        RECT  1.005000  80.530000 17.410000  80.600000 ;
        RECT  1.005000  80.600000 17.480000  80.670000 ;
        RECT  1.005000  80.670000 17.550000  80.740000 ;
        RECT  1.005000  80.740000 17.620000  80.780000 ;
        RECT  1.005000  80.780000 56.705000  89.480000 ;
        RECT  1.005000  89.480000 17.595000  89.550000 ;
        RECT  1.005000  89.550000 17.525000  89.620000 ;
        RECT  1.005000  89.620000 17.455000  89.690000 ;
        RECT  1.005000  89.690000 17.385000  89.760000 ;
        RECT  1.005000  89.760000 17.315000  89.830000 ;
        RECT  1.005000  89.830000 17.245000  89.900000 ;
        RECT  1.005000  89.900000 17.175000  89.970000 ;
        RECT  1.005000  89.970000 17.105000  90.040000 ;
        RECT  1.005000  90.040000 17.035000  90.110000 ;
        RECT  1.005000  90.110000 16.965000  90.180000 ;
        RECT  1.005000  90.180000 16.895000  90.250000 ;
        RECT  1.005000  90.250000 16.825000  90.320000 ;
        RECT  1.005000  90.320000 16.755000  90.390000 ;
        RECT  1.005000  90.390000 16.685000  90.460000 ;
        RECT  1.005000  90.460000 16.615000  90.530000 ;
        RECT  1.005000  90.530000 16.545000  90.600000 ;
        RECT  1.005000  90.600000 16.475000  90.670000 ;
        RECT  1.005000  90.670000 16.405000  90.740000 ;
        RECT  1.005000  90.740000 16.335000  90.810000 ;
        RECT  1.005000  90.810000 16.265000  90.880000 ;
        RECT  1.005000  90.880000 16.195000  90.950000 ;
        RECT  1.005000  90.950000 16.125000  91.020000 ;
        RECT  1.005000  91.020000 16.055000  91.090000 ;
        RECT  1.005000  91.090000 15.985000  91.160000 ;
        RECT  1.005000  91.160000 15.915000  91.230000 ;
        RECT  1.005000  91.230000 15.845000  91.300000 ;
        RECT  1.005000  91.300000 15.775000  91.370000 ;
        RECT  1.005000  91.370000 15.705000  91.440000 ;
        RECT  1.005000  91.440000 15.635000  91.510000 ;
        RECT  1.005000  91.510000 15.565000  91.580000 ;
        RECT  1.005000  91.580000 15.495000  91.650000 ;
        RECT  1.005000  91.650000 15.425000  91.720000 ;
        RECT  1.005000  91.720000 15.355000  91.790000 ;
        RECT  1.005000  91.790000 15.285000  91.860000 ;
        RECT  1.005000  91.860000 15.215000  91.930000 ;
        RECT  1.005000  91.930000 15.145000  92.000000 ;
        RECT  1.005000  92.000000 15.075000  92.070000 ;
        RECT  1.005000  92.070000 15.005000  92.140000 ;
        RECT  1.005000  92.140000 14.935000  92.210000 ;
        RECT  1.005000  92.210000 14.865000  92.280000 ;
        RECT  1.005000  92.280000 14.795000  92.350000 ;
        RECT  1.005000  92.350000 14.725000  92.420000 ;
        RECT  1.005000  92.420000 14.655000  92.490000 ;
        RECT  1.005000  92.490000 14.585000  92.560000 ;
        RECT  1.005000  92.560000 14.515000  92.630000 ;
        RECT  1.005000  92.630000 14.445000  92.700000 ;
        RECT  1.005000  92.700000 14.375000  92.770000 ;
        RECT  1.005000  92.770000 14.305000  92.840000 ;
        RECT  1.005000  92.840000 14.235000  92.910000 ;
        RECT  1.005000  92.910000 14.165000  92.980000 ;
        RECT  1.005000  92.980000 14.120000  93.025000 ;
        RECT  1.005000  93.025000 14.120000 100.240000 ;
        RECT  1.005000 100.240000 14.120000 100.310000 ;
        RECT  1.005000 100.310000 14.190000 100.380000 ;
        RECT  1.005000 100.380000 14.260000 100.450000 ;
        RECT  1.005000 100.450000 14.330000 100.520000 ;
        RECT  1.005000 100.520000 14.400000 100.590000 ;
        RECT  1.005000 100.590000 14.470000 100.660000 ;
        RECT  1.005000 100.660000 14.540000 100.730000 ;
        RECT  1.005000 100.730000 14.610000 100.800000 ;
        RECT  1.005000 100.800000 14.680000 100.870000 ;
        RECT  1.005000 100.870000 14.750000 100.940000 ;
        RECT  1.005000 100.940000 14.820000 101.010000 ;
        RECT  1.005000 101.010000 14.890000 101.080000 ;
        RECT  1.005000 101.080000 14.960000 101.150000 ;
        RECT  1.005000 101.150000 15.030000 101.220000 ;
        RECT  1.005000 101.220000 15.100000 101.290000 ;
        RECT  1.005000 101.290000 15.170000 101.360000 ;
        RECT  1.005000 101.360000 15.240000 101.430000 ;
        RECT  1.005000 101.430000 15.310000 101.500000 ;
        RECT  1.005000 101.500000 15.380000 101.570000 ;
        RECT  1.005000 101.570000 15.450000 101.640000 ;
        RECT  1.005000 101.640000 15.520000 101.710000 ;
        RECT  1.005000 101.710000 15.590000 101.780000 ;
        RECT  1.005000 101.780000 15.660000 101.850000 ;
        RECT  1.005000 101.850000 15.730000 101.920000 ;
        RECT  1.005000 101.920000 15.800000 101.990000 ;
        RECT  1.005000 101.990000 15.870000 102.060000 ;
        RECT  1.005000 102.060000 15.940000 102.130000 ;
        RECT  1.005000 102.130000 16.010000 102.200000 ;
        RECT  1.005000 102.200000 16.080000 102.270000 ;
        RECT  1.005000 102.270000 16.150000 102.340000 ;
        RECT  1.005000 102.340000 16.220000 102.410000 ;
        RECT  1.005000 102.410000 16.290000 102.480000 ;
        RECT  1.005000 102.480000 16.360000 102.550000 ;
        RECT  1.005000 102.550000 16.430000 102.620000 ;
        RECT  1.005000 102.620000 16.500000 102.690000 ;
        RECT  1.005000 102.690000 16.570000 102.760000 ;
        RECT  1.005000 102.760000 16.640000 102.830000 ;
        RECT  1.005000 102.830000 16.710000 102.900000 ;
        RECT  1.005000 102.900000 16.780000 102.970000 ;
        RECT  1.005000 102.970000 16.850000 103.040000 ;
        RECT  1.005000 103.040000 16.920000 103.110000 ;
        RECT  1.005000 103.110000 16.990000 103.180000 ;
        RECT  1.005000 103.180000 17.060000 103.250000 ;
        RECT  1.005000 103.250000 17.130000 103.320000 ;
        RECT  1.005000 103.320000 17.200000 103.390000 ;
        RECT  1.005000 103.390000 17.270000 103.460000 ;
        RECT  1.005000 103.460000 17.340000 103.530000 ;
        RECT  1.005000 103.530000 17.410000 103.600000 ;
        RECT  1.005000 103.600000 17.480000 103.670000 ;
        RECT  1.005000 103.670000 17.550000 103.740000 ;
        RECT  1.005000 103.740000 17.620000 103.780000 ;
        RECT  1.005000 103.780000 56.705000 112.480000 ;
        RECT  1.005000 112.480000 17.635000 112.550000 ;
        RECT  1.005000 112.550000 17.565000 112.620000 ;
        RECT  1.005000 112.620000 17.495000 112.690000 ;
        RECT  1.005000 112.690000 17.425000 112.760000 ;
        RECT  1.005000 112.760000 17.355000 112.830000 ;
        RECT  1.005000 112.830000 17.285000 112.900000 ;
        RECT  1.005000 112.900000 17.215000 112.970000 ;
        RECT  1.005000 112.970000 17.145000 113.040000 ;
        RECT  1.005000 113.040000 17.075000 113.110000 ;
        RECT  1.005000 113.110000 17.005000 113.180000 ;
        RECT  1.005000 113.180000 16.935000 113.250000 ;
        RECT  1.005000 113.250000 16.865000 113.320000 ;
        RECT  1.005000 113.320000 16.795000 113.390000 ;
        RECT  1.005000 113.390000 16.725000 113.460000 ;
        RECT  1.005000 113.460000 16.655000 113.530000 ;
        RECT  1.005000 113.530000 16.585000 113.600000 ;
        RECT  1.005000 113.600000 16.515000 113.670000 ;
        RECT  1.005000 113.670000 16.445000 113.740000 ;
        RECT  1.005000 113.740000 16.375000 113.810000 ;
        RECT  1.005000 113.810000 16.305000 113.880000 ;
        RECT  1.005000 113.880000 16.235000 113.950000 ;
        RECT  1.005000 113.950000 16.165000 114.020000 ;
        RECT  1.005000 114.020000 16.095000 114.090000 ;
        RECT  1.005000 114.090000 16.025000 114.160000 ;
        RECT  1.005000 114.160000 15.955000 114.230000 ;
        RECT  1.005000 114.230000 15.885000 114.300000 ;
        RECT  1.005000 114.300000 15.815000 114.370000 ;
        RECT  1.005000 114.370000 15.745000 114.440000 ;
        RECT  1.005000 114.440000 15.675000 114.510000 ;
        RECT  1.005000 114.510000 15.605000 114.580000 ;
        RECT  1.005000 114.580000 15.535000 114.650000 ;
        RECT  1.005000 114.650000 15.465000 114.720000 ;
        RECT  1.005000 114.720000 15.395000 114.790000 ;
        RECT  1.005000 114.790000 15.325000 114.860000 ;
        RECT  1.005000 114.860000 15.255000 114.930000 ;
        RECT  1.005000 114.930000 15.185000 115.000000 ;
        RECT  1.005000 115.000000 15.115000 115.070000 ;
        RECT  1.005000 115.070000 15.045000 115.140000 ;
        RECT  1.005000 115.140000 14.975000 115.210000 ;
        RECT  1.005000 115.210000 14.905000 115.280000 ;
        RECT  1.005000 115.280000 14.835000 115.350000 ;
        RECT  1.005000 115.350000 14.765000 115.420000 ;
        RECT  1.005000 115.420000 14.695000 115.490000 ;
        RECT  1.005000 115.490000 14.625000 115.560000 ;
        RECT  1.005000 115.560000 14.555000 115.630000 ;
        RECT  1.005000 115.630000 14.485000 115.700000 ;
        RECT  1.005000 115.700000 14.415000 115.770000 ;
        RECT  1.005000 115.770000 14.345000 115.840000 ;
        RECT  1.005000 115.840000 14.275000 115.910000 ;
        RECT  1.005000 115.910000 14.205000 115.980000 ;
        RECT  1.005000 115.980000 14.135000 116.050000 ;
        RECT  1.005000 116.050000 14.120000 116.065000 ;
        RECT  1.005000 116.065000 14.120000 123.145000 ;
        RECT  1.005000 123.145000 14.120000 123.215000 ;
        RECT  1.005000 123.215000 14.190000 123.285000 ;
        RECT  1.005000 123.285000 14.260000 123.355000 ;
        RECT  1.005000 123.355000 14.330000 123.425000 ;
        RECT  1.005000 123.425000 14.400000 123.495000 ;
        RECT  1.005000 123.495000 14.470000 123.565000 ;
        RECT  1.005000 123.565000 14.540000 123.635000 ;
        RECT  1.005000 123.635000 14.610000 123.705000 ;
        RECT  1.005000 123.705000 14.680000 123.775000 ;
        RECT  1.005000 123.775000 14.750000 123.845000 ;
        RECT  1.005000 123.845000 14.820000 123.915000 ;
        RECT  1.005000 123.915000 14.890000 123.985000 ;
        RECT  1.005000 123.985000 14.960000 124.055000 ;
        RECT  1.005000 124.055000 15.030000 124.125000 ;
        RECT  1.005000 124.125000 15.100000 124.195000 ;
        RECT  1.005000 124.195000 15.170000 124.265000 ;
        RECT  1.005000 124.265000 15.240000 124.335000 ;
        RECT  1.005000 124.335000 15.310000 124.405000 ;
        RECT  1.005000 124.405000 15.380000 124.475000 ;
        RECT  1.005000 124.475000 15.450000 124.545000 ;
        RECT  1.005000 124.545000 15.520000 124.615000 ;
        RECT  1.005000 124.615000 15.590000 124.685000 ;
        RECT  1.005000 124.685000 15.660000 124.755000 ;
        RECT  1.005000 124.755000 15.730000 124.825000 ;
        RECT  1.005000 124.825000 15.800000 124.895000 ;
        RECT  1.005000 124.895000 15.870000 124.965000 ;
        RECT  1.005000 124.965000 15.940000 125.035000 ;
        RECT  1.005000 125.035000 16.010000 125.105000 ;
        RECT  1.005000 125.105000 16.080000 125.175000 ;
        RECT  1.005000 125.175000 16.150000 125.245000 ;
        RECT  1.005000 125.245000 16.220000 125.315000 ;
        RECT  1.005000 125.315000 16.290000 125.385000 ;
        RECT  1.005000 125.385000 16.360000 125.455000 ;
        RECT  1.005000 125.455000 16.430000 125.525000 ;
        RECT  1.005000 125.525000 16.500000 125.595000 ;
        RECT  1.005000 125.595000 16.570000 125.665000 ;
        RECT  1.005000 125.665000 16.640000 125.735000 ;
        RECT  1.005000 125.735000 16.710000 125.805000 ;
        RECT  1.005000 125.805000 16.780000 125.875000 ;
        RECT  1.005000 125.875000 16.850000 125.945000 ;
        RECT  1.005000 125.945000 16.920000 126.015000 ;
        RECT  1.005000 126.015000 16.990000 126.085000 ;
        RECT  1.005000 126.085000 17.060000 126.155000 ;
        RECT  1.005000 126.155000 17.130000 126.225000 ;
        RECT  1.005000 126.225000 17.200000 126.295000 ;
        RECT  1.005000 126.295000 17.270000 126.365000 ;
        RECT  1.005000 126.365000 17.340000 126.435000 ;
        RECT  1.005000 126.435000 17.410000 126.505000 ;
        RECT  1.005000 126.505000 17.480000 126.575000 ;
        RECT  1.005000 126.575000 17.550000 126.645000 ;
        RECT  1.005000 126.645000 17.620000 126.715000 ;
        RECT  1.005000 126.715000 17.690000 126.780000 ;
        RECT  1.005000 126.780000 56.705000 135.480000 ;
        RECT  1.005000 135.480000 17.740000 135.550000 ;
        RECT  1.005000 135.550000 17.670000 135.620000 ;
        RECT  1.005000 135.620000 17.600000 135.690000 ;
        RECT  1.005000 135.690000 17.530000 135.760000 ;
        RECT  1.005000 135.760000 17.460000 135.830000 ;
        RECT  1.005000 135.830000 17.390000 135.900000 ;
        RECT  1.005000 135.900000 17.320000 135.970000 ;
        RECT  1.005000 135.970000 17.250000 136.040000 ;
        RECT  1.005000 136.040000 17.180000 136.110000 ;
        RECT  1.005000 136.110000 17.110000 136.180000 ;
        RECT  1.005000 136.180000 17.040000 136.250000 ;
        RECT  1.005000 136.250000 16.970000 136.320000 ;
        RECT  1.005000 136.320000 16.900000 136.390000 ;
        RECT  1.005000 136.390000 16.830000 136.460000 ;
        RECT  1.005000 136.460000 16.760000 136.530000 ;
        RECT  1.005000 136.530000 16.690000 136.600000 ;
        RECT  1.005000 136.600000 16.620000 136.670000 ;
        RECT  1.005000 136.670000 16.550000 136.740000 ;
        RECT  1.005000 136.740000 16.480000 136.810000 ;
        RECT  1.005000 136.810000 16.410000 136.880000 ;
        RECT  1.005000 136.880000 16.340000 136.950000 ;
        RECT  1.005000 136.950000 16.270000 137.020000 ;
        RECT  1.005000 137.020000 16.200000 137.090000 ;
        RECT  1.005000 137.090000 16.130000 137.160000 ;
        RECT  1.005000 137.160000 16.060000 137.230000 ;
        RECT  1.005000 137.230000 15.990000 137.300000 ;
        RECT  1.005000 137.300000 15.920000 137.370000 ;
        RECT  1.005000 137.370000 15.850000 137.440000 ;
        RECT  1.005000 137.440000 15.780000 137.510000 ;
        RECT  1.005000 137.510000 15.710000 137.580000 ;
        RECT  1.005000 137.580000 15.640000 137.650000 ;
        RECT  1.005000 137.650000 15.570000 137.720000 ;
        RECT  1.005000 137.720000 15.500000 137.790000 ;
        RECT  1.005000 137.790000 15.430000 137.860000 ;
        RECT  1.005000 137.860000 15.360000 137.930000 ;
        RECT  1.005000 137.930000 15.290000 138.000000 ;
        RECT  1.005000 138.000000 15.220000 138.070000 ;
        RECT  1.005000 138.070000 15.150000 138.140000 ;
        RECT  1.005000 138.140000 15.080000 138.210000 ;
        RECT  1.005000 138.210000 15.010000 138.280000 ;
        RECT  1.005000 138.280000 14.940000 138.350000 ;
        RECT  1.005000 138.350000 14.870000 138.420000 ;
        RECT  1.005000 138.420000 14.800000 138.490000 ;
        RECT  1.005000 138.490000 14.730000 138.560000 ;
        RECT  1.005000 138.560000 14.660000 138.630000 ;
        RECT  1.005000 138.630000 14.590000 138.700000 ;
        RECT  1.005000 138.700000 14.520000 138.770000 ;
        RECT  1.005000 138.770000 14.450000 138.840000 ;
        RECT  1.005000 138.840000 14.380000 138.910000 ;
        RECT  1.005000 138.910000 14.310000 138.980000 ;
        RECT  1.005000 138.980000 14.240000 139.050000 ;
        RECT  1.005000 139.050000 14.170000 139.120000 ;
        RECT  1.005000 139.120000 14.120000 139.170000 ;
        RECT  1.005000 139.170000 14.120000 146.215000 ;
        RECT  1.005000 146.215000 14.120000 146.285000 ;
        RECT  1.005000 146.285000 14.190000 146.355000 ;
        RECT  1.005000 146.355000 14.260000 146.425000 ;
        RECT  1.005000 146.425000 14.330000 146.495000 ;
        RECT  1.005000 146.495000 14.400000 146.565000 ;
        RECT  1.005000 146.565000 14.470000 146.635000 ;
        RECT  1.005000 146.635000 14.540000 146.705000 ;
        RECT  1.005000 146.705000 14.610000 146.775000 ;
        RECT  1.005000 146.775000 14.680000 146.845000 ;
        RECT  1.005000 146.845000 14.750000 146.915000 ;
        RECT  1.005000 146.915000 14.820000 146.985000 ;
        RECT  1.005000 146.985000 14.890000 147.055000 ;
        RECT  1.005000 147.055000 14.960000 147.125000 ;
        RECT  1.005000 147.125000 15.030000 147.195000 ;
        RECT  1.005000 147.195000 15.100000 147.265000 ;
        RECT  1.005000 147.265000 15.170000 147.335000 ;
        RECT  1.005000 147.335000 15.240000 147.405000 ;
        RECT  1.005000 147.405000 15.310000 147.475000 ;
        RECT  1.005000 147.475000 15.380000 147.545000 ;
        RECT  1.005000 147.545000 15.450000 147.615000 ;
        RECT  1.005000 147.615000 15.520000 147.685000 ;
        RECT  1.005000 147.685000 15.590000 147.755000 ;
        RECT  1.005000 147.755000 15.660000 147.825000 ;
        RECT  1.005000 147.825000 15.730000 147.895000 ;
        RECT  1.005000 147.895000 15.800000 147.965000 ;
        RECT  1.005000 147.965000 15.870000 148.035000 ;
        RECT  1.005000 148.035000 15.940000 148.105000 ;
        RECT  1.005000 148.105000 16.010000 148.175000 ;
        RECT  1.005000 148.175000 16.080000 148.245000 ;
        RECT  1.005000 148.245000 16.150000 148.315000 ;
        RECT  1.005000 148.315000 16.220000 148.385000 ;
        RECT  1.005000 148.385000 16.290000 148.455000 ;
        RECT  1.005000 148.455000 16.360000 148.525000 ;
        RECT  1.005000 148.525000 16.430000 148.595000 ;
        RECT  1.005000 148.595000 16.500000 148.665000 ;
        RECT  1.005000 148.665000 16.570000 148.735000 ;
        RECT  1.005000 148.735000 16.640000 148.805000 ;
        RECT  1.005000 148.805000 16.710000 148.875000 ;
        RECT  1.005000 148.875000 16.780000 148.945000 ;
        RECT  1.005000 148.945000 16.850000 149.015000 ;
        RECT  1.005000 149.015000 16.920000 149.085000 ;
        RECT  1.005000 149.085000 16.990000 149.155000 ;
        RECT  1.005000 149.155000 17.060000 149.225000 ;
        RECT  1.005000 149.225000 17.130000 149.295000 ;
        RECT  1.005000 149.295000 17.200000 149.365000 ;
        RECT  1.005000 149.365000 17.270000 149.435000 ;
        RECT  1.005000 149.435000 17.340000 149.505000 ;
        RECT  1.005000 149.505000 17.410000 149.575000 ;
        RECT  1.005000 149.575000 17.480000 149.645000 ;
        RECT  1.005000 149.645000 17.550000 149.715000 ;
        RECT  1.005000 149.715000 17.620000 149.780000 ;
        RECT  1.005000 149.780000 56.705000 158.480000 ;
        RECT  1.005000 158.480000 17.650000 158.550000 ;
        RECT  1.005000 158.550000 17.580000 158.620000 ;
        RECT  1.005000 158.620000 17.510000 158.690000 ;
        RECT  1.005000 158.690000 17.440000 158.760000 ;
        RECT  1.005000 158.760000 17.370000 158.830000 ;
        RECT  1.005000 158.830000 17.300000 158.900000 ;
        RECT  1.005000 158.900000 17.230000 158.970000 ;
        RECT  1.005000 158.970000 17.160000 159.040000 ;
        RECT  1.005000 159.040000 17.090000 159.110000 ;
        RECT  1.005000 159.110000 17.020000 159.180000 ;
        RECT  1.005000 159.180000 16.950000 159.250000 ;
        RECT  1.005000 159.250000 16.880000 159.320000 ;
        RECT  1.005000 159.320000 16.810000 159.390000 ;
        RECT  1.005000 159.390000 16.740000 159.460000 ;
        RECT  1.005000 159.460000 16.670000 159.530000 ;
        RECT  1.005000 159.530000 16.600000 159.600000 ;
        RECT  1.005000 159.600000 16.530000 159.670000 ;
        RECT  1.005000 159.670000 16.460000 159.740000 ;
        RECT  1.005000 159.740000 16.390000 159.810000 ;
        RECT  1.005000 159.810000 16.320000 159.880000 ;
        RECT  1.005000 159.880000 16.250000 159.950000 ;
        RECT  1.005000 159.950000 16.180000 160.020000 ;
        RECT  1.005000 160.020000 16.110000 160.090000 ;
        RECT  1.005000 160.090000 16.040000 160.160000 ;
        RECT  1.005000 160.160000 15.970000 160.230000 ;
        RECT  1.005000 160.230000 15.900000 160.300000 ;
        RECT  1.005000 160.300000 15.830000 160.370000 ;
        RECT  1.005000 160.370000 15.760000 160.440000 ;
        RECT  1.005000 160.440000 15.690000 160.510000 ;
        RECT  1.005000 160.510000 15.620000 160.580000 ;
        RECT  1.005000 160.580000 15.550000 160.650000 ;
        RECT  1.005000 160.650000 15.480000 160.720000 ;
        RECT  1.005000 160.720000 15.410000 160.790000 ;
        RECT  1.005000 160.790000 15.340000 160.860000 ;
        RECT  1.005000 160.860000 15.270000 160.930000 ;
        RECT  1.005000 160.930000 15.200000 161.000000 ;
        RECT  1.005000 161.000000 15.130000 161.070000 ;
        RECT  1.005000 161.070000 15.060000 161.140000 ;
        RECT  1.005000 161.140000 14.990000 161.210000 ;
        RECT  1.005000 161.210000 14.920000 161.280000 ;
        RECT  1.005000 161.280000 14.850000 161.350000 ;
        RECT  1.005000 161.350000 14.780000 161.420000 ;
        RECT  1.005000 161.420000 14.710000 161.490000 ;
        RECT  1.005000 161.490000 14.640000 161.560000 ;
        RECT  1.005000 161.560000 14.570000 161.630000 ;
        RECT  1.005000 161.630000 14.500000 161.700000 ;
        RECT  1.005000 161.700000 14.430000 161.770000 ;
        RECT  1.005000 161.770000 14.360000 161.840000 ;
        RECT  1.005000 161.840000 14.290000 161.910000 ;
        RECT  1.005000 161.910000 14.220000 161.980000 ;
        RECT  1.005000 161.980000 14.150000 162.050000 ;
        RECT  1.005000 162.050000 14.120000 162.080000 ;
        RECT  1.005000 162.080000 14.120000 169.220000 ;
        RECT  1.005000 169.220000 14.120000 169.290000 ;
        RECT  1.005000 169.290000 14.190000 169.360000 ;
        RECT  1.005000 169.360000 14.260000 169.430000 ;
        RECT  1.005000 169.430000 14.330000 169.500000 ;
        RECT  1.005000 169.500000 14.400000 169.570000 ;
        RECT  1.005000 169.570000 14.470000 169.640000 ;
        RECT  1.005000 169.640000 14.540000 169.710000 ;
        RECT  1.005000 169.710000 14.610000 169.780000 ;
        RECT  1.005000 169.780000 14.680000 169.850000 ;
        RECT  1.005000 169.850000 14.750000 169.920000 ;
        RECT  1.005000 169.920000 14.820000 169.990000 ;
        RECT  1.005000 169.990000 14.890000 170.060000 ;
        RECT  1.005000 170.060000 14.960000 170.130000 ;
        RECT  1.005000 170.130000 15.030000 170.200000 ;
        RECT  1.005000 170.200000 15.100000 170.270000 ;
        RECT  1.005000 170.270000 15.170000 170.340000 ;
        RECT  1.005000 170.340000 15.240000 170.410000 ;
        RECT  1.005000 170.410000 15.310000 170.480000 ;
        RECT  1.005000 170.480000 15.380000 170.550000 ;
        RECT  1.005000 170.550000 15.450000 170.620000 ;
        RECT  1.005000 170.620000 15.520000 170.690000 ;
        RECT  1.005000 170.690000 15.590000 170.760000 ;
        RECT  1.005000 170.760000 15.660000 170.830000 ;
        RECT  1.005000 170.830000 15.730000 170.900000 ;
        RECT  1.005000 170.900000 15.800000 170.970000 ;
        RECT  1.005000 170.970000 15.870000 171.040000 ;
        RECT  1.005000 171.040000 15.940000 171.110000 ;
        RECT  1.005000 171.110000 16.010000 171.180000 ;
        RECT  1.005000 171.180000 16.080000 171.250000 ;
        RECT  1.005000 171.250000 16.150000 171.320000 ;
        RECT  1.005000 171.320000 16.220000 171.390000 ;
        RECT  1.005000 171.390000 16.290000 171.460000 ;
        RECT  1.005000 171.460000 16.360000 171.530000 ;
        RECT  1.005000 171.530000 16.430000 171.600000 ;
        RECT  1.005000 171.600000 16.500000 171.670000 ;
        RECT  1.005000 171.670000 16.570000 171.740000 ;
        RECT  1.005000 171.740000 16.640000 171.810000 ;
        RECT  1.005000 171.810000 16.710000 171.880000 ;
        RECT  1.005000 171.880000 16.780000 171.950000 ;
        RECT  1.005000 171.950000 16.850000 172.020000 ;
        RECT  1.005000 172.020000 16.920000 172.090000 ;
        RECT  1.005000 172.090000 16.990000 172.160000 ;
        RECT  1.005000 172.160000 17.060000 172.230000 ;
        RECT  1.005000 172.230000 17.130000 172.300000 ;
        RECT  1.005000 172.300000 17.200000 172.370000 ;
        RECT  1.005000 172.370000 17.270000 172.440000 ;
        RECT  1.005000 172.440000 17.340000 172.510000 ;
        RECT  1.005000 172.510000 17.410000 172.580000 ;
        RECT  1.005000 172.580000 17.480000 172.650000 ;
        RECT  1.005000 172.650000 17.550000 172.720000 ;
        RECT  1.005000 172.720000 17.620000 172.780000 ;
        RECT  1.005000 172.780000 57.960000 181.480000 ;
        RECT  1.005000 181.480000 17.625000 181.550000 ;
        RECT  1.005000 181.550000 17.555000 181.620000 ;
        RECT  1.005000 181.620000 17.485000 181.690000 ;
        RECT  1.005000 181.690000 17.415000 181.760000 ;
        RECT  1.005000 181.760000 17.345000 181.830000 ;
        RECT  1.005000 181.830000 17.275000 181.900000 ;
        RECT  1.005000 181.900000 17.205000 181.970000 ;
        RECT  1.005000 181.970000 17.135000 182.040000 ;
        RECT  1.005000 182.040000 17.065000 182.110000 ;
        RECT  1.005000 182.110000 16.995000 182.180000 ;
        RECT  1.005000 182.180000 16.925000 182.250000 ;
        RECT  1.005000 182.250000 16.855000 182.320000 ;
        RECT  1.005000 182.320000 16.785000 182.390000 ;
        RECT  1.005000 182.390000 16.715000 182.460000 ;
        RECT  1.005000 182.460000 16.645000 182.530000 ;
        RECT  1.005000 182.530000 16.575000 182.600000 ;
        RECT  1.005000 182.600000 16.505000 182.670000 ;
        RECT  1.005000 182.670000 16.435000 182.740000 ;
        RECT  1.005000 182.740000 16.365000 182.810000 ;
        RECT  1.005000 182.810000 16.295000 182.880000 ;
        RECT  1.005000 182.880000 16.225000 182.950000 ;
        RECT  1.005000 182.950000 16.155000 183.020000 ;
        RECT  1.005000 183.020000 16.085000 183.090000 ;
        RECT  1.005000 183.090000 16.015000 183.160000 ;
        RECT  1.005000 183.160000 15.945000 183.230000 ;
        RECT  1.005000 183.230000 15.875000 183.300000 ;
        RECT  1.005000 183.300000 15.805000 183.370000 ;
        RECT  1.005000 183.370000 15.735000 183.440000 ;
        RECT  1.005000 183.440000 15.665000 183.510000 ;
        RECT  1.005000 183.510000 15.595000 183.580000 ;
        RECT  1.005000 183.580000 15.525000 183.650000 ;
        RECT  1.005000 183.650000 15.455000 183.720000 ;
        RECT  1.005000 183.720000 15.385000 183.790000 ;
        RECT  1.005000 183.790000 15.315000 183.860000 ;
        RECT  1.005000 183.860000 15.245000 183.930000 ;
        RECT  1.005000 183.930000 15.175000 184.000000 ;
        RECT  1.005000 184.000000 15.105000 184.070000 ;
        RECT  1.005000 184.070000 15.035000 184.140000 ;
        RECT  1.005000 184.140000 14.965000 184.210000 ;
        RECT  1.005000 184.210000 14.895000 184.280000 ;
        RECT  1.005000 184.280000 14.825000 184.350000 ;
        RECT  1.005000 184.350000 14.755000 184.420000 ;
        RECT  1.005000 184.420000 14.685000 184.490000 ;
        RECT  1.005000 184.490000 14.615000 184.560000 ;
        RECT  1.005000 184.560000 14.545000 184.630000 ;
        RECT  1.005000 184.630000 14.475000 184.700000 ;
        RECT  1.005000 184.700000 14.405000 184.770000 ;
        RECT  1.005000 184.770000 14.335000 184.840000 ;
        RECT  1.005000 184.840000 14.265000 184.910000 ;
        RECT  1.005000 184.910000 14.195000 184.980000 ;
        RECT  1.005000 184.980000 14.125000 185.050000 ;
        RECT  1.005000 185.050000 14.120000 185.055000 ;
        RECT  1.005000 185.055000 14.120000 189.585000 ;
        RECT  1.005000 189.585000 14.120000 189.655000 ;
        RECT  1.005000 189.655000 14.190000 189.725000 ;
        RECT  1.005000 189.725000 14.260000 189.795000 ;
        RECT  1.005000 189.795000 14.330000 189.865000 ;
        RECT  1.005000 189.865000 14.400000 189.935000 ;
        RECT  1.005000 189.935000 14.470000 190.005000 ;
        RECT  1.005000 190.005000 14.540000 190.075000 ;
        RECT  1.005000 190.075000 14.610000 190.145000 ;
        RECT  1.005000 190.145000 14.680000 190.215000 ;
        RECT  1.005000 190.215000 14.750000 190.285000 ;
        RECT  1.005000 190.285000 14.820000 190.355000 ;
        RECT  1.005000 190.355000 14.890000 190.425000 ;
        RECT  1.005000 190.425000 14.960000 190.495000 ;
        RECT  1.005000 190.495000 15.030000 190.560000 ;
        RECT  1.005000 190.560000 67.200000 195.075000 ;
        RECT  1.010000  47.125000 14.120000  47.130000 ;
        RECT  1.045000  36.640000 16.180000  36.680000 ;
        RECT  1.050000  47.085000 14.120000  47.125000 ;
        RECT  1.085000  36.680000 16.220000  36.720000 ;
        RECT  1.090000  36.720000 16.260000  36.725000 ;
        RECT  1.090000  36.725000 16.265000  36.795000 ;
        RECT  1.090000  36.795000 16.335000  36.865000 ;
        RECT  1.090000  36.865000 16.405000  36.935000 ;
        RECT  1.090000  36.935000 16.475000  37.005000 ;
        RECT  1.090000  37.005000 16.545000  37.075000 ;
        RECT  1.090000  37.075000 16.615000  37.145000 ;
        RECT  1.090000  37.145000 16.685000  37.215000 ;
        RECT  1.090000  37.215000 16.755000  37.285000 ;
        RECT  1.090000  37.285000 16.825000  37.355000 ;
        RECT  1.090000  37.355000 16.895000  37.425000 ;
        RECT  1.090000  37.425000 16.965000  37.495000 ;
        RECT  1.090000  37.495000 17.035000  37.565000 ;
        RECT  1.090000  37.565000 17.105000  37.635000 ;
        RECT  1.090000  37.635000 17.175000  37.705000 ;
        RECT  1.090000  37.705000 17.245000  37.775000 ;
        RECT  1.090000  37.775000 17.315000  37.845000 ;
        RECT  1.090000  37.845000 17.385000  37.915000 ;
        RECT  1.090000  37.915000 17.455000  37.985000 ;
        RECT  1.090000  37.985000 17.525000  38.055000 ;
        RECT  1.090000  38.055000 17.595000  38.125000 ;
        RECT  1.090000  38.125000 17.665000  38.195000 ;
        RECT  1.090000  38.195000 17.735000  38.265000 ;
        RECT  1.090000  38.265000 17.805000  38.335000 ;
        RECT  1.090000  38.335000 17.875000  38.405000 ;
        RECT  1.090000  38.405000 17.945000  38.475000 ;
        RECT  1.090000  38.475000 18.015000  38.545000 ;
        RECT  1.090000  38.545000 18.085000  38.615000 ;
        RECT  1.090000  38.615000 18.155000  38.685000 ;
        RECT  1.090000  38.685000 18.225000  38.755000 ;
        RECT  1.090000  38.755000 18.295000  38.825000 ;
        RECT  1.090000  38.825000 18.365000  38.895000 ;
        RECT  1.090000  38.895000 18.435000  38.965000 ;
        RECT  1.090000  38.965000 18.505000  39.035000 ;
        RECT  1.090000  39.035000 18.575000  39.105000 ;
        RECT  1.090000  39.105000 18.645000  39.175000 ;
        RECT  1.090000  39.175000 18.715000  39.245000 ;
        RECT  1.090000  39.245000 18.785000  39.315000 ;
        RECT  1.090000  39.315000 18.855000  39.385000 ;
        RECT  1.090000  39.385000 18.925000  39.455000 ;
        RECT  1.090000  39.455000 18.995000  39.525000 ;
        RECT  1.090000  39.525000 19.065000  39.595000 ;
        RECT  1.090000  39.595000 19.135000  39.665000 ;
        RECT  1.090000  39.665000 19.205000  39.735000 ;
        RECT  1.090000  39.735000 19.275000  39.805000 ;
        RECT  1.090000  39.805000 19.345000  39.875000 ;
        RECT  1.090000  39.875000 19.415000  39.945000 ;
        RECT  1.090000  39.945000 19.485000  40.015000 ;
        RECT  1.090000  40.015000 19.555000  40.085000 ;
        RECT  1.090000  40.085000 19.625000  40.155000 ;
        RECT  1.090000  40.155000 19.695000  40.225000 ;
        RECT  1.090000  40.225000 19.765000  40.295000 ;
        RECT  1.090000  40.295000 19.835000  40.350000 ;
        RECT  1.090000  40.350000 56.160000  40.420000 ;
        RECT  1.090000  40.420000 56.090000  40.490000 ;
        RECT  1.090000  40.490000 56.020000  40.560000 ;
        RECT  1.090000  40.560000 55.950000  40.630000 ;
        RECT  1.090000  40.630000 55.880000  40.700000 ;
        RECT  1.090000  40.700000 55.810000  40.770000 ;
        RECT  1.090000  40.770000 55.740000  40.840000 ;
        RECT  1.090000  40.840000 55.670000  40.910000 ;
        RECT  1.090000  40.910000 55.600000  40.980000 ;
        RECT  1.090000  40.980000 55.530000  41.050000 ;
        RECT  1.090000  41.050000 55.460000  41.120000 ;
        RECT  1.090000  41.120000 55.390000  41.190000 ;
        RECT  1.090000  41.190000 55.320000  41.260000 ;
        RECT  1.090000  41.260000 55.250000  41.330000 ;
        RECT  1.090000  41.330000 55.180000  41.400000 ;
        RECT  1.090000  41.400000 55.110000  41.470000 ;
        RECT  1.090000  41.470000 55.040000  41.540000 ;
        RECT  1.090000  41.540000 54.970000  41.610000 ;
        RECT  1.090000  41.610000 54.900000  41.680000 ;
        RECT  1.090000  41.680000 54.830000  41.750000 ;
        RECT  1.090000  41.750000 54.760000  41.820000 ;
        RECT  1.090000  41.820000 54.690000  41.890000 ;
        RECT  1.090000  41.890000 54.620000  41.960000 ;
        RECT  1.090000  41.960000 54.550000  42.030000 ;
        RECT  1.090000  42.030000 54.480000  42.100000 ;
        RECT  1.090000  42.100000 54.410000  42.170000 ;
        RECT  1.090000  42.170000 54.340000  42.240000 ;
        RECT  1.090000  42.240000 54.270000  42.310000 ;
        RECT  1.090000  42.310000 54.200000  42.380000 ;
        RECT  1.090000  42.380000 16.985000  42.450000 ;
        RECT  1.090000  42.450000 16.915000  42.520000 ;
        RECT  1.090000  42.520000 16.845000  42.590000 ;
        RECT  1.090000  42.590000 16.775000  42.660000 ;
        RECT  1.090000  42.660000 16.705000  42.730000 ;
        RECT  1.090000  42.730000 16.635000  42.800000 ;
        RECT  1.090000  42.800000 16.565000  42.870000 ;
        RECT  1.090000  42.870000 16.495000  42.940000 ;
        RECT  1.090000  42.940000 16.425000  43.010000 ;
        RECT  1.090000  43.010000 16.355000  43.080000 ;
        RECT  1.090000  43.080000 16.285000  43.150000 ;
        RECT  1.090000  43.150000 16.215000  43.220000 ;
        RECT  1.090000  43.220000 16.145000  43.290000 ;
        RECT  1.090000  43.290000 16.075000  43.360000 ;
        RECT  1.090000  43.360000 16.005000  43.430000 ;
        RECT  1.090000  43.430000 15.935000  43.500000 ;
        RECT  1.090000  43.500000 15.865000  43.570000 ;
        RECT  1.090000  43.570000 15.795000  43.640000 ;
        RECT  1.090000  43.640000 15.725000  43.710000 ;
        RECT  1.090000  43.710000 15.655000  43.780000 ;
        RECT  1.090000  43.780000 15.585000  43.850000 ;
        RECT  1.090000  43.850000 15.515000  43.920000 ;
        RECT  1.090000  43.920000 15.445000  43.990000 ;
        RECT  1.090000  43.990000 15.375000  44.060000 ;
        RECT  1.090000  44.060000 15.305000  44.130000 ;
        RECT  1.090000  44.130000 15.235000  44.200000 ;
        RECT  1.090000  44.200000 15.165000  44.270000 ;
        RECT  1.090000  44.270000 15.095000  44.340000 ;
        RECT  1.090000  44.340000 15.025000  44.410000 ;
        RECT  1.090000  44.410000 14.955000  44.480000 ;
        RECT  1.090000  44.480000 14.885000  44.550000 ;
        RECT  1.090000  44.550000 14.815000  44.620000 ;
        RECT  1.090000  44.620000 14.745000  44.690000 ;
        RECT  1.090000  44.690000 14.675000  44.760000 ;
        RECT  1.090000  44.760000 14.605000  44.830000 ;
        RECT  1.090000  44.830000 14.535000  44.900000 ;
        RECT  1.090000  44.900000 14.465000  44.970000 ;
        RECT  1.090000  44.970000 14.395000  45.040000 ;
        RECT  1.090000  45.040000 14.325000  45.110000 ;
        RECT  1.090000  45.110000 14.255000  45.180000 ;
        RECT  1.090000  45.180000 14.185000  45.250000 ;
        RECT  1.090000  45.250000 14.120000  45.315000 ;
        RECT  1.090000  45.315000 14.120000  47.045000 ;
        RECT  1.090000  47.045000 14.120000  47.085000 ;
        RECT 52.630000  40.295000 56.230000  40.350000 ;
        RECT 52.700000  40.225000 56.285000  40.295000 ;
        RECT 52.770000  40.155000 56.355000  40.225000 ;
        RECT 52.840000  40.085000 56.425000  40.155000 ;
        RECT 52.910000  40.015000 56.495000  40.085000 ;
        RECT 52.980000  39.945000 56.565000  40.015000 ;
        RECT 53.050000  39.875000 56.635000  39.945000 ;
        RECT 53.120000  39.805000 56.705000  39.875000 ;
        RECT 53.190000  39.735000 56.775000  39.805000 ;
        RECT 53.260000  39.665000 56.845000  39.735000 ;
        RECT 53.270000  39.655000 56.915000  39.665000 ;
        RECT 53.340000  39.585000 56.915000  39.655000 ;
        RECT 53.410000  39.515000 56.915000  39.585000 ;
        RECT 53.480000  39.445000 56.915000  39.515000 ;
        RECT 53.550000  39.375000 56.915000  39.445000 ;
        RECT 53.620000  39.305000 56.915000  39.375000 ;
        RECT 53.690000  39.235000 56.915000  39.305000 ;
        RECT 53.760000  39.165000 56.915000  39.235000 ;
        RECT 53.830000  39.095000 56.915000  39.165000 ;
        RECT 53.900000  39.025000 56.915000  39.095000 ;
        RECT 53.970000  38.955000 56.915000  39.025000 ;
        RECT 54.040000  38.885000 56.915000  38.955000 ;
        RECT 54.110000  38.815000 56.915000  38.885000 ;
        RECT 54.180000  38.745000 56.915000  38.815000 ;
        RECT 54.250000  38.675000 56.915000  38.745000 ;
        RECT 54.320000  38.605000 56.915000  38.675000 ;
        RECT 54.390000  38.535000 56.915000  38.605000 ;
        RECT 54.460000  38.465000 56.915000  38.535000 ;
        RECT 54.530000  38.395000 56.915000  38.465000 ;
        RECT 54.600000  38.325000 56.915000  38.395000 ;
        RECT 54.670000  36.115000 56.915000  38.255000 ;
        RECT 54.670000  38.255000 56.915000  38.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.050000 172.755000 25.010000 195.100000 ;
        RECT 14.055000 172.750000 25.010000 172.755000 ;
        RECT 14.110000 172.695000 25.010000 172.750000 ;
        RECT 14.165000 172.640000 25.010000 172.695000 ;
        RECT 14.300000 172.505000 24.875000 172.640000 ;
        RECT 14.450000 172.355000 24.725000 172.505000 ;
        RECT 14.600000 172.205000 24.575000 172.355000 ;
        RECT 14.750000 172.055000 24.425000 172.205000 ;
        RECT 14.900000 171.905000 24.275000 172.055000 ;
        RECT 15.050000 171.755000 24.125000 171.905000 ;
        RECT 15.200000 171.605000 23.975000 171.755000 ;
        RECT 15.350000 171.455000 23.825000 171.605000 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
        RECT 15.500000 169.130000 21.500000 169.280000 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
        RECT 15.500000 171.230000 23.600000 171.305000 ;
        RECT 15.500000 171.305000 23.675000 171.455000 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
        RECT 17.595000 100.105000 25.925000 100.255000 ;
        RECT 17.745000  99.955000 26.075000 100.105000 ;
        RECT 17.895000  99.805000 26.225000  99.955000 ;
        RECT 18.045000  99.655000 26.375000  99.805000 ;
        RECT 18.195000  99.505000 26.525000  99.655000 ;
        RECT 18.345000  99.355000 26.675000  99.505000 ;
        RECT 18.495000  99.205000 26.825000  99.355000 ;
        RECT 18.645000  99.055000 26.975000  99.205000 ;
        RECT 18.795000  98.905000 27.125000  99.055000 ;
        RECT 18.945000  98.755000 27.275000  98.905000 ;
        RECT 19.095000  98.605000 27.425000  98.755000 ;
        RECT 19.245000  98.455000 27.575000  98.605000 ;
        RECT 19.395000  98.305000 27.725000  98.455000 ;
        RECT 19.545000  98.155000 27.875000  98.305000 ;
        RECT 19.695000  98.005000 28.025000  98.155000 ;
        RECT 19.845000  97.855000 28.175000  98.005000 ;
        RECT 19.995000  97.705000 28.325000  97.855000 ;
        RECT 20.145000  97.555000 28.475000  97.705000 ;
        RECT 20.295000  97.405000 28.625000  97.555000 ;
        RECT 20.445000  97.255000 28.775000  97.405000 ;
        RECT 20.595000  97.105000 28.925000  97.255000 ;
        RECT 20.745000  96.955000 29.075000  97.105000 ;
        RECT 20.895000  96.805000 29.225000  96.955000 ;
        RECT 21.045000  96.655000 29.375000  96.805000 ;
        RECT 21.195000  96.505000 29.525000  96.655000 ;
        RECT 21.345000  96.355000 29.525000  96.505000 ;
        RECT 21.495000  96.205000 29.525000  96.355000 ;
        RECT 21.645000  96.055000 29.525000  96.205000 ;
        RECT 21.795000  95.905000 29.525000  96.055000 ;
        RECT 21.945000  95.755000 29.525000  95.905000 ;
        RECT 22.095000  95.605000 29.525000  95.755000 ;
        RECT 22.245000  95.455000 29.525000  95.605000 ;
        RECT 22.395000  95.305000 29.525000  95.455000 ;
        RECT 22.545000  95.155000 29.525000  95.305000 ;
        RECT 22.695000  95.005000 29.525000  95.155000 ;
        RECT 22.845000  94.855000 29.525000  95.005000 ;
        RECT 22.995000  94.705000 29.525000  94.855000 ;
        RECT 23.145000  94.555000 29.525000  94.705000 ;
        RECT 23.295000  94.405000 29.525000  94.555000 ;
        RECT 23.445000  94.255000 29.525000  94.405000 ;
        RECT 23.595000  94.105000 29.525000  94.255000 ;
        RECT 23.745000  92.540000 29.935000  92.690000 ;
        RECT 23.745000  92.690000 29.785000  92.840000 ;
        RECT 23.745000  92.840000 29.635000  92.990000 ;
        RECT 23.745000  92.990000 29.525000  93.100000 ;
        RECT 23.745000  93.100000 29.525000  93.955000 ;
        RECT 23.745000  93.955000 29.525000  94.105000 ;
        RECT 23.820000  92.465000 30.085000  92.540000 ;
        RECT 23.895000  92.390000 30.160000  92.465000 ;
        RECT 23.945000  92.340000 36.895000  92.390000 ;
        RECT 24.095000  92.190000 36.895000  92.340000 ;
        RECT 24.245000  92.040000 36.895000  92.190000 ;
        RECT 24.395000  91.890000 36.895000  92.040000 ;
        RECT 24.545000  91.740000 36.895000  91.890000 ;
        RECT 24.695000  91.590000 36.895000  91.740000 ;
        RECT 24.845000  91.440000 36.895000  91.590000 ;
        RECT 24.995000  91.290000 36.895000  91.440000 ;
        RECT 25.145000  91.140000 36.895000  91.290000 ;
        RECT 25.295000  90.990000 36.895000  91.140000 ;
        RECT 25.445000  90.840000 36.895000  90.990000 ;
        RECT 25.595000  90.690000 36.895000  90.840000 ;
        RECT 25.745000  90.540000 36.895000  90.690000 ;
        RECT 25.895000   0.000000 36.895000  90.390000 ;
        RECT 25.895000  90.390000 36.895000  90.540000 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
        RECT 25.930000 170.460000 31.930000 170.610000 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
        RECT 25.930000 172.710000 34.180000 172.860000 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
        RECT 25.930000 173.310000 34.780000 173.460000 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
        RECT 25.930000 174.060000 35.530000 174.210000 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
        RECT 25.930000 174.660000 36.130000 174.810000 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
        RECT 25.930000 175.260000 36.730000 175.350000 ;
        RECT 25.930000 175.350000 36.820000 195.100000 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
        RECT 27.975000 100.345000 36.295000 100.495000 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
        RECT 28.425000  99.895000 36.745000 100.045000 ;
        RECT 28.495000  99.825000 36.895000  99.895000 ;
        RECT 28.645000  99.675000 36.895000  99.825000 ;
        RECT 28.795000  99.525000 36.895000  99.675000 ;
        RECT 28.945000  99.375000 36.895000  99.525000 ;
        RECT 29.095000  99.225000 36.895000  99.375000 ;
        RECT 29.245000  99.075000 36.895000  99.225000 ;
        RECT 29.395000  98.925000 36.895000  99.075000 ;
        RECT 29.545000  98.775000 36.895000  98.925000 ;
        RECT 29.695000  98.625000 36.895000  98.775000 ;
        RECT 29.845000  98.475000 36.895000  98.625000 ;
        RECT 29.995000  98.325000 36.895000  98.475000 ;
        RECT 30.145000  98.175000 36.895000  98.325000 ;
        RECT 30.295000  98.025000 36.895000  98.175000 ;
        RECT 30.445000  97.875000 36.895000  98.025000 ;
        RECT 30.595000  97.725000 36.895000  97.875000 ;
        RECT 30.745000  97.575000 36.895000  97.725000 ;
        RECT 30.895000  97.425000 36.895000  97.575000 ;
        RECT 31.045000  97.275000 36.895000  97.425000 ;
        RECT 31.195000  97.125000 36.895000  97.275000 ;
        RECT 31.345000  96.975000 36.895000  97.125000 ;
        RECT 31.385000  92.390000 36.895000  92.540000 ;
        RECT 31.495000  96.825000 36.895000  96.975000 ;
        RECT 31.535000  92.540000 36.895000  92.690000 ;
        RECT 31.645000  96.675000 36.895000  96.825000 ;
        RECT 31.685000  92.690000 36.895000  92.840000 ;
        RECT 31.795000  96.525000 36.895000  96.675000 ;
        RECT 31.835000  92.840000 36.895000  92.990000 ;
        RECT 31.945000  92.990000 36.895000  93.100000 ;
        RECT 31.945000  93.100000 36.895000  96.375000 ;
        RECT 31.945000  96.375000 36.895000  96.525000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  1.145000  43.280000  1.315000  43.810000 ;
      RECT  3.100000  27.160000 48.200000  28.030000 ;
      RECT  3.100000  28.030000  4.020000  38.695000 ;
      RECT  3.100000  38.695000 48.200000  39.565000 ;
      RECT  3.130000  27.140000 48.200000  27.160000 ;
      RECT  3.130000  39.565000 48.200000  39.585000 ;
      RECT  4.735000  29.230000 45.955000  29.430000 ;
      RECT  4.735000  29.430000  4.905000  37.425000 ;
      RECT  4.735000  37.425000 45.955000  37.595000 ;
      RECT  6.115000  33.340000  6.285000  36.490000 ;
      RECT  6.340000  36.970000 45.060000  37.230000 ;
      RECT  6.895000  29.775000  7.065000  32.860000 ;
      RECT  7.675000  33.335000  7.845000  36.490000 ;
      RECT  8.050000  43.270000  8.580000  43.440000 ;
      RECT  8.455000  29.770000  8.625000  32.860000 ;
      RECT  8.510000 162.655000 10.360000 169.150000 ;
      RECT  9.135000  43.505000 70.125000  44.755000 ;
      RECT  9.135000  44.755000 10.385000  71.570000 ;
      RECT  9.135000  71.570000 21.085000  72.820000 ;
      RECT  9.150000 169.400000 10.400000 198.445000 ;
      RECT  9.150000 198.445000 70.125000 199.695000 ;
      RECT  9.170000 133.350000 20.990000 134.540000 ;
      RECT  9.170000 134.540000 10.360000 162.655000 ;
      RECT  9.170000 169.150000 10.360000 169.400000 ;
      RECT  9.200000 133.205000 14.190000 133.350000 ;
      RECT  9.235000  33.340000  9.405000  36.490000 ;
      RECT  9.405000  74.180000  9.935000  74.350000 ;
      RECT 10.015000  29.775000 10.185000  32.860000 ;
      RECT 10.770000 162.655000 11.975000 169.905000 ;
      RECT 10.795000  33.335000 10.965000  36.490000 ;
      RECT 11.100000 170.415000 11.990000 196.835000 ;
      RECT 11.100000 196.835000 68.155000 197.725000 ;
      RECT 11.105000  45.460000 68.155000  46.350000 ;
      RECT 11.105000  46.350000 11.995000  69.975000 ;
      RECT 11.105000  69.975000 22.680000  70.865000 ;
      RECT 11.125000 135.315000 22.660000 136.165000 ;
      RECT 11.125000 136.165000 12.100000 158.915000 ;
      RECT 11.125000 158.915000 11.975000 162.655000 ;
      RECT 11.125000 169.905000 11.975000 170.415000 ;
      RECT 11.575000  29.770000 11.745000  32.860000 ;
      RECT 12.065000   1.000000 70.650000   1.890000 ;
      RECT 12.065000   1.890000 13.045000  22.230000 ;
      RECT 12.065000  22.230000 56.085000  22.350000 ;
      RECT 12.065000  22.350000 56.105000  23.240000 ;
      RECT 12.355000  33.340000 12.525000  36.490000 ;
      RECT 12.400000 159.555000 64.500000 161.990000 ;
      RECT 12.830000 182.570000 66.685000 184.990000 ;
      RECT 13.085000  46.815000 64.500000  46.990000 ;
      RECT 13.085000  46.990000 13.255000  67.965000 ;
      RECT 13.090000  46.740000 64.500000  46.815000 ;
      RECT 13.135000  29.775000 13.305000  32.860000 ;
      RECT 13.915000  33.335000 14.085000  36.490000 ;
      RECT 14.385000  47.160000 15.415000  66.930000 ;
      RECT 14.385000 139.160000 15.415000 158.930000 ;
      RECT 14.385000 162.160000 15.415000 181.930000 ;
      RECT 14.385000 185.160000 15.435000 195.185000 ;
      RECT 14.695000  29.770000 14.865000  32.860000 ;
      RECT 15.475000  33.340000 15.645000  36.490000 ;
      RECT 15.705000  67.340000 64.500000  68.995000 ;
      RECT 15.780000 136.540000 64.500000 138.990000 ;
      RECT 15.780000 159.340000 64.500000 159.555000 ;
      RECT 15.780000 182.340000 66.685000 182.570000 ;
      RECT 15.780000 195.370000 16.490000 195.540000 ;
      RECT 16.255000  29.770000 16.425000  32.860000 ;
      RECT 17.035000  33.335000 17.205000  36.490000 ;
      RECT 17.790000 195.370000 18.500000 195.540000 ;
      RECT 17.815000  29.770000 17.985000  32.860000 ;
      RECT 17.835000 133.145000 20.990000 133.350000 ;
      RECT 18.470000  74.200000 19.000000  74.370000 ;
      RECT 18.595000  33.340000 18.765000  36.490000 ;
      RECT 18.985000  47.515000 19.875000  66.855000 ;
      RECT 18.985000 139.515000 19.875000 158.810000 ;
      RECT 18.985000 162.515000 19.875000 181.810000 ;
      RECT 18.985000 185.515000 19.875000 195.075000 ;
      RECT 19.375000  29.775000 19.545000  32.860000 ;
      RECT 19.565000  97.500000 20.990000 133.145000 ;
      RECT 19.800000  72.820000 21.085000  96.895000 ;
      RECT 19.800000  96.895000 20.990000  97.500000 ;
      RECT 20.155000  33.335000 20.325000  36.490000 ;
      RECT 20.380000 195.370000 21.090000 195.540000 ;
      RECT 20.935000  29.770000 21.105000  32.860000 ;
      RECT 21.715000  33.340000 21.885000  36.490000 ;
      RECT 21.790000  70.865000 22.680000  97.450000 ;
      RECT 21.810000  97.450000 22.660000 135.315000 ;
      RECT 22.390000 195.370000 23.100000 195.540000 ;
      RECT 22.495000  29.775000 22.665000  32.860000 ;
      RECT 23.025000  90.495000 64.500000  92.990000 ;
      RECT 23.055000 113.340000 64.500000 115.990000 ;
      RECT 23.275000  33.335000 23.445000  36.490000 ;
      RECT 23.510000  68.995000 64.500000  69.990000 ;
      RECT 23.585000  47.515000 24.475000  66.810000 ;
      RECT 23.585000  70.160000 24.615000  89.930000 ;
      RECT 23.585000  93.160000 24.615000 112.930000 ;
      RECT 23.585000 116.160000 24.615000 135.930000 ;
      RECT 23.585000 139.515000 24.475000 158.765000 ;
      RECT 23.585000 162.515000 24.475000 181.765000 ;
      RECT 23.585000 185.515000 24.475000 195.030000 ;
      RECT 24.055000  29.770000 24.225000  32.860000 ;
      RECT 24.835000  33.340000 25.005000  36.490000 ;
      RECT 24.980000  90.370000 64.500000  90.495000 ;
      RECT 24.980000 136.370000 64.500000 136.540000 ;
      RECT 24.980000 195.370000 25.690000 195.540000 ;
      RECT 25.615000  29.775000 25.785000  32.860000 ;
      RECT 25.670000  90.340000 64.500000  90.370000 ;
      RECT 25.670000 136.340000 64.500000 136.370000 ;
      RECT 26.395000  33.335000 26.565000  36.490000 ;
      RECT 26.990000 195.370000 27.700000 195.540000 ;
      RECT 27.175000  29.770000 27.345000  32.860000 ;
      RECT 27.955000  33.340000 28.125000  36.490000 ;
      RECT 28.185000  47.515000 29.075000  66.810000 ;
      RECT 28.185000  70.515000 29.075000  89.810000 ;
      RECT 28.185000  93.515000 29.075000 112.855000 ;
      RECT 28.185000 116.515000 29.075000 135.810000 ;
      RECT 28.185000 139.515000 29.075000 158.765000 ;
      RECT 28.185000 162.515000 29.075000 181.765000 ;
      RECT 28.185000 185.515000 29.075000 195.030000 ;
      RECT 28.735000  29.775000 28.905000  32.860000 ;
      RECT 29.515000  33.335000 29.685000  36.490000 ;
      RECT 29.580000 195.370000 30.290000 195.540000 ;
      RECT 30.295000  29.770000 30.465000  32.860000 ;
      RECT 31.075000  33.340000 31.245000  36.490000 ;
      RECT 31.590000 195.370000 32.300000 195.540000 ;
      RECT 31.855000  29.775000 32.025000  32.860000 ;
      RECT 32.635000  33.335000 32.805000  36.490000 ;
      RECT 32.785000  47.515000 33.675000  66.810000 ;
      RECT 32.785000  70.515000 33.675000  89.765000 ;
      RECT 32.785000  93.515000 33.675000 112.810000 ;
      RECT 32.785000 116.515000 33.675000 135.765000 ;
      RECT 32.785000 139.515000 33.675000 158.765000 ;
      RECT 32.785000 162.515000 33.675000 181.765000 ;
      RECT 32.785000 185.515000 33.675000 195.030000 ;
      RECT 33.415000  29.770000 33.585000  32.860000 ;
      RECT 34.180000 195.370000 34.890000 195.540000 ;
      RECT 34.195000  33.340000 34.365000  36.490000 ;
      RECT 34.975000  29.775000 35.145000  32.860000 ;
      RECT 35.755000  33.335000 35.925000  36.490000 ;
      RECT 36.190000 195.370000 36.900000 195.540000 ;
      RECT 36.535000  29.770000 36.705000  32.860000 ;
      RECT 37.315000  33.340000 37.485000  36.490000 ;
      RECT 37.385000  47.515000 38.275000  66.810000 ;
      RECT 37.385000  70.515000 38.275000  89.765000 ;
      RECT 37.385000  93.515000 38.275000 112.810000 ;
      RECT 37.385000 116.515000 38.275000 135.765000 ;
      RECT 37.385000 139.515000 38.275000 158.765000 ;
      RECT 37.385000 162.515000 38.275000 181.765000 ;
      RECT 37.385000 185.515000 38.275000 195.030000 ;
      RECT 38.095000  29.775000 38.265000  32.860000 ;
      RECT 38.780000 195.370000 39.490000 195.540000 ;
      RECT 38.875000  33.335000 39.045000  36.490000 ;
      RECT 39.655000  29.770000 39.825000  32.860000 ;
      RECT 40.435000  33.335000 40.605000  36.490000 ;
      RECT 40.790000 195.370000 41.500000 195.540000 ;
      RECT 41.215000  29.770000 41.385000  32.860000 ;
      RECT 41.985000  47.515000 42.875000  66.810000 ;
      RECT 41.985000  70.515000 42.875000  89.765000 ;
      RECT 41.985000  93.515000 42.875000 112.810000 ;
      RECT 41.985000 116.515000 42.875000 135.765000 ;
      RECT 41.985000 139.515000 42.875000 158.765000 ;
      RECT 41.985000 162.515000 42.875000 181.765000 ;
      RECT 41.985000 185.515000 42.875000 195.030000 ;
      RECT 41.995000  33.340000 42.165000  36.490000 ;
      RECT 42.775000  29.775000 42.945000  32.860000 ;
      RECT 43.380000 195.370000 44.090000 195.540000 ;
      RECT 43.555000  33.335000 43.725000  36.490000 ;
      RECT 44.335000  29.770000 44.505000  32.860000 ;
      RECT 45.115000  33.340000 45.285000  36.490000 ;
      RECT 45.390000 195.370000 46.100000 195.540000 ;
      RECT 45.755000  29.430000 45.955000  37.425000 ;
      RECT 46.585000  47.515000 47.475000  66.810000 ;
      RECT 46.585000  70.515000 47.475000  89.765000 ;
      RECT 46.585000  93.515000 47.475000 112.810000 ;
      RECT 46.585000 116.515000 47.475000 135.765000 ;
      RECT 46.585000 139.515000 47.475000 158.765000 ;
      RECT 46.585000 162.515000 47.475000 181.765000 ;
      RECT 46.585000 185.515000 47.475000 195.030000 ;
      RECT 47.310000  28.030000 48.200000  29.215000 ;
      RECT 47.310000  29.525000 48.200000  38.695000 ;
      RECT 47.330000  29.215000 48.180000  29.525000 ;
      RECT 47.980000 195.370000 48.690000 195.540000 ;
      RECT 49.990000 195.370000 50.700000 195.540000 ;
      RECT 51.185000  47.515000 52.075000  66.810000 ;
      RECT 51.185000  70.515000 52.075000  89.765000 ;
      RECT 51.185000  93.515000 52.075000 112.810000 ;
      RECT 51.185000 116.515000 52.075000 135.765000 ;
      RECT 51.185000 139.515000 52.075000 158.765000 ;
      RECT 51.185000 162.515000 52.075000 181.765000 ;
      RECT 51.185000 185.515000 52.075000 195.030000 ;
      RECT 52.320000  29.300000 68.865000  31.060000 ;
      RECT 52.320000  31.060000 53.210000  41.455000 ;
      RECT 52.320000  41.455000 68.865000  42.495000 ;
      RECT 52.580000 195.370000 53.290000 195.540000 ;
      RECT 53.960000  31.835000 67.140000  32.005000 ;
      RECT 53.960000  32.005000 54.130000  40.410000 ;
      RECT 53.960000  40.410000 67.140000  40.580000 ;
      RECT 54.590000 195.370000 55.300000 195.540000 ;
      RECT 54.695000  36.190000 54.865000  39.290000 ;
      RECT 54.940000  39.770000 66.335000  39.940000 ;
      RECT 55.215000  23.240000 56.105000  28.345000 ;
      RECT 55.215000  28.345000 70.630000  29.300000 ;
      RECT 55.465000  32.620000 55.635000  35.770000 ;
      RECT 55.785000  47.515000 56.675000  66.810000 ;
      RECT 55.785000  70.515000 56.675000  89.765000 ;
      RECT 55.785000  93.515000 56.675000 112.810000 ;
      RECT 55.785000 116.515000 56.675000 135.765000 ;
      RECT 55.785000 139.515000 56.675000 158.765000 ;
      RECT 55.785000 162.515000 56.675000 181.765000 ;
      RECT 55.785000 185.515000 56.675000 195.140000 ;
      RECT 56.255000  36.190000 56.425000  39.290000 ;
      RECT 56.820000  23.480000 57.050000  27.485000 ;
      RECT 56.820000  27.485000 62.810000  27.715000 ;
      RECT 56.850000  21.465000 57.020000  23.480000 ;
      RECT 57.025000  32.620000 57.195000  35.770000 ;
      RECT 57.180000 195.370000 57.890000 195.540000 ;
      RECT 57.555000  23.480000 57.785000  26.430000 ;
      RECT 57.815000  21.735000 61.815000  21.965000 ;
      RECT 57.815000  36.190000 57.985000  39.290000 ;
      RECT 58.585000  32.620000 58.755000  35.770000 ;
      RECT 59.190000 195.370000 59.900000 195.540000 ;
      RECT 59.375000  36.190000 59.545000  39.290000 ;
      RECT 60.145000  32.620000 60.315000  35.770000 ;
      RECT 60.385000  47.515000 61.275000  66.810000 ;
      RECT 60.385000  70.515000 61.275000  89.765000 ;
      RECT 60.385000  93.515000 61.275000 112.810000 ;
      RECT 60.385000 116.515000 61.275000 135.765000 ;
      RECT 60.385000 139.515000 61.275000 158.765000 ;
      RECT 60.385000 162.515000 61.275000 181.765000 ;
      RECT 60.385000 185.515000 61.275000 195.140000 ;
      RECT 60.935000  36.190000 61.105000  39.290000 ;
      RECT 61.705000  32.620000 61.875000  35.770000 ;
      RECT 61.780000 195.370000 62.490000 195.540000 ;
      RECT 61.850000  23.480000 62.080000  26.430000 ;
      RECT 62.495000  36.190000 62.665000  39.290000 ;
      RECT 62.580000  23.480000 62.810000  27.485000 ;
      RECT 62.610000  21.465000 62.780000  23.480000 ;
      RECT 63.265000  32.620000 63.435000  35.770000 ;
      RECT 63.790000 195.370000 64.500000 195.540000 ;
      RECT 64.055000  36.190000 64.225000  39.290000 ;
      RECT 64.825000  32.620000 64.995000  35.770000 ;
      RECT 64.845000  47.160000 65.875000  66.930000 ;
      RECT 64.845000  70.160000 65.875000  72.950000 ;
      RECT 64.845000  87.140000 65.875000  89.930000 ;
      RECT 64.845000  93.160000 65.875000  95.950000 ;
      RECT 64.845000 110.145000 65.875000 112.935000 ;
      RECT 64.845000 116.160000 65.875000 118.950000 ;
      RECT 64.845000 133.140000 65.875000 135.930000 ;
      RECT 64.845000 139.160000 65.875000 158.930000 ;
      RECT 64.845000 162.160000 65.875000 181.930000 ;
      RECT 64.845000 185.160000 65.875000 195.180000 ;
      RECT 64.985000  72.950000 65.875000  87.140000 ;
      RECT 64.985000  95.950000 65.875000 110.145000 ;
      RECT 64.985000 118.950000 65.875000 133.140000 ;
      RECT 65.615000  36.190000 65.785000  39.290000 ;
      RECT 66.385000  32.620000 66.555000  35.770000 ;
      RECT 66.935000  32.005000 67.140000  36.065000 ;
      RECT 66.935000  36.275000 67.140000  40.410000 ;
      RECT 66.970000  36.065000 67.140000  36.275000 ;
      RECT 67.265000  46.350000 68.155000 101.315000 ;
      RECT 67.265000 166.045000 68.155000 196.835000 ;
      RECT 67.290000 101.315000 68.140000 101.710000 ;
      RECT 67.290000 101.710000 68.155000 165.645000 ;
      RECT 67.290000 165.645000 68.140000 166.045000 ;
      RECT 67.975000  31.060000 68.865000  40.480000 ;
      RECT 67.975000  41.315000 68.865000  41.455000 ;
      RECT 68.000000  40.480000 68.830000  41.315000 ;
      RECT 68.875000  44.755000 70.125000  45.995000 ;
      RECT 68.875000  46.185000 70.125000 198.445000 ;
      RECT 68.905000  45.995000 70.095000  46.185000 ;
      RECT 69.740000  22.520000 70.630000  28.345000 ;
      RECT 69.760000   1.890000 70.650000   2.770000 ;
      RECT 69.765000   3.845000 70.630000   8.915000 ;
      RECT 69.765000   9.845000 70.630000  14.915000 ;
      RECT 69.765000  16.165000 70.630000  21.235000 ;
      RECT 69.780000   2.770000 70.630000   3.845000 ;
      RECT 69.780000   8.915000 70.630000   9.845000 ;
      RECT 69.780000  14.915000 70.630000  16.165000 ;
      RECT 69.780000  21.235000 70.630000  22.520000 ;
      RECT 70.470000  42.820000 71.055000  42.990000 ;
      RECT 70.725000  42.735000 71.055000  42.820000 ;
      RECT 72.245000 199.210000 72.775000 199.380000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   2.170000  0.215000   2.240000 ;
      RECT  0.000000   2.170000  0.725000   2.680000 ;
      RECT  0.000000   2.240000  0.285000   2.310000 ;
      RECT  0.000000   2.310000  0.355000   2.380000 ;
      RECT  0.000000   2.380000  0.425000   2.450000 ;
      RECT  0.000000   2.450000  0.495000   2.520000 ;
      RECT  0.000000   2.520000  0.565000   2.590000 ;
      RECT  0.000000   2.590000  0.635000   2.660000 ;
      RECT  0.000000   2.660000  0.705000   2.680000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000  36.755000  0.725000  36.800000 ;
      RECT  0.000000  36.755000  0.810000  36.840000 ;
      RECT  0.000000  36.800000  0.770000  36.840000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  46.930000  0.725000  47.015000 ;
      RECT  0.000000  46.930000  0.770000  46.970000 ;
      RECT  0.000000  46.970000  0.730000  47.010000 ;
      RECT  0.000000  47.010000  0.725000  47.015000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000 195.355000 67.480000 200.000000 ;
      RECT  0.000000 195.355000 75.000000 200.000000 ;
      RECT 14.400000  45.430000 57.415000  47.315000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.175000 16.525000  54.100000 ;
      RECT 14.400000  47.315000 16.665000  54.100000 ;
      RECT 14.400000  54.100000 16.665000  54.905000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.445000  70.315000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.175000 24.540000  72.870000 ;
      RECT 14.400000  70.315000 24.680000  72.925000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.925000 23.590000  74.015000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.875000 18.130000  74.695000 ;
      RECT 14.400000  74.015000 18.270000  74.555000 ;
      RECT 14.400000  74.555000 24.680000  75.675000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.680000  77.125000 ;
      RECT 14.400000  75.730000 24.540000  77.125000 ;
      RECT 14.400000  77.125000 24.680000  79.295000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.505000  93.315000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.175000 24.540000 100.125000 ;
      RECT 14.400000  93.315000 24.680000 100.125000 ;
      RECT 14.400000 100.125000 24.680000 102.295000 ;
      RECT 14.400000 116.180000 24.540000 123.030000 ;
      RECT 14.400000 116.180000 57.415000 116.315000 ;
      RECT 14.400000 116.315000 24.680000 123.030000 ;
      RECT 14.400000 123.030000 24.680000 125.295000 ;
      RECT 14.400000 139.285000 16.525000 146.100000 ;
      RECT 14.400000 139.285000 57.450000 139.315000 ;
      RECT 14.400000 139.315000 16.665000 146.100000 ;
      RECT 14.400000 146.100000 16.665000 146.770000 ;
      RECT 14.400000 162.195000 16.525000 169.105000 ;
      RECT 14.400000 162.195000 57.465000 162.315000 ;
      RECT 14.400000 162.315000 16.665000 169.105000 ;
      RECT 14.400000 169.105000 16.665000 171.295000 ;
      RECT 14.400000 185.170000 15.340000 189.470000 ;
      RECT 14.400000 185.170000 15.480000 189.470000 ;
      RECT 14.400000 189.470000 15.480000 190.155000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.410000 162.185000 16.525000 162.195000 ;
      RECT 14.415000 185.155000 15.340000 185.170000 ;
      RECT 14.415000 185.155000 15.480000 185.170000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000 162.175000 16.525000 162.185000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000 139.230000 16.525000 139.285000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.470000  54.100000 16.525000  54.170000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 146.100000 16.525000 146.170000 ;
      RECT 14.470000 169.105000 16.525000 169.175000 ;
      RECT 14.470000 189.470000 15.340000 189.540000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.485000 185.085000 15.340000 185.155000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.510000 139.175000 16.525000 139.230000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.540000  54.170000 16.525000  54.240000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 146.170000 16.525000 146.240000 ;
      RECT 14.540000 169.175000 16.525000 169.245000 ;
      RECT 14.540000 189.540000 15.340000 189.610000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.555000 185.015000 15.340000 185.085000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 185.005000 58.580000 185.015000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.610000  54.240000 16.525000  54.310000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 146.240000 16.525000 146.310000 ;
      RECT 14.610000 169.245000 16.525000 169.315000 ;
      RECT 14.610000 189.610000 15.340000 189.680000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 184.935000 58.590000 185.005000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.680000  54.310000 16.525000  54.380000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 146.310000 16.525000 146.380000 ;
      RECT 14.680000 169.315000 16.525000 169.385000 ;
      RECT 14.680000 189.680000 15.340000 189.750000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 184.865000 58.660000 184.935000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.750000  54.380000 16.525000  54.450000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 146.380000 16.525000 146.450000 ;
      RECT 14.750000 169.385000 16.525000 169.455000 ;
      RECT 14.750000 189.750000 15.340000 189.820000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 184.795000 58.730000 184.865000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.820000  54.450000 16.525000  54.520000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 146.450000 16.525000 146.520000 ;
      RECT 14.820000 169.455000 16.525000 169.525000 ;
      RECT 14.820000 189.820000 15.340000 189.890000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 184.725000 58.800000 184.795000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.890000  54.520000 16.525000  54.590000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 146.520000 16.525000 146.590000 ;
      RECT 14.890000 169.525000 16.525000 169.595000 ;
      RECT 14.890000 189.890000 15.340000 189.960000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 184.655000 58.870000 184.725000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.960000  54.590000 16.525000  54.660000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 146.590000 16.525000 146.660000 ;
      RECT 14.960000 169.595000 16.525000 169.665000 ;
      RECT 14.960000 189.960000 15.340000 190.030000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 184.585000 58.940000 184.655000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.030000  54.660000 16.525000  54.730000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 146.660000 16.525000 146.730000 ;
      RECT 15.030000 169.665000 16.525000 169.735000 ;
      RECT 15.030000 190.030000 15.340000 190.100000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 184.515000 59.010000 184.585000 ;
      RECT 15.070000 146.770000 18.190000 148.295000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000 190.155000 75.000000 190.280000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.100000  54.730000 16.525000  54.800000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 146.730000 16.525000 146.800000 ;
      RECT 15.100000 169.735000 16.525000 169.805000 ;
      RECT 15.100000 190.100000 15.340000 190.170000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 146.800000 16.525000 146.825000 ;
      RECT 15.125000 184.445000 59.080000 184.515000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.170000  54.800000 16.525000  54.870000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 169.805000 16.525000 169.875000 ;
      RECT 15.170000 190.170000 15.340000 190.240000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 146.825000 16.525000 146.895000 ;
      RECT 15.195000 184.375000 59.150000 184.445000 ;
      RECT 15.205000  54.905000 18.790000  56.295000 ;
      RECT 15.210000 190.240000 15.340000 190.280000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.240000  54.870000 16.525000  54.940000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 169.875000 16.525000 169.945000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 146.895000 16.595000 146.965000 ;
      RECT 15.265000 184.305000 59.220000 184.375000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.310000  54.940000 16.525000  55.010000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 169.945000 16.525000 170.015000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 146.965000 16.665000 147.035000 ;
      RECT 15.335000 184.235000 59.290000 184.305000 ;
      RECT 15.345000  55.010000 16.525000  55.045000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 170.015000 16.525000 170.085000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 147.035000 16.735000 147.105000 ;
      RECT 15.405000 184.165000 59.360000 184.235000 ;
      RECT 15.415000  55.045000 17.345000  55.115000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 170.085000 16.525000 170.155000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 147.105000 16.805000 147.175000 ;
      RECT 15.475000 184.095000 59.430000 184.165000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 60.970000  31.015000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  31.015000 60.970000  35.550000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.070000 60.830000  35.550000 ;
      RECT 15.485000  35.550000 60.970000  35.975000 ;
      RECT 15.485000  55.115000 17.415000  55.185000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 170.155000 16.525000 170.225000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 147.175000 16.875000 147.245000 ;
      RECT 15.545000 184.025000 59.500000 184.095000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  55.185000 17.485000  55.255000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 170.225000 16.525000 170.295000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 147.245000 16.945000 147.315000 ;
      RECT 15.615000 183.955000 59.570000 184.025000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  55.255000 17.555000  55.325000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 170.295000 16.525000 170.365000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 147.315000 17.015000 147.385000 ;
      RECT 15.685000 183.885000 59.640000 183.955000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  55.325000 17.625000  55.395000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 170.365000 16.525000 170.435000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 147.385000 17.085000 147.455000 ;
      RECT 15.755000 183.815000 59.710000 183.885000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  55.395000 17.695000  55.465000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 170.435000 16.525000 170.505000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 147.455000 17.155000 147.525000 ;
      RECT 15.825000 183.745000 59.780000 183.815000 ;
      RECT 15.835000  55.465000 17.765000  55.535000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 170.505000 16.525000 170.575000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 147.525000 17.225000 147.595000 ;
      RECT 15.895000 183.675000 59.850000 183.745000 ;
      RECT 15.905000  55.535000 17.835000  55.605000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.975000 54.530000  38.195000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 170.575000 16.525000 170.645000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 147.595000 17.295000 147.665000 ;
      RECT 15.965000 183.605000 59.920000 183.675000 ;
      RECT 15.975000  55.605000 17.905000  55.675000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 170.645000 16.525000 170.715000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 147.665000 17.365000 147.735000 ;
      RECT 16.035000 183.535000 59.990000 183.605000 ;
      RECT 16.045000  55.675000 17.975000  55.745000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.070000  43.760000 59.300000  45.430000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 170.715000 16.525000 170.785000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 147.735000 17.435000 147.805000 ;
      RECT 16.105000 183.465000 60.060000 183.535000 ;
      RECT 16.115000  55.745000 18.045000  55.815000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 170.785000 16.525000 170.855000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 147.805000 17.505000 147.875000 ;
      RECT 16.175000 183.395000 60.130000 183.465000 ;
      RECT 16.185000  55.815000 18.115000  55.885000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 170.855000 16.525000 170.925000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 147.875000 17.575000 147.945000 ;
      RECT 16.245000 183.325000 60.200000 183.395000 ;
      RECT 16.255000  55.885000 18.185000  55.955000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 170.925000 16.525000 170.995000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 147.945000 17.645000 148.015000 ;
      RECT 16.315000 183.255000 60.270000 183.325000 ;
      RECT 16.325000  55.955000 18.255000  56.025000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 170.995000 16.525000 171.065000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 148.015000 17.715000 148.085000 ;
      RECT 16.385000 183.185000 60.340000 183.255000 ;
      RECT 16.395000  56.025000 18.325000  56.095000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 171.065000 16.525000 171.135000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 148.085000 17.785000 148.155000 ;
      RECT 16.455000 183.115000 60.410000 183.185000 ;
      RECT 16.465000  56.095000 18.395000  56.165000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 171.135000 16.525000 171.205000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 148.155000 17.855000 148.225000 ;
      RECT 16.525000 183.045000 60.480000 183.115000 ;
      RECT 16.535000  56.165000 18.465000  56.235000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.295000 58.700000  80.500000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.295000 58.700000 103.500000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000 171.295000 58.710000 172.500000 ;
      RECT 16.595000  56.295000 58.670000  57.500000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 148.225000 17.925000 148.295000 ;
      RECT 16.595000 148.295000 58.630000 149.500000 ;
      RECT 16.595000 182.975000 60.550000 183.045000 ;
      RECT 16.605000  56.235000 18.535000  56.305000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.665000 125.295000 58.700000 126.500000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 148.295000 17.995000 148.365000 ;
      RECT 16.665000 182.905000 60.620000 182.975000 ;
      RECT 16.675000  56.305000 18.605000  56.375000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.735000  56.375000 18.675000  56.435000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 148.365000 18.065000 148.435000 ;
      RECT 16.735000 182.835000 60.690000 182.905000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000 182.820000 58.635000 185.155000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 57.440000  79.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 57.440000 102.505000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000 171.435000 57.450000 171.505000 ;
      RECT 16.805000  56.435000 57.410000  56.505000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 148.435000 57.370000 148.505000 ;
      RECT 16.805000 182.765000 60.760000 182.835000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.830000 182.740000 60.830000 182.765000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 57.510000  79.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 57.510000 102.575000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000 171.505000 57.520000 171.575000 ;
      RECT 16.875000  56.505000 57.480000  56.575000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 57.440000 125.505000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 148.505000 57.440000 148.575000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.900000 182.670000 60.830000 182.740000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 57.580000  79.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 57.580000 102.645000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000 171.575000 57.590000 171.645000 ;
      RECT 16.945000  56.575000 57.550000  56.645000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 57.510000 125.575000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 148.575000 57.510000 148.645000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.970000 182.600000 60.830000 182.670000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 57.650000  79.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 57.650000 102.715000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000 171.645000 57.660000 171.715000 ;
      RECT 17.015000  56.645000 57.620000  56.715000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 57.580000 125.645000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 148.645000 57.580000 148.715000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.040000 182.530000 60.830000 182.600000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 57.720000  79.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 57.720000 102.785000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000 171.715000 57.730000 171.785000 ;
      RECT 17.085000  56.715000 57.690000  56.785000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 57.650000 125.715000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 148.715000 57.650000 148.785000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.110000 182.460000 60.830000 182.530000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 57.790000  79.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 57.790000 102.855000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000 171.785000 57.800000 171.855000 ;
      RECT 17.155000  56.785000 57.760000  56.855000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 57.720000 125.785000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 148.785000 57.720000 148.855000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.970000  43.760000 ;
      RECT 17.180000 182.390000 60.830000 182.460000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 57.860000  79.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 57.860000 102.925000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000 171.855000 57.870000 171.925000 ;
      RECT 17.225000  56.855000 57.830000  56.925000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 57.790000 125.855000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 148.855000 57.790000 148.925000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.250000 182.320000 60.830000 182.390000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 57.930000  79.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 57.930000 102.995000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000 171.925000 57.940000 171.995000 ;
      RECT 17.295000  56.925000 57.900000  56.995000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 57.860000 125.925000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 148.925000 57.860000 148.995000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.320000 182.250000 60.830000 182.320000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 58.000000  80.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 58.000000 103.065000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000 171.995000 58.010000 172.065000 ;
      RECT 17.365000  56.995000 57.970000  57.065000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 57.930000 125.995000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 148.995000 57.930000 149.065000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.390000 182.180000 60.830000 182.250000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 58.070000  80.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 58.070000 103.135000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000 172.065000 58.080000 172.135000 ;
      RECT 17.435000  57.065000 58.040000  57.135000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 58.000000 126.065000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 149.065000 58.000000 149.135000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.460000 182.110000 60.830000 182.180000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 58.140000  80.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 58.140000 103.205000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000 172.135000 58.150000 172.205000 ;
      RECT 17.505000  57.135000 58.110000  57.205000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 58.070000 126.135000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 149.135000 58.070000 149.205000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.530000 182.040000 60.830000 182.110000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 58.210000  80.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 58.210000 103.275000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000 172.205000 58.220000 172.275000 ;
      RECT 17.575000  57.205000 58.180000  57.275000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 58.140000 126.205000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 149.205000 58.140000 149.275000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.600000 181.970000 60.830000 182.040000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 58.280000  80.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 58.280000 103.345000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000 172.275000 58.290000 172.345000 ;
      RECT 17.645000  57.275000 58.250000  57.345000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 58.210000 126.275000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 149.275000 58.210000 149.345000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.670000 181.900000 60.830000 181.970000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 58.350000  80.415000 ;
      RECT 17.690000  89.850000 57.680000  93.140000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 58.350000 103.415000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000 172.345000 58.360000 172.415000 ;
      RECT 17.715000  57.345000 58.320000  57.415000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 58.280000 126.345000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 149.345000 58.280000 149.415000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.740000 181.830000 60.830000 181.900000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.750000  66.790000 57.620000  70.140000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 58.420000  80.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 58.420000 103.485000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 58.490000  80.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 58.490000 103.500000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.970000  66.790000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.970000  89.850000 ;
      RECT 17.780000 172.415000 58.430000 172.485000 ;
      RECT 17.785000  57.415000 58.390000  57.485000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 58.350000 126.415000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 149.415000 58.350000 149.485000 ;
      RECT 17.785000 158.810000 57.585000 162.195000 ;
      RECT 17.795000 172.485000 58.500000 172.500000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  57.485000 58.460000  57.500000 ;
      RECT 17.800000 149.485000 58.420000 149.500000 ;
      RECT 17.810000 181.760000 60.830000 181.830000 ;
      RECT 17.810000 181.760000 60.970000 182.820000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.820000 112.760000 57.550000 116.180000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.970000 112.760000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.970000 158.810000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 58.420000 126.485000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 58.490000 126.500000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.890000 135.795000 57.480000 139.285000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.970000 135.795000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.130000  38.195000 52.655000  40.070000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 59.390000  29.430000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.400000  40.070000 52.515000  40.210000 ;
      RECT 22.850000  42.520000 60.970000  42.660000 ;
      RECT 24.675000   0.000000 25.615000   0.815000 ;
      RECT 24.675000   0.000000 25.755000   0.675000 ;
      RECT 24.675000   0.675000 50.250000   8.480000 ;
      RECT 24.675000   0.815000 50.110000   8.480000 ;
      RECT 24.675000   8.480000 50.250000   8.565000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.765000   8.565000 46.695000  12.120000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 28.035000   0.000000 50.250000   0.675000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.175000   0.000000 50.110000   0.815000 ;
      RECT 28.175000   0.000000 50.110000   8.480000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 37.175000  12.120000 37.610000  25.940000 ;
      RECT 37.175000  12.120000 46.660000  12.155000 ;
      RECT 37.175000  12.155000 37.750000  25.800000 ;
      RECT 37.175000  25.800000 55.935000  25.980000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 60.970000  82.770000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.770000 60.970000  89.760000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.825000 60.830000  89.760000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 60.970000 105.770000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.770000 60.970000 112.760000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.825000 60.830000 112.705000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 60.970000 128.770000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.770000 60.970000 135.760000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.825000 60.830000 135.740000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 60.970000 151.840000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.840000 60.970000 158.760000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.895000 60.830000 158.755000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 60.970000  59.800000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.800000 60.970000  66.760000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.855000 60.830000  66.735000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 57.055000  35.975000 60.970000  39.725000 ;
      RECT 57.055000  39.725000 60.970000  42.520000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.195000  35.835000 60.830000  39.780000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 58.240000 172.500000 58.515000 172.570000 ;
      RECT 58.240000 172.500000 60.970000 174.760000 ;
      RECT 58.240000 172.570000 58.585000 172.640000 ;
      RECT 58.240000 172.640000 58.655000 172.710000 ;
      RECT 58.240000 172.710000 58.725000 172.780000 ;
      RECT 58.240000 172.780000 58.795000 172.850000 ;
      RECT 58.240000 172.850000 58.865000 172.920000 ;
      RECT 58.240000 172.920000 58.935000 172.990000 ;
      RECT 58.240000 172.990000 59.005000 173.060000 ;
      RECT 58.240000 173.060000 59.075000 173.130000 ;
      RECT 58.240000 173.130000 59.145000 173.200000 ;
      RECT 58.240000 173.200000 59.215000 173.270000 ;
      RECT 58.240000 173.270000 59.285000 173.340000 ;
      RECT 58.240000 173.340000 59.355000 173.410000 ;
      RECT 58.240000 173.410000 59.425000 173.480000 ;
      RECT 58.240000 173.480000 59.495000 173.550000 ;
      RECT 58.240000 173.550000 59.565000 173.620000 ;
      RECT 58.240000 173.620000 59.635000 173.690000 ;
      RECT 58.240000 173.690000 59.705000 173.760000 ;
      RECT 58.240000 173.760000 59.775000 173.830000 ;
      RECT 58.240000 173.830000 59.845000 173.900000 ;
      RECT 58.240000 173.900000 59.915000 173.970000 ;
      RECT 58.240000 173.970000 59.985000 174.040000 ;
      RECT 58.240000 174.040000 60.055000 174.110000 ;
      RECT 58.240000 174.110000 60.125000 174.180000 ;
      RECT 58.240000 174.180000 60.195000 174.250000 ;
      RECT 58.240000 174.250000 60.265000 174.320000 ;
      RECT 58.240000 174.320000 60.335000 174.390000 ;
      RECT 58.240000 174.390000 60.405000 174.460000 ;
      RECT 58.240000 174.460000 60.475000 174.530000 ;
      RECT 58.240000 174.530000 60.545000 174.600000 ;
      RECT 58.240000 174.600000 60.615000 174.670000 ;
      RECT 58.240000 174.670000 60.685000 174.740000 ;
      RECT 58.240000 174.740000 60.755000 174.810000 ;
      RECT 58.240000 174.760000 60.970000 181.760000 ;
      RECT 58.240000 174.810000 60.825000 174.815000 ;
      RECT 58.240000 174.815000 60.830000 181.760000 ;
      RECT 67.480000 190.280000 75.000000 195.355000 ;
      RECT 67.480000 190.295000 75.000000 200.000000 ;
      RECT 70.480000 193.295000 72.000000 197.000000 ;
      RECT 74.430000   0.000000 75.000000 190.155000 ;
      RECT 74.570000   0.000000 75.000000 190.295000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.195000  36.635000 ;
      RECT  0.000000  36.635000  0.670000  37.110000 ;
      RECT  0.000000  36.730000  0.150000  36.880000 ;
      RECT  0.000000  36.880000  0.300000  37.030000 ;
      RECT  0.000000  37.030000  0.450000  37.150000 ;
      RECT  0.000000  37.110000  0.670000  46.360000 ;
      RECT  0.000000  37.150000  0.570000  46.320000 ;
      RECT  0.000000  46.320000  0.420000  46.470000 ;
      RECT  0.000000  46.360000  0.195000  46.835000 ;
      RECT  0.000000  46.470000  0.270000  46.620000 ;
      RECT  0.000000  46.620000  0.120000  46.770000 ;
      RECT  0.000000  46.835000  0.195000 173.455000 ;
      RECT  0.000000 173.455000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT 13.800000 101.520000 15.100000 102.035000 ;
      RECT 13.800000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 101.560000 15.425000 101.710000 ;
      RECT 13.900000 101.710000 15.275000 101.860000 ;
      RECT 13.900000 101.860000 15.125000 102.010000 ;
      RECT 13.900000 102.010000 15.100000 102.035000 ;
      RECT 13.900000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 171.140000 14.950000 171.290000 ;
      RECT 13.900000 171.290000 14.800000 171.440000 ;
      RECT 13.900000 171.440000 14.650000 171.590000 ;
      RECT 13.900000 171.590000 14.500000 171.740000 ;
      RECT 13.900000 171.740000 14.350000 171.890000 ;
      RECT 13.900000 171.890000 14.200000 172.040000 ;
      RECT 13.900000 172.040000 14.050000 172.190000 ;
      RECT 14.020000 101.440000 15.575000 101.560000 ;
      RECT 14.170000 101.290000 15.695000 101.440000 ;
      RECT 14.320000 101.140000 15.845000 101.290000 ;
      RECT 14.470000 100.990000 15.995000 101.140000 ;
      RECT 14.620000 100.840000 16.145000 100.990000 ;
      RECT 14.770000 100.690000 16.295000 100.840000 ;
      RECT 14.920000 100.540000 16.445000 100.690000 ;
      RECT 15.070000 100.390000 16.595000 100.540000 ;
      RECT 15.220000 100.240000 16.745000 100.390000 ;
      RECT 15.370000 100.090000 16.895000 100.240000 ;
      RECT 15.520000  99.940000 17.045000 100.090000 ;
      RECT 15.670000  99.790000 17.195000  99.940000 ;
      RECT 15.820000  99.640000 17.345000  99.790000 ;
      RECT 15.970000  99.490000 17.495000  99.640000 ;
      RECT 16.120000  99.340000 17.645000  99.490000 ;
      RECT 16.270000  99.190000 17.795000  99.340000 ;
      RECT 16.420000  99.040000 17.945000  99.190000 ;
      RECT 16.570000  98.890000 18.095000  99.040000 ;
      RECT 16.720000  98.740000 18.245000  98.890000 ;
      RECT 16.870000  98.590000 18.395000  98.740000 ;
      RECT 17.020000  98.440000 18.545000  98.590000 ;
      RECT 17.170000  98.290000 18.695000  98.440000 ;
      RECT 17.320000  98.140000 18.845000  98.290000 ;
      RECT 17.470000  97.990000 18.995000  98.140000 ;
      RECT 17.620000  97.840000 19.145000  97.990000 ;
      RECT 17.770000  97.690000 19.295000  97.840000 ;
      RECT 17.920000  97.540000 19.445000  97.690000 ;
      RECT 18.070000  97.390000 19.595000  97.540000 ;
      RECT 18.220000  97.240000 19.745000  97.390000 ;
      RECT 18.370000  97.090000 19.895000  97.240000 ;
      RECT 18.520000  96.940000 20.045000  97.090000 ;
      RECT 18.670000  96.790000 20.195000  96.940000 ;
      RECT 18.820000  96.640000 20.345000  96.790000 ;
      RECT 18.970000  96.490000 20.495000  96.640000 ;
      RECT 19.120000  96.340000 20.645000  96.490000 ;
      RECT 19.270000  96.190000 20.795000  96.340000 ;
      RECT 19.420000  96.040000 20.945000  96.190000 ;
      RECT 19.570000  95.890000 21.095000  96.040000 ;
      RECT 19.720000  95.740000 21.245000  95.890000 ;
      RECT 19.870000  95.590000 21.395000  95.740000 ;
      RECT 20.020000  95.440000 21.545000  95.590000 ;
      RECT 20.170000  95.290000 21.695000  95.440000 ;
      RECT 20.320000  95.140000 21.845000  95.290000 ;
      RECT 20.470000  94.990000 21.995000  95.140000 ;
      RECT 20.620000  94.840000 22.145000  94.990000 ;
      RECT 20.770000  94.690000 22.295000  94.840000 ;
      RECT 20.920000  94.540000 22.445000  94.690000 ;
      RECT 21.070000  94.390000 22.595000  94.540000 ;
      RECT 21.220000  94.240000 22.745000  94.390000 ;
      RECT 21.370000  94.090000 22.895000  94.240000 ;
      RECT 21.520000  93.940000 23.045000  94.090000 ;
      RECT 21.670000  93.790000 23.195000  93.940000 ;
      RECT 21.695000  93.765000 23.345000  93.790000 ;
      RECT 21.845000  93.615000 23.345000  93.765000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 168.965000 25.530000 172.475000 ;
      RECT 21.970000 104.775000 25.530000 104.845000 ;
      RECT 21.995000  93.465000 23.345000  93.615000 ;
      RECT 22.050000 168.965000 25.530000 169.115000 ;
      RECT 22.120000 104.625000 25.530000 104.775000 ;
      RECT 22.145000  93.315000 23.345000  93.465000 ;
      RECT 22.200000 169.115000 25.530000 169.265000 ;
      RECT 22.270000 104.475000 25.530000 104.625000 ;
      RECT 22.295000  93.165000 23.345000  93.315000 ;
      RECT 22.350000 169.265000 25.530000 169.415000 ;
      RECT 22.420000 104.325000 25.530000 104.475000 ;
      RECT 22.445000  93.015000 23.345000  93.165000 ;
      RECT 22.500000 169.415000 25.530000 169.565000 ;
      RECT 22.570000 104.175000 25.530000 104.325000 ;
      RECT 22.595000  92.865000 23.345000  93.015000 ;
      RECT 22.650000 169.565000 25.530000 169.715000 ;
      RECT 22.720000 104.025000 25.530000 104.175000 ;
      RECT 22.745000  92.715000 23.345000  92.865000 ;
      RECT 22.800000 169.715000 25.530000 169.865000 ;
      RECT 22.870000 103.875000 25.530000 104.025000 ;
      RECT 22.895000  92.565000 23.345000  92.715000 ;
      RECT 22.945000  92.375000 23.345000  93.790000 ;
      RECT 22.950000 169.865000 25.530000 170.015000 ;
      RECT 23.020000 103.725000 25.530000 103.875000 ;
      RECT 23.045000  92.415000 23.345000  92.565000 ;
      RECT 23.100000 170.015000 25.530000 170.165000 ;
      RECT 23.170000 103.575000 25.530000 103.725000 ;
      RECT 23.195000  92.265000 23.345000  92.415000 ;
      RECT 23.250000 170.165000 25.530000 170.315000 ;
      RECT 23.320000 103.425000 25.530000 103.575000 ;
      RECT 23.400000 170.315000 25.530000 170.465000 ;
      RECT 23.470000 103.275000 25.530000 103.425000 ;
      RECT 23.550000 170.465000 25.530000 170.615000 ;
      RECT 23.620000 103.125000 25.530000 103.275000 ;
      RECT 23.700000 170.615000 25.530000 170.765000 ;
      RECT 23.770000 102.975000 25.530000 103.125000 ;
      RECT 23.850000 170.765000 25.530000 170.915000 ;
      RECT 23.920000 102.825000 25.530000 102.975000 ;
      RECT 24.000000 170.915000 25.530000 171.065000 ;
      RECT 24.070000 102.675000 25.530000 102.825000 ;
      RECT 24.150000 171.065000 25.530000 171.215000 ;
      RECT 24.220000 102.525000 25.530000 102.675000 ;
      RECT 24.300000 171.215000 25.530000 171.365000 ;
      RECT 24.370000 102.375000 25.530000 102.525000 ;
      RECT 24.450000 171.365000 25.530000 171.515000 ;
      RECT 24.520000 102.225000 25.530000 102.375000 ;
      RECT 24.520000 102.225000 25.530000 104.845000 ;
      RECT 24.525000 102.220000 25.530000 102.225000 ;
      RECT 24.600000 171.515000 25.530000 171.665000 ;
      RECT 24.675000 102.070000 25.535000 102.220000 ;
      RECT 24.695000   0.000000 25.495000  90.225000 ;
      RECT 24.695000  90.225000 25.095000  90.625000 ;
      RECT 24.750000 171.665000 25.530000 171.815000 ;
      RECT 24.795000   0.000000 25.495000  90.225000 ;
      RECT 24.795000  90.225000 25.345000  90.375000 ;
      RECT 24.795000  90.375000 25.195000  90.525000 ;
      RECT 24.795000  90.525000 25.045000  90.675000 ;
      RECT 24.795000  90.675000 24.895000  90.825000 ;
      RECT 24.825000 101.920000 25.685000 102.070000 ;
      RECT 24.900000 171.815000 25.530000 171.965000 ;
      RECT 24.975000 101.770000 25.835000 101.920000 ;
      RECT 25.050000 171.965000 25.530000 172.115000 ;
      RECT 25.125000 101.620000 25.985000 101.770000 ;
      RECT 25.200000 172.115000 25.530000 172.265000 ;
      RECT 25.275000 101.470000 26.135000 101.620000 ;
      RECT 25.350000 172.265000 25.530000 172.415000 ;
      RECT 25.410000 172.475000 25.530000 195.500000 ;
      RECT 25.425000 101.320000 26.285000 101.470000 ;
      RECT 25.500000 172.415000 25.530000 172.565000 ;
      RECT 25.575000 101.170000 26.435000 101.320000 ;
      RECT 25.725000 101.020000 26.585000 101.170000 ;
      RECT 25.875000 100.870000 26.735000 101.020000 ;
      RECT 26.025000 100.720000 26.885000 100.870000 ;
      RECT 26.175000 100.570000 27.035000 100.720000 ;
      RECT 26.325000 100.420000 27.185000 100.570000 ;
      RECT 26.475000 100.270000 27.335000 100.420000 ;
      RECT 26.625000 100.120000 27.485000 100.270000 ;
      RECT 26.775000  99.970000 27.635000 100.120000 ;
      RECT 26.925000  99.820000 27.785000  99.970000 ;
      RECT 27.075000  99.670000 27.935000  99.820000 ;
      RECT 27.225000  99.520000 28.085000  99.670000 ;
      RECT 27.375000  99.370000 28.235000  99.520000 ;
      RECT 27.525000  99.220000 28.385000  99.370000 ;
      RECT 27.675000  99.070000 28.535000  99.220000 ;
      RECT 27.825000  98.920000 28.685000  99.070000 ;
      RECT 27.975000  98.770000 28.835000  98.920000 ;
      RECT 28.125000  98.620000 28.985000  98.770000 ;
      RECT 28.275000  98.470000 29.135000  98.620000 ;
      RECT 28.425000  98.320000 29.285000  98.470000 ;
      RECT 28.575000  98.170000 29.435000  98.320000 ;
      RECT 28.725000  98.020000 29.585000  98.170000 ;
      RECT 28.875000  97.870000 29.735000  98.020000 ;
      RECT 29.025000  97.720000 29.885000  97.870000 ;
      RECT 29.175000  97.570000 30.035000  97.720000 ;
      RECT 29.325000  97.420000 30.185000  97.570000 ;
      RECT 29.475000  97.270000 30.335000  97.420000 ;
      RECT 29.625000  97.120000 30.485000  97.270000 ;
      RECT 29.775000  96.970000 30.635000  97.120000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  96.210000 30.935000  96.820000 ;
      RECT 29.925000  96.210000 31.395000  96.360000 ;
      RECT 29.925000  96.360000 31.245000  96.510000 ;
      RECT 29.925000  96.510000 31.095000  96.660000 ;
      RECT 29.925000  96.660000 30.945000  96.810000 ;
      RECT 29.925000  96.810000 30.935000  96.820000 ;
      RECT 29.925000  96.820000 30.785000  96.970000 ;
      RECT 29.950000  93.240000 31.520000  93.265000 ;
      RECT 30.100000  93.090000 31.370000  93.240000 ;
      RECT 30.250000  92.940000 31.220000  93.090000 ;
      RECT 30.400000  92.790000 31.070000  92.940000 ;
      RECT 30.400000  92.790000 31.545000  93.265000 ;
      RECT 32.330000  99.865000 37.490000 110.785000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 42.455000 110.785000 ;
      RECT 32.330000 105.820000 42.455000 175.185000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 170.295000 37.565000 175.185000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.220000 175.185000 37.565000 190.420000 ;
      RECT 37.220000 175.270000 37.305000 175.355000 ;
      RECT 37.220000 175.355000 37.565000 190.420000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.295000   0.000000 37.490000 100.060000 ;
      RECT 37.295000 100.060000 37.490000 105.025000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.480000 175.270000 37.565000 175.355000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 101.970000 44.860000 102.580000 ;
      RECT 43.265000 100.355000 44.835000 100.380000 ;
      RECT 43.390000 101.970000 44.860000 102.120000 ;
      RECT 43.415000 100.205000 44.685000 100.355000 ;
      RECT 43.540000 102.120000 44.860000 102.270000 ;
      RECT 43.565000 100.055000 44.535000 100.205000 ;
      RECT 43.690000 102.270000 44.860000 102.420000 ;
      RECT 43.715000  99.905000 44.385000 100.055000 ;
      RECT 43.715000  99.905000 44.860000 100.380000 ;
      RECT 43.840000 102.420000 44.860000 102.570000 ;
      RECT 43.850000 102.570000 44.860000 102.580000 ;
      RECT 43.850000 102.580000 50.265000 107.985000 ;
      RECT 44.000000 102.580000 44.860000 102.730000 ;
      RECT 44.150000 102.730000 45.010000 102.880000 ;
      RECT 44.300000 102.880000 45.160000 103.030000 ;
      RECT 44.450000 103.030000 45.310000 103.180000 ;
      RECT 44.600000 103.180000 45.460000 103.330000 ;
      RECT 44.750000 103.330000 45.610000 103.480000 ;
      RECT 44.900000 103.480000 45.760000 103.630000 ;
      RECT 45.050000 103.630000 45.910000 103.780000 ;
      RECT 45.200000 103.780000 46.060000 103.930000 ;
      RECT 45.350000 103.930000 46.210000 104.080000 ;
      RECT 45.500000 104.080000 46.360000 104.230000 ;
      RECT 45.650000 104.230000 46.510000 104.380000 ;
      RECT 45.800000 104.380000 46.660000 104.530000 ;
      RECT 45.950000 104.530000 46.810000 104.680000 ;
      RECT 46.100000 104.680000 46.960000 104.830000 ;
      RECT 46.250000 104.830000 47.110000 104.980000 ;
      RECT 46.400000 104.980000 47.260000 105.130000 ;
      RECT 46.550000 105.130000 47.410000 105.280000 ;
      RECT 46.700000 105.280000 47.560000 105.430000 ;
      RECT 46.850000 105.430000 47.710000 105.580000 ;
      RECT 47.000000 105.580000 47.860000 105.730000 ;
      RECT 47.150000 105.730000 48.010000 105.880000 ;
      RECT 47.300000 105.880000 48.160000 106.030000 ;
      RECT 47.450000 106.030000 48.310000 106.180000 ;
      RECT 47.600000 106.180000 48.460000 106.330000 ;
      RECT 47.750000 106.330000 48.610000 106.480000 ;
      RECT 47.900000 106.480000 48.760000 106.630000 ;
      RECT 48.050000 106.630000 48.910000 106.780000 ;
      RECT 48.200000 106.780000 49.060000 106.930000 ;
      RECT 48.350000 106.930000 49.210000 107.080000 ;
      RECT 48.500000 107.080000 49.360000 107.230000 ;
      RECT 48.650000 107.230000 49.510000 107.380000 ;
      RECT 48.800000 107.380000 49.660000 107.530000 ;
      RECT 48.950000 107.530000 49.810000 107.680000 ;
      RECT 49.100000 107.680000 49.960000 107.830000 ;
      RECT 49.250000 107.830000 50.110000 107.980000 ;
      RECT 49.255000 107.980000 50.260000 107.985000 ;
      RECT 49.255000 107.985000 50.265000 108.135000 ;
      RECT 49.255000 107.985000 52.885000 110.605000 ;
      RECT 49.255000 108.135000 50.415000 108.285000 ;
      RECT 49.255000 108.285000 50.565000 108.435000 ;
      RECT 49.255000 108.435000 50.715000 108.585000 ;
      RECT 49.255000 108.585000 50.865000 108.735000 ;
      RECT 49.255000 108.735000 51.015000 108.885000 ;
      RECT 49.255000 108.885000 51.165000 109.035000 ;
      RECT 49.255000 109.035000 51.315000 109.185000 ;
      RECT 49.255000 109.185000 51.465000 109.335000 ;
      RECT 49.255000 109.335000 51.615000 109.485000 ;
      RECT 49.255000 109.485000 51.765000 109.635000 ;
      RECT 49.255000 109.635000 51.915000 109.785000 ;
      RECT 49.255000 109.785000 52.065000 109.935000 ;
      RECT 49.255000 109.935000 52.215000 110.085000 ;
      RECT 49.255000 110.085000 52.365000 110.235000 ;
      RECT 49.255000 110.235000 52.515000 110.385000 ;
      RECT 49.255000 110.385000 52.665000 110.535000 ;
      RECT 49.255000 110.535000 52.815000 110.605000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 168.970000 49.375000 172.480000 ;
      RECT 49.255000 168.970000 52.735000 169.120000 ;
      RECT 49.255000 169.120000 52.585000 169.270000 ;
      RECT 49.255000 169.270000 52.435000 169.420000 ;
      RECT 49.255000 169.420000 52.285000 169.570000 ;
      RECT 49.255000 169.570000 52.135000 169.720000 ;
      RECT 49.255000 169.720000 51.985000 169.870000 ;
      RECT 49.255000 169.870000 51.835000 170.020000 ;
      RECT 49.255000 170.020000 51.685000 170.170000 ;
      RECT 49.255000 170.170000 51.535000 170.320000 ;
      RECT 49.255000 170.320000 51.385000 170.470000 ;
      RECT 49.255000 170.470000 51.235000 170.620000 ;
      RECT 49.255000 170.620000 51.085000 170.770000 ;
      RECT 49.255000 170.770000 50.935000 170.920000 ;
      RECT 49.255000 170.920000 50.785000 171.070000 ;
      RECT 49.255000 171.070000 50.635000 171.220000 ;
      RECT 49.255000 171.220000 50.485000 171.370000 ;
      RECT 49.255000 171.370000 50.335000 171.520000 ;
      RECT 49.255000 171.520000 50.185000 171.670000 ;
      RECT 49.255000 171.670000 50.035000 171.820000 ;
      RECT 49.255000 171.820000 49.885000 171.970000 ;
      RECT 49.255000 171.970000 49.735000 172.120000 ;
      RECT 49.255000 172.120000 49.585000 172.270000 ;
      RECT 49.255000 172.270000 49.435000 172.420000 ;
      RECT 49.255000 172.420000 49.285000 172.570000 ;
      RECT 49.255000 172.480000 49.375000 190.420000 ;
      RECT 49.290000   0.000000 49.990000  89.650000 ;
      RECT 49.290000   0.000000 50.090000  90.310000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.310000 55.765000  95.985000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.985000 57.915000  98.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 59.330000  99.550000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.550000 61.200000 101.420000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.310000 101.420000 61.200000 107.795000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.685000 107.795000 61.200000 172.855000 ;
      RECT 59.685000 107.945000 59.835000 108.095000 ;
      RECT 59.685000 108.095000 59.985000 108.245000 ;
      RECT 59.685000 108.245000 60.135000 108.395000 ;
      RECT 59.685000 108.395000 60.285000 108.545000 ;
      RECT 59.685000 108.545000 60.435000 108.695000 ;
      RECT 59.685000 108.695000 60.585000 108.845000 ;
      RECT 59.685000 108.845000 60.735000 108.995000 ;
      RECT 59.685000 108.995000 60.885000 109.145000 ;
      RECT 59.685000 109.145000 61.035000 109.210000 ;
      RECT 59.685000 109.210000 61.100000 172.855000 ;
      RECT 59.685000 172.855000 61.200000 173.620000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.835000 172.855000 61.100000 173.005000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.985000 173.005000 61.100000 173.155000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.135000 173.155000 61.100000 173.305000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.285000 173.305000 61.100000 173.455000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.435000 173.455000 61.100000 173.605000 ;
      RECT 60.450000 173.620000 75.000000 174.515000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 173.605000 61.100000 173.720000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.345000 173.720000 75.000000 190.440000 ;
      RECT 61.345000 173.720000 75.000000 200.000000 ;
      RECT 61.345000 174.470000 75.000000 174.515000 ;
      RECT 61.345000 174.515000 75.000000 190.440000 ;
      RECT 74.590000   0.000000 75.000000 173.620000 ;
      RECT 74.690000   0.000000 75.000000 173.720000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   0.535000 ;
      RECT  0.000000  96.585000 75.000000 137.725000 ;
      RECT  0.000000 137.725000 35.045000 147.535000 ;
      RECT  0.000000 147.535000 75.000000 174.185000 ;
      RECT  2.565000  15.035000 72.435000  18.285000 ;
      RECT  2.870000   0.000000 72.130000  15.035000 ;
      RECT  2.870000  18.285000 72.130000  96.585000 ;
      RECT  2.870000 174.185000 72.130000 200.000000 ;
      RECT 39.570000 137.725000 75.000000 147.535000 ;
  END
END sky130_fd_io__top_ground_hvc_wpad
MACRO sky130_fd_io__top_power_hvc_wpad
  CLASS PAD ;
  ORIGIN  0.000000  0.000000 ;
  FOREIGN sky130_fd_io__top_power_hvc_wpad  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN P_PAD
    ANTENNAPARTIALMETALSIDEAREA  284.1730 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT  4.800000 104.230000 70.200000 166.570000 ;
        RECT  4.930000 104.100000 70.070000 104.230000 ;
        RECT  5.200000 166.570000 69.800000 166.970000 ;
        RECT  5.330000 103.700000 69.670000 104.100000 ;
        RECT  5.600000 166.970000 69.400000 167.370000 ;
        RECT  5.730000 103.300000 69.270000 103.700000 ;
        RECT  6.000000 167.370000 69.000000 167.770000 ;
        RECT  6.130000 102.900000 68.870000 103.300000 ;
        RECT  6.400000 167.770000 68.600000 168.170000 ;
        RECT  6.530000 102.500000 68.470000 102.900000 ;
        RECT  6.800000 168.170000 68.200000 168.570000 ;
        RECT  6.930000 102.100000 68.070000 102.500000 ;
        RECT  7.200000 168.570000 67.800000 168.970000 ;
        RECT  7.330000 101.700000 67.670000 102.100000 ;
        RECT  7.600000 168.970000 67.400000 169.370000 ;
        RECT  7.730000 101.300000 67.270000 101.700000 ;
        RECT  8.000000 169.370000 67.000000 169.770000 ;
        RECT  8.130000 100.900000 66.870000 101.300000 ;
        RECT  8.400000 169.770000 66.600000 170.170000 ;
        RECT  8.530000 100.500000 66.470000 100.900000 ;
        RECT  8.800000 170.170000 66.200000 170.570000 ;
        RECT  8.930000 100.100000 66.070000 100.500000 ;
        RECT  9.200000 170.570000 65.800000 170.970000 ;
        RECT  9.330000  99.700000 65.670000 100.100000 ;
        RECT  9.600000 170.970000 65.400000 171.370000 ;
        RECT  9.730000  99.300000 65.270000  99.700000 ;
        RECT 10.000000 171.370000 65.000000 171.770000 ;
        RECT 10.130000  98.900000 64.870000  99.300000 ;
        RECT 10.400000 171.770000 64.600000 172.170000 ;
        RECT 10.530000  98.500000 64.470000  98.900000 ;
        RECT 10.800000 172.170000 64.200000 172.570000 ;
        RECT 10.930000  98.100000 64.070000  98.500000 ;
        RECT 11.200000 172.570000 63.800000 172.970000 ;
        RECT 11.330000  97.700000 63.670000  98.100000 ;
        RECT 11.330000 172.970000 63.670000 173.100000 ;
    END
  END P_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.620000 185.295000 74.290000 190.015000 ;
        RECT 16.805000  47.455000 74.290000  54.765000 ;
        RECT 16.805000 139.455000 74.290000 146.710000 ;
        RECT 16.805000 162.455000 74.290000 171.155000 ;
        RECT 16.875000 146.710000 74.290000 146.780000 ;
        RECT 16.945000 146.780000 74.290000 146.850000 ;
        RECT 17.015000 146.850000 74.290000 146.920000 ;
        RECT 17.085000 146.920000 74.290000 146.990000 ;
        RECT 17.155000 146.990000 74.290000 147.060000 ;
        RECT 17.225000 147.060000 74.290000 147.130000 ;
        RECT 17.295000 147.130000 74.290000 147.200000 ;
        RECT 17.365000 147.200000 74.290000 147.270000 ;
        RECT 17.435000 147.270000 74.290000 147.340000 ;
        RECT 17.505000 147.340000 74.290000 147.410000 ;
        RECT 17.530000  54.765000 74.290000  54.835000 ;
        RECT 17.575000 147.410000 74.290000 147.480000 ;
        RECT 17.600000  54.835000 74.290000  54.905000 ;
        RECT 17.645000 147.480000 74.290000 147.550000 ;
        RECT 17.670000  54.905000 74.290000  54.975000 ;
        RECT 17.715000 147.550000 74.290000 147.620000 ;
        RECT 17.740000  54.975000 74.290000  55.045000 ;
        RECT 17.785000 147.620000 74.290000 147.690000 ;
        RECT 17.810000  55.045000 74.290000  55.115000 ;
        RECT 17.855000 147.690000 74.290000 147.760000 ;
        RECT 17.880000  55.115000 74.290000  55.185000 ;
        RECT 17.925000 147.760000 74.290000 147.830000 ;
        RECT 17.950000  55.185000 74.290000  55.255000 ;
        RECT 17.995000 147.830000 74.290000 147.900000 ;
        RECT 18.020000  55.255000 74.290000  55.325000 ;
        RECT 18.065000 147.900000 74.290000 147.970000 ;
        RECT 18.090000  55.325000 74.290000  55.395000 ;
        RECT 18.135000 147.970000 74.290000 148.040000 ;
        RECT 18.160000  55.395000 74.290000  55.465000 ;
        RECT 18.205000 148.040000 74.290000 148.110000 ;
        RECT 18.230000  55.465000 74.290000  55.535000 ;
        RECT 18.250000 148.110000 74.290000 148.155000 ;
        RECT 18.300000  55.535000 74.290000  55.605000 ;
        RECT 18.370000  55.605000 74.290000  55.675000 ;
        RECT 18.410000  74.155000 74.290000  74.415000 ;
        RECT 18.440000  55.675000 74.290000  55.745000 ;
        RECT 18.510000  55.745000 74.290000  55.815000 ;
        RECT 18.580000  55.815000 74.290000  55.885000 ;
        RECT 18.650000  55.885000 74.290000  55.955000 ;
        RECT 18.720000  55.955000 74.290000  56.025000 ;
        RECT 18.790000  56.025000 74.290000  56.095000 ;
        RECT 18.850000  56.095000 74.290000  56.155000 ;
        RECT 23.690000  74.415000 74.290000  74.485000 ;
        RECT 23.700000  74.105000 74.290000  74.155000 ;
        RECT 23.760000  74.485000 74.290000  74.555000 ;
        RECT 23.770000  74.035000 74.290000  74.105000 ;
        RECT 23.830000  74.555000 74.290000  74.625000 ;
        RECT 23.840000  73.965000 74.290000  74.035000 ;
        RECT 23.900000  74.625000 74.290000  74.695000 ;
        RECT 23.910000  73.895000 74.290000  73.965000 ;
        RECT 23.970000  74.695000 74.290000  74.765000 ;
        RECT 23.980000  73.825000 74.290000  73.895000 ;
        RECT 24.040000  74.765000 74.290000  74.835000 ;
        RECT 24.050000  73.755000 74.290000  73.825000 ;
        RECT 24.110000  74.835000 74.290000  74.905000 ;
        RECT 24.120000  73.685000 74.290000  73.755000 ;
        RECT 24.180000  74.905000 74.290000  74.975000 ;
        RECT 24.190000  73.615000 74.290000  73.685000 ;
        RECT 24.250000  74.975000 74.290000  75.045000 ;
        RECT 24.260000  73.545000 74.290000  73.615000 ;
        RECT 24.320000  75.045000 74.290000  75.115000 ;
        RECT 24.330000  73.475000 74.290000  73.545000 ;
        RECT 24.390000  75.115000 74.290000  75.185000 ;
        RECT 24.400000  73.405000 74.290000  73.475000 ;
        RECT 24.460000  75.185000 74.290000  75.255000 ;
        RECT 24.470000  73.335000 74.290000  73.405000 ;
        RECT 24.530000  75.255000 74.290000  75.325000 ;
        RECT 24.540000  73.265000 74.290000  73.335000 ;
        RECT 24.600000  75.325000 74.290000  75.395000 ;
        RECT 24.610000  73.195000 74.290000  73.265000 ;
        RECT 24.670000  75.395000 74.290000  75.465000 ;
        RECT 24.680000  73.125000 74.290000  73.195000 ;
        RECT 24.740000  75.465000 74.290000  75.535000 ;
        RECT 24.750000  73.055000 74.290000  73.125000 ;
        RECT 24.810000  75.535000 74.290000  75.605000 ;
        RECT 24.820000  70.455000 74.290000  72.985000 ;
        RECT 24.820000  72.985000 74.290000  73.055000 ;
        RECT 24.820000  75.605000 74.290000  75.615000 ;
        RECT 24.820000  75.615000 74.290000  79.155000 ;
        RECT 24.820000  93.455000 74.290000 102.155000 ;
        RECT 24.820000 116.455000 74.290000 125.155000 ;
        RECT 37.890000  12.295000 74.290000  25.660000 ;
        RECT 46.750000  12.265000 74.290000  12.295000 ;
        RECT 46.820000  12.195000 74.290000  12.265000 ;
        RECT 46.890000  12.125000 74.290000  12.195000 ;
        RECT 46.960000  12.055000 74.290000  12.125000 ;
        RECT 47.030000  11.985000 74.290000  12.055000 ;
        RECT 47.100000  11.915000 74.290000  11.985000 ;
        RECT 47.170000  11.845000 74.290000  11.915000 ;
        RECT 47.240000  11.775000 74.290000  11.845000 ;
        RECT 47.310000  11.705000 74.290000  11.775000 ;
        RECT 47.380000  11.635000 74.290000  11.705000 ;
        RECT 47.450000  11.565000 74.290000  11.635000 ;
        RECT 47.520000  11.495000 74.290000  11.565000 ;
        RECT 47.590000  11.425000 74.290000  11.495000 ;
        RECT 47.660000  11.355000 74.290000  11.425000 ;
        RECT 47.730000  11.285000 74.290000  11.355000 ;
        RECT 47.800000  11.215000 74.290000  11.285000 ;
        RECT 47.870000  11.145000 74.290000  11.215000 ;
        RECT 47.940000  11.075000 74.290000  11.145000 ;
        RECT 48.010000  11.005000 74.290000  11.075000 ;
        RECT 48.080000  10.935000 74.290000  11.005000 ;
        RECT 48.150000  10.865000 74.290000  10.935000 ;
        RECT 48.220000  10.795000 74.290000  10.865000 ;
        RECT 48.290000  10.725000 74.290000  10.795000 ;
        RECT 48.360000  10.655000 74.290000  10.725000 ;
        RECT 48.430000  10.585000 74.290000  10.655000 ;
        RECT 48.500000  10.515000 74.290000  10.585000 ;
        RECT 48.570000  10.445000 74.290000  10.515000 ;
        RECT 48.640000  10.375000 74.290000  10.445000 ;
        RECT 48.710000  10.305000 74.290000  10.375000 ;
        RECT 48.780000  10.235000 74.290000  10.305000 ;
        RECT 48.850000  10.165000 74.290000  10.235000 ;
        RECT 48.920000  10.095000 74.290000  10.165000 ;
        RECT 48.990000  10.025000 74.290000  10.095000 ;
        RECT 49.060000   9.955000 74.290000  10.025000 ;
        RECT 49.130000   9.885000 74.290000   9.955000 ;
        RECT 49.200000   9.815000 74.290000   9.885000 ;
        RECT 49.270000   9.745000 74.290000   9.815000 ;
        RECT 49.340000   9.675000 74.290000   9.745000 ;
        RECT 49.410000   9.605000 74.290000   9.675000 ;
        RECT 49.480000   9.535000 74.290000   9.605000 ;
        RECT 49.550000   9.465000 74.290000   9.535000 ;
        RECT 49.620000   9.395000 74.290000   9.465000 ;
        RECT 49.690000   9.325000 74.290000   9.395000 ;
        RECT 49.760000   9.255000 74.290000   9.325000 ;
        RECT 49.830000   9.185000 74.290000   9.255000 ;
        RECT 49.900000   9.115000 74.290000   9.185000 ;
        RECT 49.970000   9.045000 74.290000   9.115000 ;
        RECT 50.040000   8.975000 74.290000   9.045000 ;
        RECT 50.110000   8.905000 74.290000   8.975000 ;
        RECT 50.180000   8.835000 74.290000   8.905000 ;
        RECT 50.250000   8.765000 74.290000   8.835000 ;
        RECT 50.320000   8.695000 74.290000   8.765000 ;
        RECT 50.390000   0.000000 74.290000   8.625000 ;
        RECT 50.390000   8.625000 74.290000   8.695000 ;
        RECT 55.885000  25.660000 74.290000  25.730000 ;
        RECT 55.955000  25.730000 74.290000  25.800000 ;
        RECT 56.025000  25.800000 74.290000  25.870000 ;
        RECT 56.095000  25.870000 74.290000  25.940000 ;
        RECT 56.165000  25.940000 74.290000  26.010000 ;
        RECT 56.235000  26.010000 74.290000  26.080000 ;
        RECT 56.305000  26.080000 74.290000  26.150000 ;
        RECT 56.375000  26.150000 74.290000  26.220000 ;
        RECT 56.445000  26.220000 74.290000  26.290000 ;
        RECT 56.515000  26.290000 74.290000  26.360000 ;
        RECT 56.585000  26.360000 74.290000  26.430000 ;
        RECT 56.655000  26.430000 74.290000  26.500000 ;
        RECT 56.725000  26.500000 74.290000  26.570000 ;
        RECT 56.795000  26.570000 74.290000  26.640000 ;
        RECT 56.865000  26.640000 74.290000  26.710000 ;
        RECT 56.935000  26.710000 74.290000  26.780000 ;
        RECT 57.005000  26.780000 74.290000  26.850000 ;
        RECT 57.075000  26.850000 74.290000  26.920000 ;
        RECT 57.145000  26.920000 74.290000  26.990000 ;
        RECT 57.215000  26.990000 74.290000  27.060000 ;
        RECT 57.285000  27.060000 74.290000  27.130000 ;
        RECT 57.355000  27.130000 74.290000  27.200000 ;
        RECT 57.425000  27.200000 74.290000  27.270000 ;
        RECT 57.495000  27.270000 74.290000  27.340000 ;
        RECT 57.540000  47.390000 74.290000  47.455000 ;
        RECT 57.540000  70.420000 74.290000  70.455000 ;
        RECT 57.540000 116.390000 74.290000 116.455000 ;
        RECT 57.540000 139.425000 74.290000 139.455000 ;
        RECT 57.540000 162.440000 74.290000 162.455000 ;
        RECT 57.555000 148.155000 74.290000 148.225000 ;
        RECT 57.565000  27.340000 74.290000  27.410000 ;
        RECT 57.595000  56.155000 74.290000  56.225000 ;
        RECT 57.610000  47.320000 74.290000  47.390000 ;
        RECT 57.610000  70.350000 74.290000  70.420000 ;
        RECT 57.610000  93.410000 74.290000  93.455000 ;
        RECT 57.610000 116.320000 74.290000 116.390000 ;
        RECT 57.610000 139.355000 74.290000 139.425000 ;
        RECT 57.610000 162.370000 74.290000 162.440000 ;
        RECT 57.625000  79.155000 74.290000  79.225000 ;
        RECT 57.625000 102.155000 74.290000 102.225000 ;
        RECT 57.625000 125.155000 74.290000 125.225000 ;
        RECT 57.625000 148.225000 74.290000 148.295000 ;
        RECT 57.635000  27.410000 74.290000  27.480000 ;
        RECT 57.635000 171.155000 74.290000 171.225000 ;
        RECT 57.665000  56.225000 74.290000  56.295000 ;
        RECT 57.680000  47.250000 74.290000  47.320000 ;
        RECT 57.680000  70.280000 74.290000  70.350000 ;
        RECT 57.680000  93.340000 74.290000  93.410000 ;
        RECT 57.680000 116.250000 74.290000 116.320000 ;
        RECT 57.680000 139.285000 74.290000 139.355000 ;
        RECT 57.680000 162.300000 74.290000 162.370000 ;
        RECT 57.695000  79.225000 74.290000  79.295000 ;
        RECT 57.695000 102.225000 74.290000 102.295000 ;
        RECT 57.695000 125.225000 74.290000 125.295000 ;
        RECT 57.695000 148.295000 74.290000 148.365000 ;
        RECT 57.705000  27.480000 74.290000  27.550000 ;
        RECT 57.705000 171.225000 74.290000 171.295000 ;
        RECT 57.735000  56.295000 74.290000  56.365000 ;
        RECT 57.750000  47.180000 74.290000  47.250000 ;
        RECT 57.750000  70.210000 74.290000  70.280000 ;
        RECT 57.750000  93.270000 74.290000  93.340000 ;
        RECT 57.750000 116.180000 74.290000 116.250000 ;
        RECT 57.750000 139.215000 74.290000 139.285000 ;
        RECT 57.750000 162.230000 74.290000 162.300000 ;
        RECT 57.765000  79.295000 74.290000  79.365000 ;
        RECT 57.765000 102.295000 74.290000 102.365000 ;
        RECT 57.765000 125.295000 74.290000 125.365000 ;
        RECT 57.765000 148.365000 74.290000 148.435000 ;
        RECT 57.775000  27.550000 74.290000  27.620000 ;
        RECT 57.775000 171.295000 74.290000 171.365000 ;
        RECT 57.805000  56.365000 74.290000  56.435000 ;
        RECT 57.820000  47.110000 74.290000  47.180000 ;
        RECT 57.820000  70.140000 74.290000  70.210000 ;
        RECT 57.820000  93.200000 74.290000  93.270000 ;
        RECT 57.820000 116.110000 74.290000 116.180000 ;
        RECT 57.820000 139.145000 74.290000 139.215000 ;
        RECT 57.820000 162.160000 74.290000 162.230000 ;
        RECT 57.835000  79.365000 74.290000  79.435000 ;
        RECT 57.835000 102.365000 74.290000 102.435000 ;
        RECT 57.835000 125.365000 74.290000 125.435000 ;
        RECT 57.835000 148.435000 74.290000 148.505000 ;
        RECT 57.845000  27.620000 74.290000  27.690000 ;
        RECT 57.845000 171.365000 74.290000 171.435000 ;
        RECT 57.875000  56.435000 74.290000  56.505000 ;
        RECT 57.890000  47.040000 74.290000  47.110000 ;
        RECT 57.890000  70.070000 74.290000  70.140000 ;
        RECT 57.890000  93.130000 74.290000  93.200000 ;
        RECT 57.890000 116.040000 74.290000 116.110000 ;
        RECT 57.890000 139.075000 74.290000 139.145000 ;
        RECT 57.890000 162.090000 74.290000 162.160000 ;
        RECT 57.905000  79.435000 74.290000  79.505000 ;
        RECT 57.905000 102.435000 74.290000 102.505000 ;
        RECT 57.905000 125.435000 74.290000 125.505000 ;
        RECT 57.905000 148.505000 74.290000 148.575000 ;
        RECT 57.915000  27.690000 74.290000  27.760000 ;
        RECT 57.915000 171.435000 74.290000 171.505000 ;
        RECT 57.945000  56.505000 74.290000  56.575000 ;
        RECT 57.960000  46.970000 74.290000  47.040000 ;
        RECT 57.960000  70.000000 74.290000  70.070000 ;
        RECT 57.960000  93.060000 74.290000  93.130000 ;
        RECT 57.960000 115.970000 74.290000 116.040000 ;
        RECT 57.960000 139.005000 74.290000 139.075000 ;
        RECT 57.960000 162.020000 74.290000 162.090000 ;
        RECT 57.975000  79.505000 74.290000  79.575000 ;
        RECT 57.975000 102.505000 74.290000 102.575000 ;
        RECT 57.975000 125.505000 74.290000 125.575000 ;
        RECT 57.975000 148.575000 74.290000 148.645000 ;
        RECT 57.985000  27.760000 74.290000  27.830000 ;
        RECT 57.985000 171.505000 74.290000 171.575000 ;
        RECT 58.015000  56.575000 74.290000  56.645000 ;
        RECT 58.030000  46.900000 74.290000  46.970000 ;
        RECT 58.030000  69.930000 74.290000  70.000000 ;
        RECT 58.030000  92.990000 74.290000  93.060000 ;
        RECT 58.030000 115.900000 74.290000 115.970000 ;
        RECT 58.030000 138.935000 74.290000 139.005000 ;
        RECT 58.030000 161.950000 74.290000 162.020000 ;
        RECT 58.045000  79.575000 74.290000  79.645000 ;
        RECT 58.045000 102.575000 74.290000 102.645000 ;
        RECT 58.045000 125.575000 74.290000 125.645000 ;
        RECT 58.045000 148.645000 74.290000 148.715000 ;
        RECT 58.055000  27.830000 74.290000  27.900000 ;
        RECT 58.055000 171.575000 74.290000 171.645000 ;
        RECT 58.085000  56.645000 74.290000  56.715000 ;
        RECT 58.100000  46.830000 74.290000  46.900000 ;
        RECT 58.100000  69.860000 74.290000  69.930000 ;
        RECT 58.100000  92.920000 74.290000  92.990000 ;
        RECT 58.100000 115.830000 74.290000 115.900000 ;
        RECT 58.100000 138.865000 74.290000 138.935000 ;
        RECT 58.100000 161.880000 74.290000 161.950000 ;
        RECT 58.115000  79.645000 74.290000  79.715000 ;
        RECT 58.115000 102.645000 74.290000 102.715000 ;
        RECT 58.115000 125.645000 74.290000 125.715000 ;
        RECT 58.115000 148.715000 74.290000 148.785000 ;
        RECT 58.125000  27.900000 74.290000  27.970000 ;
        RECT 58.125000 171.645000 74.290000 171.715000 ;
        RECT 58.155000  56.715000 74.290000  56.785000 ;
        RECT 58.170000  46.760000 74.290000  46.830000 ;
        RECT 58.170000  69.790000 74.290000  69.860000 ;
        RECT 58.170000  92.850000 74.290000  92.920000 ;
        RECT 58.170000 115.760000 74.290000 115.830000 ;
        RECT 58.170000 138.795000 74.290000 138.865000 ;
        RECT 58.170000 161.810000 74.290000 161.880000 ;
        RECT 58.185000  79.715000 74.290000  79.785000 ;
        RECT 58.185000 102.715000 74.290000 102.785000 ;
        RECT 58.185000 125.715000 74.290000 125.785000 ;
        RECT 58.185000 148.785000 74.290000 148.855000 ;
        RECT 58.195000  27.970000 74.290000  28.040000 ;
        RECT 58.195000 171.715000 74.290000 171.785000 ;
        RECT 58.225000  56.785000 74.290000  56.855000 ;
        RECT 58.240000  46.690000 74.290000  46.760000 ;
        RECT 58.240000  69.720000 74.290000  69.790000 ;
        RECT 58.240000  92.780000 74.290000  92.850000 ;
        RECT 58.240000 115.690000 74.290000 115.760000 ;
        RECT 58.240000 138.725000 74.290000 138.795000 ;
        RECT 58.240000 161.740000 74.290000 161.810000 ;
        RECT 58.255000  79.785000 74.290000  79.855000 ;
        RECT 58.255000 102.785000 74.290000 102.855000 ;
        RECT 58.255000 125.785000 74.290000 125.855000 ;
        RECT 58.255000 148.855000 74.290000 148.925000 ;
        RECT 58.265000  28.040000 74.290000  28.110000 ;
        RECT 58.265000 171.785000 74.290000 171.855000 ;
        RECT 58.295000  56.855000 74.290000  56.925000 ;
        RECT 58.310000  46.620000 74.290000  46.690000 ;
        RECT 58.310000  69.650000 74.290000  69.720000 ;
        RECT 58.310000  92.710000 74.290000  92.780000 ;
        RECT 58.310000 115.620000 74.290000 115.690000 ;
        RECT 58.310000 138.655000 74.290000 138.725000 ;
        RECT 58.310000 161.670000 74.290000 161.740000 ;
        RECT 58.325000  79.855000 74.290000  79.925000 ;
        RECT 58.325000 102.855000 74.290000 102.925000 ;
        RECT 58.325000 125.855000 74.290000 125.925000 ;
        RECT 58.325000 148.925000 74.290000 148.995000 ;
        RECT 58.335000  28.110000 74.290000  28.180000 ;
        RECT 58.335000 171.855000 74.290000 171.925000 ;
        RECT 58.365000  56.925000 74.290000  56.995000 ;
        RECT 58.380000  46.550000 74.290000  46.620000 ;
        RECT 58.380000  69.580000 74.290000  69.650000 ;
        RECT 58.380000  92.640000 74.290000  92.710000 ;
        RECT 58.380000 115.550000 74.290000 115.620000 ;
        RECT 58.380000 138.585000 74.290000 138.655000 ;
        RECT 58.380000 161.600000 74.290000 161.670000 ;
        RECT 58.395000  79.925000 74.290000  79.995000 ;
        RECT 58.395000 102.925000 74.290000 102.995000 ;
        RECT 58.395000 125.925000 74.290000 125.995000 ;
        RECT 58.395000 148.995000 74.290000 149.065000 ;
        RECT 58.405000  28.180000 74.290000  28.250000 ;
        RECT 58.405000 171.925000 74.290000 171.995000 ;
        RECT 58.435000  56.995000 74.290000  57.065000 ;
        RECT 58.450000  46.480000 74.290000  46.550000 ;
        RECT 58.450000  69.510000 74.290000  69.580000 ;
        RECT 58.450000  92.570000 74.290000  92.640000 ;
        RECT 58.450000 115.480000 74.290000 115.550000 ;
        RECT 58.450000 138.515000 74.290000 138.585000 ;
        RECT 58.450000 161.530000 74.290000 161.600000 ;
        RECT 58.465000  79.995000 74.290000  80.065000 ;
        RECT 58.465000 102.995000 74.290000 103.065000 ;
        RECT 58.465000 125.995000 74.290000 126.065000 ;
        RECT 58.465000 149.065000 74.290000 149.135000 ;
        RECT 58.475000  28.250000 74.290000  28.320000 ;
        RECT 58.475000 171.995000 74.290000 172.065000 ;
        RECT 58.505000  57.065000 74.290000  57.135000 ;
        RECT 58.520000  46.410000 74.290000  46.480000 ;
        RECT 58.520000  69.440000 74.290000  69.510000 ;
        RECT 58.520000  92.500000 74.290000  92.570000 ;
        RECT 58.520000 115.410000 74.290000 115.480000 ;
        RECT 58.520000 138.445000 74.290000 138.515000 ;
        RECT 58.520000 161.460000 74.290000 161.530000 ;
        RECT 58.535000  80.065000 74.290000  80.135000 ;
        RECT 58.535000 103.065000 74.290000 103.135000 ;
        RECT 58.535000 126.065000 74.290000 126.135000 ;
        RECT 58.535000 149.135000 74.290000 149.205000 ;
        RECT 58.545000  28.320000 74.290000  28.390000 ;
        RECT 58.545000 172.065000 74.290000 172.135000 ;
        RECT 58.575000  57.135000 74.290000  57.205000 ;
        RECT 58.590000  46.340000 74.290000  46.410000 ;
        RECT 58.590000  69.370000 74.290000  69.440000 ;
        RECT 58.590000  92.430000 74.290000  92.500000 ;
        RECT 58.590000 115.340000 74.290000 115.410000 ;
        RECT 58.590000 138.375000 74.290000 138.445000 ;
        RECT 58.590000 161.390000 74.290000 161.460000 ;
        RECT 58.605000  80.135000 74.290000  80.205000 ;
        RECT 58.605000 103.135000 74.290000 103.205000 ;
        RECT 58.605000 126.135000 74.290000 126.205000 ;
        RECT 58.605000 149.205000 74.290000 149.275000 ;
        RECT 58.615000  28.390000 74.290000  28.460000 ;
        RECT 58.615000 172.135000 74.290000 172.205000 ;
        RECT 58.645000  57.205000 74.290000  57.275000 ;
        RECT 58.660000  46.270000 74.290000  46.340000 ;
        RECT 58.660000  69.300000 74.290000  69.370000 ;
        RECT 58.660000  92.360000 74.290000  92.430000 ;
        RECT 58.660000 115.270000 74.290000 115.340000 ;
        RECT 58.660000 138.305000 74.290000 138.375000 ;
        RECT 58.660000 161.320000 74.290000 161.390000 ;
        RECT 58.675000  80.205000 74.290000  80.275000 ;
        RECT 58.675000 103.205000 74.290000 103.275000 ;
        RECT 58.675000 126.205000 74.290000 126.275000 ;
        RECT 58.675000 149.275000 74.290000 149.345000 ;
        RECT 58.685000  28.460000 74.290000  28.530000 ;
        RECT 58.685000 172.205000 74.290000 172.275000 ;
        RECT 58.715000  57.275000 74.290000  57.345000 ;
        RECT 58.730000  46.200000 74.290000  46.270000 ;
        RECT 58.730000  69.230000 74.290000  69.300000 ;
        RECT 58.730000  92.290000 74.290000  92.360000 ;
        RECT 58.730000 115.200000 74.290000 115.270000 ;
        RECT 58.730000 138.235000 74.290000 138.305000 ;
        RECT 58.730000 161.250000 74.290000 161.320000 ;
        RECT 58.730000 185.260000 74.290000 185.295000 ;
        RECT 58.745000  80.275000 74.290000  80.345000 ;
        RECT 58.745000 103.275000 74.290000 103.345000 ;
        RECT 58.745000 126.275000 74.290000 126.345000 ;
        RECT 58.745000 149.345000 74.290000 149.415000 ;
        RECT 58.755000  28.530000 74.290000  28.600000 ;
        RECT 58.755000 172.275000 74.290000 172.345000 ;
        RECT 58.785000  57.345000 74.290000  57.415000 ;
        RECT 58.800000  46.130000 74.290000  46.200000 ;
        RECT 58.800000  69.160000 74.290000  69.230000 ;
        RECT 58.800000  92.220000 74.290000  92.290000 ;
        RECT 58.800000 115.130000 74.290000 115.200000 ;
        RECT 58.800000 138.165000 74.290000 138.235000 ;
        RECT 58.800000 161.180000 74.290000 161.250000 ;
        RECT 58.800000 185.190000 74.290000 185.260000 ;
        RECT 58.815000  80.345000 74.290000  80.415000 ;
        RECT 58.815000 103.345000 74.290000 103.415000 ;
        RECT 58.815000 126.345000 74.290000 126.415000 ;
        RECT 58.815000 149.415000 74.290000 149.485000 ;
        RECT 58.825000  28.600000 74.290000  28.670000 ;
        RECT 58.825000 172.345000 74.290000 172.415000 ;
        RECT 58.855000  57.415000 74.290000  57.485000 ;
        RECT 58.870000  46.060000 74.290000  46.130000 ;
        RECT 58.870000  69.090000 74.290000  69.160000 ;
        RECT 58.870000  92.150000 74.290000  92.220000 ;
        RECT 58.870000 115.060000 74.290000 115.130000 ;
        RECT 58.870000 138.095000 74.290000 138.165000 ;
        RECT 58.870000 161.110000 74.290000 161.180000 ;
        RECT 58.870000 185.120000 74.290000 185.190000 ;
        RECT 58.885000  80.415000 74.290000  80.485000 ;
        RECT 58.885000 103.415000 74.290000 103.485000 ;
        RECT 58.885000 126.415000 74.290000 126.485000 ;
        RECT 58.885000 149.485000 74.290000 149.555000 ;
        RECT 58.895000  28.670000 74.290000  28.740000 ;
        RECT 58.895000 172.415000 74.290000 172.485000 ;
        RECT 58.925000  57.485000 74.290000  57.555000 ;
        RECT 58.940000  45.990000 74.290000  46.060000 ;
        RECT 58.940000  69.020000 74.290000  69.090000 ;
        RECT 58.940000  92.080000 74.290000  92.150000 ;
        RECT 58.940000 114.990000 74.290000 115.060000 ;
        RECT 58.940000 138.025000 74.290000 138.095000 ;
        RECT 58.940000 161.040000 74.290000 161.110000 ;
        RECT 58.940000 185.050000 74.290000 185.120000 ;
        RECT 58.955000  80.485000 74.290000  80.555000 ;
        RECT 58.955000 103.485000 74.290000 103.555000 ;
        RECT 58.955000 126.485000 74.290000 126.555000 ;
        RECT 58.955000 149.555000 74.290000 149.625000 ;
        RECT 58.965000  28.740000 74.290000  28.810000 ;
        RECT 58.965000 172.485000 74.290000 172.555000 ;
        RECT 58.995000  57.555000 74.290000  57.625000 ;
        RECT 59.010000  45.920000 74.290000  45.990000 ;
        RECT 59.010000  68.950000 74.290000  69.020000 ;
        RECT 59.010000  92.010000 74.290000  92.080000 ;
        RECT 59.010000 114.920000 74.290000 114.990000 ;
        RECT 59.010000 137.955000 74.290000 138.025000 ;
        RECT 59.010000 160.970000 74.290000 161.040000 ;
        RECT 59.010000 184.980000 74.290000 185.050000 ;
        RECT 59.025000  80.555000 74.290000  80.625000 ;
        RECT 59.025000 103.555000 74.290000 103.625000 ;
        RECT 59.025000 126.555000 74.290000 126.625000 ;
        RECT 59.025000 149.625000 74.290000 149.695000 ;
        RECT 59.035000  28.810000 74.290000  28.880000 ;
        RECT 59.035000 172.555000 74.290000 172.625000 ;
        RECT 59.065000  57.625000 74.290000  57.695000 ;
        RECT 59.080000  45.850000 74.290000  45.920000 ;
        RECT 59.080000  68.880000 74.290000  68.950000 ;
        RECT 59.080000  91.940000 74.290000  92.010000 ;
        RECT 59.080000 114.850000 74.290000 114.920000 ;
        RECT 59.080000 137.885000 74.290000 137.955000 ;
        RECT 59.080000 160.900000 74.290000 160.970000 ;
        RECT 59.080000 184.910000 74.290000 184.980000 ;
        RECT 59.095000  80.625000 74.290000  80.695000 ;
        RECT 59.095000 103.625000 74.290000 103.695000 ;
        RECT 59.095000 126.625000 74.290000 126.695000 ;
        RECT 59.095000 149.695000 74.290000 149.765000 ;
        RECT 59.105000  28.880000 74.290000  28.950000 ;
        RECT 59.105000 172.625000 74.290000 172.695000 ;
        RECT 59.135000  57.695000 74.290000  57.765000 ;
        RECT 59.150000  45.780000 74.290000  45.850000 ;
        RECT 59.150000  68.810000 74.290000  68.880000 ;
        RECT 59.150000  91.870000 74.290000  91.940000 ;
        RECT 59.150000 114.780000 74.290000 114.850000 ;
        RECT 59.150000 137.815000 74.290000 137.885000 ;
        RECT 59.150000 160.830000 74.290000 160.900000 ;
        RECT 59.150000 184.840000 74.290000 184.910000 ;
        RECT 59.165000  80.695000 74.290000  80.765000 ;
        RECT 59.165000 103.695000 74.290000 103.765000 ;
        RECT 59.165000 126.695000 74.290000 126.765000 ;
        RECT 59.165000 149.765000 74.290000 149.835000 ;
        RECT 59.175000  28.950000 74.290000  29.020000 ;
        RECT 59.175000 172.695000 74.290000 172.765000 ;
        RECT 59.205000  57.765000 74.290000  57.835000 ;
        RECT 59.220000  45.710000 74.290000  45.780000 ;
        RECT 59.220000  68.740000 74.290000  68.810000 ;
        RECT 59.220000  91.800000 74.290000  91.870000 ;
        RECT 59.220000 114.710000 74.290000 114.780000 ;
        RECT 59.220000 137.745000 74.290000 137.815000 ;
        RECT 59.220000 160.760000 74.290000 160.830000 ;
        RECT 59.220000 184.770000 74.290000 184.840000 ;
        RECT 59.235000  80.765000 74.290000  80.835000 ;
        RECT 59.235000 103.765000 74.290000 103.835000 ;
        RECT 59.235000 126.765000 74.290000 126.835000 ;
        RECT 59.235000 149.835000 74.290000 149.905000 ;
        RECT 59.245000  29.020000 74.290000  29.090000 ;
        RECT 59.245000 172.765000 74.290000 172.835000 ;
        RECT 59.275000  57.835000 74.290000  57.905000 ;
        RECT 59.290000  45.640000 74.290000  45.710000 ;
        RECT 59.290000  68.670000 74.290000  68.740000 ;
        RECT 59.290000  91.730000 74.290000  91.800000 ;
        RECT 59.290000 114.640000 74.290000 114.710000 ;
        RECT 59.290000 137.675000 74.290000 137.745000 ;
        RECT 59.290000 160.690000 74.290000 160.760000 ;
        RECT 59.290000 184.700000 74.290000 184.770000 ;
        RECT 59.305000  80.835000 74.290000  80.905000 ;
        RECT 59.305000 103.835000 74.290000 103.905000 ;
        RECT 59.305000 126.835000 74.290000 126.905000 ;
        RECT 59.305000 149.905000 74.290000 149.975000 ;
        RECT 59.315000  29.090000 74.290000  29.160000 ;
        RECT 59.315000 172.835000 74.290000 172.905000 ;
        RECT 59.345000  57.905000 74.290000  57.975000 ;
        RECT 59.360000  45.570000 74.290000  45.640000 ;
        RECT 59.360000  68.600000 74.290000  68.670000 ;
        RECT 59.360000  91.660000 74.290000  91.730000 ;
        RECT 59.360000 114.570000 74.290000 114.640000 ;
        RECT 59.360000 137.605000 74.290000 137.675000 ;
        RECT 59.360000 160.620000 74.290000 160.690000 ;
        RECT 59.360000 184.630000 74.290000 184.700000 ;
        RECT 59.375000  80.905000 74.290000  80.975000 ;
        RECT 59.375000 103.905000 74.290000 103.975000 ;
        RECT 59.375000 126.905000 74.290000 126.975000 ;
        RECT 59.375000 149.975000 74.290000 150.045000 ;
        RECT 59.385000  29.160000 74.290000  29.230000 ;
        RECT 59.385000 172.905000 74.290000 172.975000 ;
        RECT 59.415000  57.975000 74.290000  58.045000 ;
        RECT 59.430000  45.500000 74.290000  45.570000 ;
        RECT 59.430000  68.530000 74.290000  68.600000 ;
        RECT 59.430000  91.590000 74.290000  91.660000 ;
        RECT 59.430000 114.500000 74.290000 114.570000 ;
        RECT 59.430000 137.535000 74.290000 137.605000 ;
        RECT 59.430000 160.550000 74.290000 160.620000 ;
        RECT 59.430000 184.560000 74.290000 184.630000 ;
        RECT 59.445000  80.975000 74.290000  81.045000 ;
        RECT 59.445000 103.975000 74.290000 104.045000 ;
        RECT 59.445000 126.975000 74.290000 127.045000 ;
        RECT 59.445000 150.045000 74.290000 150.115000 ;
        RECT 59.455000  29.230000 74.290000  29.300000 ;
        RECT 59.455000 172.975000 74.290000 173.045000 ;
        RECT 59.485000  58.045000 74.290000  58.115000 ;
        RECT 59.500000  45.430000 74.290000  45.500000 ;
        RECT 59.500000  68.460000 74.290000  68.530000 ;
        RECT 59.500000  91.520000 74.290000  91.590000 ;
        RECT 59.500000 114.430000 74.290000 114.500000 ;
        RECT 59.500000 137.465000 74.290000 137.535000 ;
        RECT 59.500000 160.480000 74.290000 160.550000 ;
        RECT 59.500000 184.490000 74.290000 184.560000 ;
        RECT 59.515000  81.045000 74.290000  81.115000 ;
        RECT 59.515000 104.045000 74.290000 104.115000 ;
        RECT 59.515000 127.045000 74.290000 127.115000 ;
        RECT 59.515000 150.115000 74.290000 150.185000 ;
        RECT 59.525000  29.300000 74.290000  29.370000 ;
        RECT 59.525000 173.045000 74.290000 173.115000 ;
        RECT 59.555000  58.115000 74.290000  58.185000 ;
        RECT 59.570000  45.360000 74.290000  45.430000 ;
        RECT 59.570000  68.390000 74.290000  68.460000 ;
        RECT 59.570000  91.450000 74.290000  91.520000 ;
        RECT 59.570000 114.360000 74.290000 114.430000 ;
        RECT 59.570000 137.395000 74.290000 137.465000 ;
        RECT 59.570000 160.410000 74.290000 160.480000 ;
        RECT 59.570000 184.420000 74.290000 184.490000 ;
        RECT 59.585000  81.115000 74.290000  81.185000 ;
        RECT 59.585000 104.115000 74.290000 104.185000 ;
        RECT 59.585000 127.115000 74.290000 127.185000 ;
        RECT 59.585000 150.185000 74.290000 150.255000 ;
        RECT 59.595000  29.370000 74.290000  29.440000 ;
        RECT 59.595000 173.115000 74.290000 173.185000 ;
        RECT 59.625000  58.185000 74.290000  58.255000 ;
        RECT 59.640000  45.290000 74.290000  45.360000 ;
        RECT 59.640000  68.320000 74.290000  68.390000 ;
        RECT 59.640000  91.380000 74.290000  91.450000 ;
        RECT 59.640000 114.290000 74.290000 114.360000 ;
        RECT 59.640000 137.325000 74.290000 137.395000 ;
        RECT 59.640000 160.340000 74.290000 160.410000 ;
        RECT 59.640000 184.350000 74.290000 184.420000 ;
        RECT 59.655000  81.185000 74.290000  81.255000 ;
        RECT 59.655000 104.185000 74.290000 104.255000 ;
        RECT 59.655000 127.185000 74.290000 127.255000 ;
        RECT 59.655000 150.255000 74.290000 150.325000 ;
        RECT 59.665000  29.440000 74.290000  29.510000 ;
        RECT 59.665000 173.185000 74.290000 173.255000 ;
        RECT 59.695000  58.255000 74.290000  58.325000 ;
        RECT 59.710000  45.220000 74.290000  45.290000 ;
        RECT 59.710000  68.250000 74.290000  68.320000 ;
        RECT 59.710000  91.310000 74.290000  91.380000 ;
        RECT 59.710000 114.220000 74.290000 114.290000 ;
        RECT 59.710000 137.255000 74.290000 137.325000 ;
        RECT 59.710000 160.270000 74.290000 160.340000 ;
        RECT 59.710000 184.280000 74.290000 184.350000 ;
        RECT 59.725000  81.255000 74.290000  81.325000 ;
        RECT 59.725000 104.255000 74.290000 104.325000 ;
        RECT 59.725000 127.255000 74.290000 127.325000 ;
        RECT 59.725000 150.325000 74.290000 150.395000 ;
        RECT 59.735000  29.510000 74.290000  29.580000 ;
        RECT 59.735000 173.255000 74.290000 173.325000 ;
        RECT 59.765000  58.325000 74.290000  58.395000 ;
        RECT 59.780000  45.150000 74.290000  45.220000 ;
        RECT 59.780000  68.180000 74.290000  68.250000 ;
        RECT 59.780000  91.240000 74.290000  91.310000 ;
        RECT 59.780000 114.150000 74.290000 114.220000 ;
        RECT 59.780000 137.185000 74.290000 137.255000 ;
        RECT 59.780000 160.200000 74.290000 160.270000 ;
        RECT 59.780000 184.210000 74.290000 184.280000 ;
        RECT 59.795000  81.325000 74.290000  81.395000 ;
        RECT 59.795000 104.325000 74.290000 104.395000 ;
        RECT 59.795000 127.325000 74.290000 127.395000 ;
        RECT 59.795000 150.395000 74.290000 150.465000 ;
        RECT 59.805000  29.580000 74.290000  29.650000 ;
        RECT 59.805000 173.325000 74.290000 173.395000 ;
        RECT 59.835000  58.395000 74.290000  58.465000 ;
        RECT 59.850000  45.080000 74.290000  45.150000 ;
        RECT 59.850000  68.110000 74.290000  68.180000 ;
        RECT 59.850000  91.170000 74.290000  91.240000 ;
        RECT 59.850000 114.080000 74.290000 114.150000 ;
        RECT 59.850000 137.115000 74.290000 137.185000 ;
        RECT 59.850000 160.130000 74.290000 160.200000 ;
        RECT 59.850000 184.140000 74.290000 184.210000 ;
        RECT 59.865000  81.395000 74.290000  81.465000 ;
        RECT 59.865000 104.395000 74.290000 104.465000 ;
        RECT 59.865000 127.395000 74.290000 127.465000 ;
        RECT 59.865000 150.465000 74.290000 150.535000 ;
        RECT 59.875000  29.650000 74.290000  29.720000 ;
        RECT 59.875000 173.395000 74.290000 173.465000 ;
        RECT 59.905000  58.465000 74.290000  58.535000 ;
        RECT 59.920000  45.010000 74.290000  45.080000 ;
        RECT 59.920000  68.040000 74.290000  68.110000 ;
        RECT 59.920000  91.100000 74.290000  91.170000 ;
        RECT 59.920000 114.010000 74.290000 114.080000 ;
        RECT 59.920000 137.045000 74.290000 137.115000 ;
        RECT 59.920000 160.060000 74.290000 160.130000 ;
        RECT 59.920000 184.070000 74.290000 184.140000 ;
        RECT 59.935000  81.465000 74.290000  81.535000 ;
        RECT 59.935000 104.465000 74.290000 104.535000 ;
        RECT 59.935000 127.465000 74.290000 127.535000 ;
        RECT 59.935000 150.535000 74.290000 150.605000 ;
        RECT 59.945000  29.720000 74.290000  29.790000 ;
        RECT 59.945000 173.465000 74.290000 173.535000 ;
        RECT 59.975000  58.535000 74.290000  58.605000 ;
        RECT 59.990000  44.940000 74.290000  45.010000 ;
        RECT 59.990000  67.970000 74.290000  68.040000 ;
        RECT 59.990000  91.030000 74.290000  91.100000 ;
        RECT 59.990000 113.940000 74.290000 114.010000 ;
        RECT 59.990000 136.975000 74.290000 137.045000 ;
        RECT 59.990000 159.990000 74.290000 160.060000 ;
        RECT 59.990000 184.000000 74.290000 184.070000 ;
        RECT 60.005000  81.535000 74.290000  81.605000 ;
        RECT 60.005000 104.535000 74.290000 104.605000 ;
        RECT 60.005000 127.535000 74.290000 127.605000 ;
        RECT 60.005000 150.605000 74.290000 150.675000 ;
        RECT 60.015000  29.790000 74.290000  29.860000 ;
        RECT 60.015000 173.535000 74.290000 173.605000 ;
        RECT 60.045000  58.605000 74.290000  58.675000 ;
        RECT 60.060000  44.870000 74.290000  44.940000 ;
        RECT 60.060000  67.900000 74.290000  67.970000 ;
        RECT 60.060000  90.960000 74.290000  91.030000 ;
        RECT 60.060000 113.870000 74.290000 113.940000 ;
        RECT 60.060000 136.905000 74.290000 136.975000 ;
        RECT 60.060000 159.920000 74.290000 159.990000 ;
        RECT 60.060000 183.930000 74.290000 184.000000 ;
        RECT 60.075000  81.605000 74.290000  81.675000 ;
        RECT 60.075000 104.605000 74.290000 104.675000 ;
        RECT 60.075000 127.605000 74.290000 127.675000 ;
        RECT 60.075000 150.675000 74.290000 150.745000 ;
        RECT 60.085000  29.860000 74.290000  29.930000 ;
        RECT 60.085000 173.605000 74.290000 173.675000 ;
        RECT 60.115000  58.675000 74.290000  58.745000 ;
        RECT 60.130000  44.800000 74.290000  44.870000 ;
        RECT 60.130000  67.830000 74.290000  67.900000 ;
        RECT 60.130000  90.890000 74.290000  90.960000 ;
        RECT 60.130000 113.800000 74.290000 113.870000 ;
        RECT 60.130000 136.835000 74.290000 136.905000 ;
        RECT 60.130000 159.850000 74.290000 159.920000 ;
        RECT 60.130000 183.860000 74.290000 183.930000 ;
        RECT 60.145000  81.675000 74.290000  81.745000 ;
        RECT 60.145000 104.675000 74.290000 104.745000 ;
        RECT 60.145000 127.675000 74.290000 127.745000 ;
        RECT 60.145000 150.745000 74.290000 150.815000 ;
        RECT 60.155000  29.930000 74.290000  30.000000 ;
        RECT 60.155000 173.675000 74.290000 173.745000 ;
        RECT 60.185000  58.745000 74.290000  58.815000 ;
        RECT 60.200000  44.730000 74.290000  44.800000 ;
        RECT 60.200000  67.760000 74.290000  67.830000 ;
        RECT 60.200000  90.820000 74.290000  90.890000 ;
        RECT 60.200000 113.730000 74.290000 113.800000 ;
        RECT 60.200000 136.765000 74.290000 136.835000 ;
        RECT 60.200000 159.780000 74.290000 159.850000 ;
        RECT 60.200000 183.790000 74.290000 183.860000 ;
        RECT 60.215000  81.745000 74.290000  81.815000 ;
        RECT 60.215000 104.745000 74.290000 104.815000 ;
        RECT 60.215000 127.745000 74.290000 127.815000 ;
        RECT 60.215000 150.815000 74.290000 150.885000 ;
        RECT 60.225000  30.000000 74.290000  30.070000 ;
        RECT 60.225000 173.745000 74.290000 173.815000 ;
        RECT 60.255000  58.815000 74.290000  58.885000 ;
        RECT 60.270000  44.660000 74.290000  44.730000 ;
        RECT 60.270000  67.690000 74.290000  67.760000 ;
        RECT 60.270000  90.750000 74.290000  90.820000 ;
        RECT 60.270000 113.660000 74.290000 113.730000 ;
        RECT 60.270000 136.695000 74.290000 136.765000 ;
        RECT 60.270000 159.710000 74.290000 159.780000 ;
        RECT 60.270000 183.720000 74.290000 183.790000 ;
        RECT 60.285000  81.815000 74.290000  81.885000 ;
        RECT 60.285000 104.815000 74.290000 104.885000 ;
        RECT 60.285000 127.815000 74.290000 127.885000 ;
        RECT 60.285000 150.885000 74.290000 150.955000 ;
        RECT 60.295000  30.070000 74.290000  30.140000 ;
        RECT 60.295000 173.815000 74.290000 173.885000 ;
        RECT 60.325000  58.885000 74.290000  58.955000 ;
        RECT 60.340000  44.590000 74.290000  44.660000 ;
        RECT 60.340000  67.620000 74.290000  67.690000 ;
        RECT 60.340000  90.680000 74.290000  90.750000 ;
        RECT 60.340000 113.590000 74.290000 113.660000 ;
        RECT 60.340000 136.625000 74.290000 136.695000 ;
        RECT 60.340000 159.640000 74.290000 159.710000 ;
        RECT 60.340000 183.650000 74.290000 183.720000 ;
        RECT 60.355000  81.885000 74.290000  81.955000 ;
        RECT 60.355000 104.885000 74.290000 104.955000 ;
        RECT 60.355000 127.885000 74.290000 127.955000 ;
        RECT 60.355000 150.955000 74.290000 151.025000 ;
        RECT 60.365000  30.140000 74.290000  30.210000 ;
        RECT 60.365000 173.885000 74.290000 173.955000 ;
        RECT 60.395000  58.955000 74.290000  59.025000 ;
        RECT 60.410000  44.520000 74.290000  44.590000 ;
        RECT 60.410000  67.550000 74.290000  67.620000 ;
        RECT 60.410000  90.610000 74.290000  90.680000 ;
        RECT 60.410000 113.520000 74.290000 113.590000 ;
        RECT 60.410000 136.555000 74.290000 136.625000 ;
        RECT 60.410000 159.570000 74.290000 159.640000 ;
        RECT 60.410000 183.580000 74.290000 183.650000 ;
        RECT 60.425000  81.955000 74.290000  82.025000 ;
        RECT 60.425000 104.955000 74.290000 105.025000 ;
        RECT 60.425000 127.955000 74.290000 128.025000 ;
        RECT 60.425000 151.025000 74.290000 151.095000 ;
        RECT 60.435000  30.210000 74.290000  30.280000 ;
        RECT 60.435000 173.955000 74.290000 174.025000 ;
        RECT 60.465000  59.025000 74.290000  59.095000 ;
        RECT 60.480000  44.450000 74.290000  44.520000 ;
        RECT 60.480000  67.480000 74.290000  67.550000 ;
        RECT 60.480000  90.540000 74.290000  90.610000 ;
        RECT 60.480000 113.450000 74.290000 113.520000 ;
        RECT 60.480000 136.485000 74.290000 136.555000 ;
        RECT 60.480000 159.500000 74.290000 159.570000 ;
        RECT 60.480000 183.510000 74.290000 183.580000 ;
        RECT 60.495000  82.025000 74.290000  82.095000 ;
        RECT 60.495000 105.025000 74.290000 105.095000 ;
        RECT 60.495000 128.025000 74.290000 128.095000 ;
        RECT 60.495000 151.095000 74.290000 151.165000 ;
        RECT 60.505000  30.280000 74.290000  30.350000 ;
        RECT 60.505000 174.025000 74.290000 174.095000 ;
        RECT 60.535000  59.095000 74.290000  59.165000 ;
        RECT 60.550000  44.380000 74.290000  44.450000 ;
        RECT 60.550000  67.410000 74.290000  67.480000 ;
        RECT 60.550000  90.470000 74.290000  90.540000 ;
        RECT 60.550000 113.380000 74.290000 113.450000 ;
        RECT 60.550000 136.415000 74.290000 136.485000 ;
        RECT 60.550000 159.430000 74.290000 159.500000 ;
        RECT 60.550000 183.440000 74.290000 183.510000 ;
        RECT 60.565000  82.095000 74.290000  82.165000 ;
        RECT 60.565000 105.095000 74.290000 105.165000 ;
        RECT 60.565000 128.095000 74.290000 128.165000 ;
        RECT 60.565000 151.165000 74.290000 151.235000 ;
        RECT 60.575000  30.350000 74.290000  30.420000 ;
        RECT 60.575000 174.095000 74.290000 174.165000 ;
        RECT 60.605000  59.165000 74.290000  59.235000 ;
        RECT 60.620000  44.310000 74.290000  44.380000 ;
        RECT 60.620000  67.340000 74.290000  67.410000 ;
        RECT 60.620000  90.400000 74.290000  90.470000 ;
        RECT 60.620000 113.310000 74.290000 113.380000 ;
        RECT 60.620000 136.345000 74.290000 136.415000 ;
        RECT 60.620000 159.360000 74.290000 159.430000 ;
        RECT 60.620000 183.370000 74.290000 183.440000 ;
        RECT 60.635000  82.165000 74.290000  82.235000 ;
        RECT 60.635000 105.165000 74.290000 105.235000 ;
        RECT 60.635000 128.165000 74.290000 128.235000 ;
        RECT 60.635000 151.235000 74.290000 151.305000 ;
        RECT 60.645000  30.420000 74.290000  30.490000 ;
        RECT 60.645000 174.165000 74.290000 174.235000 ;
        RECT 60.675000  59.235000 74.290000  59.305000 ;
        RECT 60.690000  44.240000 74.290000  44.310000 ;
        RECT 60.690000  67.270000 74.290000  67.340000 ;
        RECT 60.690000  90.330000 74.290000  90.400000 ;
        RECT 60.690000 113.240000 74.290000 113.310000 ;
        RECT 60.690000 136.275000 74.290000 136.345000 ;
        RECT 60.690000 159.290000 74.290000 159.360000 ;
        RECT 60.690000 183.300000 74.290000 183.370000 ;
        RECT 60.705000  82.235000 74.290000  82.305000 ;
        RECT 60.705000 105.235000 74.290000 105.305000 ;
        RECT 60.705000 128.235000 74.290000 128.305000 ;
        RECT 60.705000 151.305000 74.290000 151.375000 ;
        RECT 60.715000  30.490000 74.290000  30.560000 ;
        RECT 60.715000 174.235000 74.290000 174.305000 ;
        RECT 60.745000  59.305000 74.290000  59.375000 ;
        RECT 60.760000  44.170000 74.290000  44.240000 ;
        RECT 60.760000  67.200000 74.290000  67.270000 ;
        RECT 60.760000  90.260000 74.290000  90.330000 ;
        RECT 60.760000 113.170000 74.290000 113.240000 ;
        RECT 60.760000 136.205000 74.290000 136.275000 ;
        RECT 60.760000 159.220000 74.290000 159.290000 ;
        RECT 60.760000 183.230000 74.290000 183.300000 ;
        RECT 60.775000  82.305000 74.290000  82.375000 ;
        RECT 60.775000 105.305000 74.290000 105.375000 ;
        RECT 60.775000 128.305000 74.290000 128.375000 ;
        RECT 60.775000 151.375000 74.290000 151.445000 ;
        RECT 60.785000  30.560000 74.290000  30.630000 ;
        RECT 60.785000 174.305000 74.290000 174.375000 ;
        RECT 60.815000  59.375000 74.290000  59.445000 ;
        RECT 60.830000  44.100000 74.290000  44.170000 ;
        RECT 60.830000  67.130000 74.290000  67.200000 ;
        RECT 60.830000  90.190000 74.290000  90.260000 ;
        RECT 60.830000 113.100000 74.290000 113.170000 ;
        RECT 60.830000 136.135000 74.290000 136.205000 ;
        RECT 60.830000 159.150000 74.290000 159.220000 ;
        RECT 60.830000 183.160000 74.290000 183.230000 ;
        RECT 60.845000  82.375000 74.290000  82.445000 ;
        RECT 60.845000 105.375000 74.290000 105.445000 ;
        RECT 60.845000 128.375000 74.290000 128.445000 ;
        RECT 60.845000 151.445000 74.290000 151.515000 ;
        RECT 60.855000  30.630000 74.290000  30.700000 ;
        RECT 60.855000 174.375000 74.290000 174.445000 ;
        RECT 60.885000  59.445000 74.290000  59.515000 ;
        RECT 60.900000  44.030000 74.290000  44.100000 ;
        RECT 60.900000  67.060000 74.290000  67.130000 ;
        RECT 60.900000  90.120000 74.290000  90.190000 ;
        RECT 60.900000 113.030000 74.290000 113.100000 ;
        RECT 60.900000 136.065000 74.290000 136.135000 ;
        RECT 60.900000 159.080000 74.290000 159.150000 ;
        RECT 60.900000 183.090000 74.290000 183.160000 ;
        RECT 60.915000  82.445000 74.290000  82.515000 ;
        RECT 60.915000 105.445000 74.290000 105.515000 ;
        RECT 60.915000 128.445000 74.290000 128.515000 ;
        RECT 60.915000 151.515000 74.290000 151.585000 ;
        RECT 60.925000  30.700000 74.290000  30.770000 ;
        RECT 60.925000 174.445000 74.290000 174.515000 ;
        RECT 60.955000  59.515000 74.290000  59.585000 ;
        RECT 60.970000  43.960000 74.290000  44.030000 ;
        RECT 60.970000  66.990000 74.290000  67.060000 ;
        RECT 60.970000  90.050000 74.290000  90.120000 ;
        RECT 60.970000 112.960000 74.290000 113.030000 ;
        RECT 60.970000 135.995000 74.290000 136.065000 ;
        RECT 60.970000 159.010000 74.290000 159.080000 ;
        RECT 60.970000 183.020000 74.290000 183.090000 ;
        RECT 60.985000  82.515000 74.290000  82.585000 ;
        RECT 60.985000 105.515000 74.290000 105.585000 ;
        RECT 60.985000 128.515000 74.290000 128.585000 ;
        RECT 60.985000 151.585000 74.290000 151.655000 ;
        RECT 60.995000  30.770000 74.290000  30.840000 ;
        RECT 60.995000 174.515000 74.290000 174.585000 ;
        RECT 61.025000  59.585000 74.290000  59.655000 ;
        RECT 61.040000  43.890000 74.290000  43.960000 ;
        RECT 61.040000  66.920000 74.290000  66.990000 ;
        RECT 61.040000  89.980000 74.290000  90.050000 ;
        RECT 61.040000 112.890000 74.290000 112.960000 ;
        RECT 61.040000 135.925000 74.290000 135.995000 ;
        RECT 61.040000 158.940000 74.290000 159.010000 ;
        RECT 61.040000 182.950000 74.290000 183.020000 ;
        RECT 61.055000  82.585000 74.290000  82.655000 ;
        RECT 61.055000 105.585000 74.290000 105.655000 ;
        RECT 61.055000 128.585000 74.290000 128.655000 ;
        RECT 61.055000 151.655000 74.290000 151.725000 ;
        RECT 61.065000  30.840000 74.290000  30.910000 ;
        RECT 61.065000 174.585000 74.290000 174.655000 ;
        RECT 61.095000  59.655000 74.290000  59.725000 ;
        RECT 61.110000  30.910000 74.290000  30.955000 ;
        RECT 61.110000  30.955000 74.290000  43.820000 ;
        RECT 61.110000  43.820000 74.290000  43.890000 ;
        RECT 61.110000  59.725000 74.290000  59.740000 ;
        RECT 61.110000  59.740000 74.290000  66.850000 ;
        RECT 61.110000  66.850000 74.290000  66.920000 ;
        RECT 61.110000  82.655000 74.290000  82.710000 ;
        RECT 61.110000  82.710000 74.290000  89.910000 ;
        RECT 61.110000  89.910000 74.290000  89.980000 ;
        RECT 61.110000 105.655000 74.290000 105.710000 ;
        RECT 61.110000 105.710000 74.290000 112.820000 ;
        RECT 61.110000 112.820000 74.290000 112.890000 ;
        RECT 61.110000 128.655000 74.290000 128.710000 ;
        RECT 61.110000 128.710000 74.290000 135.855000 ;
        RECT 61.110000 135.855000 74.290000 135.925000 ;
        RECT 61.110000 151.725000 74.290000 151.780000 ;
        RECT 61.110000 151.780000 74.290000 158.870000 ;
        RECT 61.110000 158.870000 74.290000 158.940000 ;
        RECT 61.110000 174.655000 74.290000 174.700000 ;
        RECT 61.110000 174.700000 74.290000 182.880000 ;
        RECT 61.110000 182.880000 74.290000 182.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000   0.000000 48.890000  96.150000 ;
        RECT 37.890000  96.150000 48.890000  96.300000 ;
        RECT 37.890000  96.300000 49.040000  96.450000 ;
        RECT 37.890000  96.450000 49.190000  96.600000 ;
        RECT 37.890000  96.600000 49.340000  96.750000 ;
        RECT 37.890000  96.750000 49.490000  96.900000 ;
        RECT 37.890000  96.900000 49.640000  97.050000 ;
        RECT 37.890000  97.050000 49.790000  97.200000 ;
        RECT 37.890000  97.200000 49.940000  97.350000 ;
        RECT 37.890000  97.350000 50.090000  97.500000 ;
        RECT 37.890000  97.500000 50.240000  97.650000 ;
        RECT 37.890000  97.650000 50.390000  97.800000 ;
        RECT 37.890000  97.800000 50.540000  97.950000 ;
        RECT 37.890000  97.950000 50.690000  98.100000 ;
        RECT 37.890000  98.100000 50.840000  98.250000 ;
        RECT 37.890000  98.250000 50.990000  98.300000 ;
        RECT 37.890000  98.300000 51.040000  99.505000 ;
        RECT 37.890000  99.505000 43.400000  99.655000 ;
        RECT 37.890000  99.655000 43.250000  99.805000 ;
        RECT 37.890000  99.805000 43.100000  99.955000 ;
        RECT 37.890000  99.955000 42.950000 100.105000 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
        RECT 37.890000 104.385000 45.090000 104.535000 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
        RECT 38.340000 105.955000 46.660000 106.105000 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
        RECT 40.385000 108.055000 48.760000 108.150000 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
        RECT 42.705000 170.610000 48.855000 170.760000 ;
        RECT 42.785000 110.400000 48.855000 110.550000 ;
        RECT 42.855000 110.550000 48.855000 110.620000 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
        RECT 44.655000  99.505000 51.040000  99.610000 ;
        RECT 44.760000  99.610000 51.040000  99.715000 ;
        RECT 44.910000  99.715000 51.040000  99.865000 ;
        RECT 45.060000  99.865000 51.190000 100.015000 ;
        RECT 45.210000 100.015000 51.340000 100.165000 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
        RECT 47.360000 104.365000 55.690000 104.515000 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
        RECT 48.710000 105.715000 57.040000 105.865000 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
        RECT 49.775000 173.020000 59.285000 173.170000 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
        RECT 49.775000 174.670000 60.935000 174.820000 ;
        RECT 49.775000 174.820000 61.085000 174.970000 ;
        RECT 49.775000 174.970000 61.235000 175.120000 ;
        RECT 49.775000 175.120000 61.385000 175.270000 ;
        RECT 49.775000 175.270000 61.535000 175.420000 ;
        RECT 49.775000 175.420000 61.685000 175.570000 ;
        RECT 49.775000 175.570000 61.835000 175.720000 ;
        RECT 49.775000 175.720000 61.985000 175.870000 ;
        RECT 49.775000 175.870000 62.135000 176.020000 ;
        RECT 49.775000 176.020000 62.285000 176.170000 ;
        RECT 49.775000 176.170000 62.435000 176.320000 ;
        RECT 49.775000 176.320000 62.585000 176.470000 ;
        RECT 49.775000 176.470000 62.735000 176.620000 ;
        RECT 49.775000 176.620000 62.885000 176.770000 ;
        RECT 49.775000 176.770000 63.035000 176.920000 ;
        RECT 49.775000 176.920000 63.185000 177.070000 ;
        RECT 49.775000 177.070000 63.335000 177.220000 ;
        RECT 49.775000 177.220000 63.485000 177.370000 ;
        RECT 49.775000 177.370000 63.635000 177.520000 ;
        RECT 49.775000 177.520000 63.785000 177.670000 ;
        RECT 49.775000 177.670000 63.935000 177.820000 ;
        RECT 49.775000 177.820000 64.085000 177.970000 ;
        RECT 49.775000 177.970000 64.235000 178.120000 ;
        RECT 49.775000 178.120000 64.385000 178.270000 ;
        RECT 49.775000 178.270000 64.535000 178.420000 ;
        RECT 49.775000 178.420000 64.685000 178.570000 ;
        RECT 49.775000 178.570000 64.835000 178.720000 ;
        RECT 49.775000 178.720000 64.985000 178.870000 ;
        RECT 49.775000 178.870000 65.135000 179.020000 ;
        RECT 49.775000 179.020000 65.285000 179.170000 ;
        RECT 49.775000 179.170000 65.435000 179.320000 ;
        RECT 49.775000 179.320000 65.585000 179.470000 ;
        RECT 49.775000 179.470000 65.735000 179.620000 ;
        RECT 49.775000 179.620000 65.885000 179.770000 ;
        RECT 49.775000 179.770000 66.035000 179.920000 ;
        RECT 49.775000 179.920000 66.185000 180.070000 ;
        RECT 49.775000 180.070000 66.335000 180.220000 ;
        RECT 49.775000 180.220000 66.485000 180.370000 ;
        RECT 49.775000 180.370000 66.635000 180.520000 ;
        RECT 49.775000 180.520000 66.785000 180.670000 ;
        RECT 49.775000 180.670000 66.935000 180.820000 ;
        RECT 49.775000 180.820000 67.085000 180.970000 ;
        RECT 49.775000 180.970000 67.235000 181.120000 ;
        RECT 49.775000 181.120000 67.385000 181.270000 ;
        RECT 49.775000 181.270000 67.535000 181.420000 ;
        RECT 49.775000 181.420000 67.685000 181.570000 ;
        RECT 49.775000 181.570000 67.835000 181.720000 ;
        RECT 49.775000 181.720000 67.985000 181.870000 ;
        RECT 49.775000 181.870000 68.135000 182.020000 ;
        RECT 49.775000 182.020000 68.285000 182.170000 ;
        RECT 49.775000 182.170000 68.435000 182.320000 ;
        RECT 49.775000 182.320000 68.585000 182.470000 ;
        RECT 49.775000 182.470000 68.735000 182.620000 ;
        RECT 49.775000 182.620000 68.885000 182.770000 ;
        RECT 49.775000 182.770000 69.035000 182.920000 ;
        RECT 49.775000 182.920000 69.185000 183.070000 ;
        RECT 49.775000 183.070000 69.335000 183.220000 ;
        RECT 49.775000 183.220000 69.485000 183.370000 ;
        RECT 49.775000 183.370000 69.635000 183.520000 ;
        RECT 49.775000 183.520000 69.785000 183.670000 ;
        RECT 49.775000 183.670000 69.935000 183.820000 ;
        RECT 49.775000 183.820000 70.085000 183.970000 ;
        RECT 49.775000 183.970000 70.235000 184.120000 ;
        RECT 49.775000 184.120000 70.385000 184.270000 ;
        RECT 49.775000 184.270000 70.535000 184.420000 ;
        RECT 49.775000 184.420000 70.685000 184.570000 ;
        RECT 49.775000 184.570000 70.835000 184.720000 ;
        RECT 49.775000 184.720000 70.985000 184.870000 ;
        RECT 49.775000 184.870000 71.135000 185.020000 ;
        RECT 49.775000 185.020000 71.285000 185.170000 ;
        RECT 49.775000 185.170000 71.435000 185.320000 ;
        RECT 49.775000 185.320000 71.585000 185.360000 ;
        RECT 49.775000 185.360000 71.625000 190.040000 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
        RECT 50.805000 107.815000 59.140000 107.960000 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
        RECT 50.955000 107.960000 59.285000 108.110000 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
        RECT 53.135000 169.285000 59.285000 169.435000 ;
        RECT 53.205000 110.210000 59.285000 110.360000 ;
        RECT 53.285000 110.360000 59.285000 110.440000 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
  END DRN_HVC
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000   0.000000 24.395000  36.510000 ;
        RECT 0.495000  46.960000 24.395000  90.500000 ;
        RECT 0.495000  90.500000 24.245000  90.650000 ;
        RECT 0.495000  90.650000 24.095000  90.800000 ;
        RECT 0.495000  90.800000 23.945000  90.950000 ;
        RECT 0.495000  90.950000 23.795000  91.100000 ;
        RECT 0.495000  91.100000 23.645000  91.250000 ;
        RECT 0.495000  91.250000 23.495000  91.400000 ;
        RECT 0.495000  91.400000 23.345000  91.550000 ;
        RECT 0.495000  91.550000 23.195000  91.700000 ;
        RECT 0.495000  91.700000 23.045000  91.850000 ;
        RECT 0.495000  91.850000 22.895000  92.000000 ;
        RECT 0.495000  92.000000 22.745000  92.150000 ;
        RECT 0.495000  92.150000 22.595000  92.300000 ;
        RECT 0.495000  92.300000 22.445000  92.450000 ;
        RECT 0.495000  92.450000 22.295000  92.600000 ;
        RECT 0.495000  92.600000 22.145000  92.750000 ;
        RECT 0.495000  92.750000 21.995000  92.900000 ;
        RECT 0.495000  92.900000 21.845000  93.050000 ;
        RECT 0.495000  93.050000 21.695000  93.200000 ;
        RECT 0.495000  93.200000 21.545000  93.350000 ;
        RECT 0.495000  93.350000 21.395000  93.500000 ;
        RECT 0.495000  93.500000 21.245000  93.650000 ;
        RECT 0.495000  93.650000 21.095000  93.800000 ;
        RECT 0.495000  93.800000 20.945000  93.950000 ;
        RECT 0.495000  93.950000 20.795000  94.100000 ;
        RECT 0.495000  94.100000 20.645000  94.250000 ;
        RECT 0.495000  94.250000 20.495000  94.400000 ;
        RECT 0.495000  94.400000 20.345000  94.550000 ;
        RECT 0.495000  94.550000 20.195000  94.700000 ;
        RECT 0.495000  94.700000 20.045000  94.850000 ;
        RECT 0.495000  94.850000 19.895000  95.000000 ;
        RECT 0.495000  95.000000 19.745000  95.150000 ;
        RECT 0.495000  95.150000 19.595000  95.300000 ;
        RECT 0.495000  95.300000 19.445000  95.450000 ;
        RECT 0.495000  95.450000 19.295000  95.600000 ;
        RECT 0.495000  95.600000 19.145000  95.750000 ;
        RECT 0.495000  95.750000 18.995000  95.900000 ;
        RECT 0.495000  95.900000 18.845000  96.050000 ;
        RECT 0.495000  96.050000 18.695000  96.200000 ;
        RECT 0.495000  96.200000 18.545000  96.350000 ;
        RECT 0.495000  96.350000 18.395000  96.500000 ;
        RECT 0.495000  96.500000 18.245000  96.650000 ;
        RECT 0.495000  96.650000 18.095000  96.800000 ;
        RECT 0.495000  96.800000 17.945000  96.950000 ;
        RECT 0.495000  96.950000 17.795000  97.100000 ;
        RECT 0.495000  97.100000 17.645000  97.250000 ;
        RECT 0.495000  97.250000 17.495000  97.400000 ;
        RECT 0.495000  97.400000 17.345000  97.550000 ;
        RECT 0.495000  97.550000 17.195000  97.700000 ;
        RECT 0.495000  97.700000 17.045000  97.850000 ;
        RECT 0.495000  97.850000 16.895000  98.000000 ;
        RECT 0.495000  98.000000 16.745000  98.150000 ;
        RECT 0.495000  98.150000 16.595000  98.300000 ;
        RECT 0.495000  98.300000 16.445000  98.450000 ;
        RECT 0.495000  98.450000 16.295000  98.600000 ;
        RECT 0.495000  98.600000 16.145000  98.750000 ;
        RECT 0.495000  98.750000 15.995000  98.900000 ;
        RECT 0.495000  98.900000 15.845000  99.050000 ;
        RECT 0.495000  99.050000 15.695000  99.200000 ;
        RECT 0.495000  99.200000 15.545000  99.350000 ;
        RECT 0.495000  99.350000 15.395000  99.500000 ;
        RECT 0.495000  99.500000 15.245000  99.650000 ;
        RECT 0.495000  99.650000 15.095000  99.800000 ;
        RECT 0.495000  99.800000 14.945000  99.950000 ;
        RECT 0.495000  99.950000 14.795000 100.100000 ;
        RECT 0.495000 100.100000 14.645000 100.250000 ;
        RECT 0.495000 100.250000 14.495000 100.400000 ;
        RECT 0.495000 100.400000 14.345000 100.550000 ;
        RECT 0.495000 100.550000 14.195000 100.700000 ;
        RECT 0.495000 100.700000 14.045000 100.850000 ;
        RECT 0.495000 100.850000 13.895000 101.000000 ;
        RECT 0.495000 101.000000 13.745000 101.150000 ;
        RECT 0.495000 101.150000 13.595000 101.300000 ;
        RECT 0.495000 101.300000 13.500000 101.395000 ;
        RECT 0.495000 101.395000 13.500000 173.155000 ;
        RECT 0.510000  46.945000 24.395000  46.960000 ;
        RECT 0.645000  36.510000 24.395000  36.660000 ;
        RECT 0.660000  46.795000 24.395000  46.945000 ;
        RECT 0.795000  36.660000 24.395000  36.810000 ;
        RECT 0.810000  46.645000 24.395000  46.795000 ;
        RECT 0.945000  36.810000 24.395000  36.960000 ;
        RECT 0.960000  46.495000 24.395000  46.645000 ;
        RECT 1.095000  36.960000 24.395000  37.110000 ;
        RECT 1.110000  37.110000 24.395000  37.125000 ;
        RECT 1.110000  37.125000 24.395000  46.345000 ;
        RECT 1.110000  46.345000 24.395000  46.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000   0.000000 74.290000  90.185000 ;
        RECT 50.540000  90.185000 74.290000  90.335000 ;
        RECT 50.690000  90.335000 74.290000  90.485000 ;
        RECT 50.840000  90.485000 74.290000  90.635000 ;
        RECT 50.990000  90.635000 74.290000  90.785000 ;
        RECT 51.140000  90.785000 74.290000  90.935000 ;
        RECT 51.290000  90.935000 74.290000  91.085000 ;
        RECT 51.440000  91.085000 74.290000  91.235000 ;
        RECT 51.590000  91.235000 74.290000  91.385000 ;
        RECT 51.740000  91.385000 74.290000  91.535000 ;
        RECT 51.890000  91.535000 74.290000  91.685000 ;
        RECT 52.040000  91.685000 74.290000  91.835000 ;
        RECT 52.190000  91.835000 74.290000  91.985000 ;
        RECT 52.340000  91.985000 74.290000  92.135000 ;
        RECT 52.490000  92.135000 74.290000  92.285000 ;
        RECT 52.640000  92.285000 74.290000  92.435000 ;
        RECT 52.790000  92.435000 74.290000  92.585000 ;
        RECT 52.940000  92.585000 74.290000  92.735000 ;
        RECT 53.090000  92.735000 74.290000  92.885000 ;
        RECT 53.240000  92.885000 74.290000  93.035000 ;
        RECT 53.390000  93.035000 74.290000  93.185000 ;
        RECT 53.540000  93.185000 74.290000  93.335000 ;
        RECT 53.690000  93.335000 74.290000  93.485000 ;
        RECT 53.840000  93.485000 74.290000  93.635000 ;
        RECT 53.990000  93.635000 74.290000  93.785000 ;
        RECT 54.140000  93.785000 74.290000  93.935000 ;
        RECT 54.290000  93.935000 74.290000  94.085000 ;
        RECT 54.440000  94.085000 74.290000  94.235000 ;
        RECT 54.590000  94.235000 74.290000  94.385000 ;
        RECT 54.740000  94.385000 74.290000  94.535000 ;
        RECT 54.890000  94.535000 74.290000  94.685000 ;
        RECT 55.040000  94.685000 74.290000  94.835000 ;
        RECT 55.190000  94.835000 74.290000  94.985000 ;
        RECT 55.340000  94.985000 74.290000  95.135000 ;
        RECT 55.490000  95.135000 74.290000  95.285000 ;
        RECT 55.640000  95.285000 74.290000  95.435000 ;
        RECT 55.790000  95.435000 74.290000  95.585000 ;
        RECT 55.940000  95.585000 74.290000  95.735000 ;
        RECT 56.090000  95.735000 74.290000  95.885000 ;
        RECT 56.240000  95.885000 74.290000  96.035000 ;
        RECT 56.390000  96.035000 74.290000  96.185000 ;
        RECT 56.540000  96.185000 74.290000  96.335000 ;
        RECT 56.690000  96.335000 74.290000  96.485000 ;
        RECT 56.840000  96.485000 74.290000  96.635000 ;
        RECT 56.990000  96.635000 74.290000  96.785000 ;
        RECT 57.140000  96.785000 74.290000  96.935000 ;
        RECT 57.290000  96.935000 74.290000  97.085000 ;
        RECT 57.440000  97.085000 74.290000  97.235000 ;
        RECT 57.590000  97.235000 74.290000  97.385000 ;
        RECT 57.740000  97.385000 74.290000  97.535000 ;
        RECT 57.890000  97.535000 74.290000  97.685000 ;
        RECT 58.040000  97.685000 74.290000  97.835000 ;
        RECT 58.190000  97.835000 74.290000  97.985000 ;
        RECT 58.340000  97.985000 74.290000  98.135000 ;
        RECT 58.490000  98.135000 74.290000  98.285000 ;
        RECT 58.640000  98.285000 74.290000  98.435000 ;
        RECT 58.790000  98.435000 74.290000  98.585000 ;
        RECT 58.940000  98.585000 74.290000  98.735000 ;
        RECT 59.090000  98.735000 74.290000  98.885000 ;
        RECT 59.240000  98.885000 74.290000  99.035000 ;
        RECT 59.390000  99.035000 74.290000  99.185000 ;
        RECT 59.540000  99.185000 74.290000  99.335000 ;
        RECT 59.690000  99.335000 74.290000  99.485000 ;
        RECT 59.840000  99.485000 74.290000  99.635000 ;
        RECT 59.990000  99.635000 74.290000  99.785000 ;
        RECT 60.140000  99.785000 74.290000  99.935000 ;
        RECT 60.290000  99.935000 74.290000 100.085000 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
        RECT 61.490000 101.135000 74.290000 101.285000 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END P_CORE
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.495000   0.000000 24.395000   2.055000 ;
        RECT  0.565000   2.055000 24.395000   2.125000 ;
        RECT  0.635000   2.125000 24.395000   2.195000 ;
        RECT  0.705000   2.195000 24.395000   2.265000 ;
        RECT  0.775000   2.265000 24.395000   2.335000 ;
        RECT  0.845000   2.335000 24.395000   2.405000 ;
        RECT  0.915000   2.405000 24.395000   2.475000 ;
        RECT  0.985000   2.475000 24.395000   2.545000 ;
        RECT  1.005000   2.545000 24.395000   2.565000 ;
        RECT  1.005000   2.565000 24.395000   8.595000 ;
        RECT  1.005000   8.595000 24.395000   8.665000 ;
        RECT  1.005000   8.665000 24.465000   8.735000 ;
        RECT  1.005000   8.735000 24.535000   8.805000 ;
        RECT  1.005000   8.805000 24.605000   8.875000 ;
        RECT  1.005000   8.875000 24.675000   8.945000 ;
        RECT  1.005000   8.945000 24.745000   9.015000 ;
        RECT  1.005000   9.015000 24.815000   9.085000 ;
        RECT  1.005000   9.085000 24.885000   9.155000 ;
        RECT  1.005000   9.155000 24.955000   9.225000 ;
        RECT  1.005000   9.225000 25.025000   9.295000 ;
        RECT  1.005000   9.295000 25.095000   9.365000 ;
        RECT  1.005000   9.365000 25.165000   9.435000 ;
        RECT  1.005000   9.435000 25.235000   9.505000 ;
        RECT  1.005000   9.505000 25.305000   9.575000 ;
        RECT  1.005000   9.575000 25.375000   9.645000 ;
        RECT  1.005000   9.645000 25.445000   9.715000 ;
        RECT  1.005000   9.715000 25.515000   9.785000 ;
        RECT  1.005000   9.785000 25.585000   9.855000 ;
        RECT  1.005000   9.855000 25.655000   9.925000 ;
        RECT  1.005000   9.925000 25.725000   9.995000 ;
        RECT  1.005000   9.995000 25.795000  10.065000 ;
        RECT  1.005000  10.065000 25.865000  10.135000 ;
        RECT  1.005000  10.135000 25.935000  10.205000 ;
        RECT  1.005000  10.205000 26.005000  10.275000 ;
        RECT  1.005000  10.275000 26.075000  10.345000 ;
        RECT  1.005000  10.345000 26.145000  10.415000 ;
        RECT  1.005000  10.415000 26.215000  10.485000 ;
        RECT  1.005000  10.485000 26.285000  10.555000 ;
        RECT  1.005000  10.555000 26.355000  10.625000 ;
        RECT  1.005000  10.625000 26.425000  10.695000 ;
        RECT  1.005000  10.695000 26.495000  10.765000 ;
        RECT  1.005000  10.765000 26.565000  10.835000 ;
        RECT  1.005000  10.835000 26.635000  10.905000 ;
        RECT  1.005000  10.905000 26.705000  10.975000 ;
        RECT  1.005000  10.975000 26.775000  11.045000 ;
        RECT  1.005000  11.045000 26.845000  11.115000 ;
        RECT  1.005000  11.115000 26.915000  11.185000 ;
        RECT  1.005000  11.185000 26.985000  11.255000 ;
        RECT  1.005000  11.255000 27.055000  11.325000 ;
        RECT  1.005000  11.325000 27.125000  11.395000 ;
        RECT  1.005000  11.395000 27.195000  11.465000 ;
        RECT  1.005000  11.465000 27.265000  11.535000 ;
        RECT  1.005000  11.535000 27.335000  11.605000 ;
        RECT  1.005000  11.605000 27.405000  11.675000 ;
        RECT  1.005000  11.675000 27.475000  11.745000 ;
        RECT  1.005000  11.745000 27.545000  11.815000 ;
        RECT  1.005000  11.815000 27.615000  11.885000 ;
        RECT  1.005000  11.885000 27.685000  11.955000 ;
        RECT  1.005000  11.955000 27.755000  12.025000 ;
        RECT  1.005000  12.025000 27.825000  12.095000 ;
        RECT  1.005000  12.095000 27.895000  12.165000 ;
        RECT  1.005000  12.165000 27.965000  12.235000 ;
        RECT  1.005000  12.235000 28.035000  12.305000 ;
        RECT  1.005000  12.305000 28.105000  12.375000 ;
        RECT  1.005000  12.375000 28.175000  12.400000 ;
        RECT  1.005000  12.400000 36.895000  25.700000 ;
        RECT  1.005000  25.700000 18.750000  25.770000 ;
        RECT  1.005000  25.770000 18.680000  25.840000 ;
        RECT  1.005000  25.840000 18.610000  25.910000 ;
        RECT  1.005000  25.910000 18.540000  25.980000 ;
        RECT  1.005000  25.980000 18.470000  26.050000 ;
        RECT  1.005000  26.050000 18.400000  26.120000 ;
        RECT  1.005000  26.120000 18.330000  26.190000 ;
        RECT  1.005000  26.190000 18.260000  26.260000 ;
        RECT  1.005000  26.260000 18.190000  26.330000 ;
        RECT  1.005000  26.330000 18.120000  26.400000 ;
        RECT  1.005000  26.400000 18.050000  26.470000 ;
        RECT  1.005000  26.470000 17.980000  26.540000 ;
        RECT  1.005000  26.540000 17.910000  26.610000 ;
        RECT  1.005000  26.610000 17.840000  26.680000 ;
        RECT  1.005000  26.680000 17.770000  26.750000 ;
        RECT  1.005000  26.750000 17.700000  26.820000 ;
        RECT  1.005000  26.820000 17.630000  26.890000 ;
        RECT  1.005000  26.890000 17.560000  26.960000 ;
        RECT  1.005000  26.960000 17.490000  27.030000 ;
        RECT  1.005000  27.030000 17.420000  27.100000 ;
        RECT  1.005000  27.100000 17.350000  27.170000 ;
        RECT  1.005000  27.170000 17.280000  27.240000 ;
        RECT  1.005000  27.240000 17.210000  27.310000 ;
        RECT  1.005000  27.310000 17.140000  27.380000 ;
        RECT  1.005000  27.380000 17.070000  27.450000 ;
        RECT  1.005000  27.450000 17.000000  27.520000 ;
        RECT  1.005000  27.520000 16.930000  27.590000 ;
        RECT  1.005000  27.590000 16.860000  27.660000 ;
        RECT  1.005000  27.660000 16.790000  27.730000 ;
        RECT  1.005000  27.730000 16.720000  27.800000 ;
        RECT  1.005000  27.800000 16.650000  27.870000 ;
        RECT  1.005000  27.870000 16.580000  27.940000 ;
        RECT  1.005000  27.940000 16.510000  28.010000 ;
        RECT  1.005000  28.010000 16.440000  28.080000 ;
        RECT  1.005000  28.080000 16.370000  28.150000 ;
        RECT  1.005000  28.150000 16.300000  28.220000 ;
        RECT  1.005000  28.220000 16.230000  28.290000 ;
        RECT  1.005000  28.290000 16.160000  28.360000 ;
        RECT  1.005000  28.360000 16.090000  28.430000 ;
        RECT  1.005000  28.430000 16.020000  28.500000 ;
        RECT  1.005000  28.500000 15.950000  28.570000 ;
        RECT  1.005000  28.570000 15.880000  28.640000 ;
        RECT  1.005000  28.640000 15.810000  28.710000 ;
        RECT  1.005000  28.710000 15.740000  28.780000 ;
        RECT  1.005000  28.780000 15.670000  28.850000 ;
        RECT  1.005000  28.850000 15.600000  28.920000 ;
        RECT  1.005000  28.920000 15.530000  28.990000 ;
        RECT  1.005000  28.990000 15.460000  29.060000 ;
        RECT  1.005000  29.060000 15.390000  29.130000 ;
        RECT  1.005000  29.130000 15.320000  29.200000 ;
        RECT  1.005000  29.200000 15.250000  29.270000 ;
        RECT  1.005000  29.270000 15.205000  29.315000 ;
        RECT  1.005000  29.315000 15.205000  35.665000 ;
        RECT  1.005000  35.665000 15.205000  35.735000 ;
        RECT  1.005000  35.735000 15.275000  35.805000 ;
        RECT  1.005000  35.805000 15.345000  35.875000 ;
        RECT  1.005000  35.875000 15.415000  35.945000 ;
        RECT  1.005000  35.945000 15.485000  36.015000 ;
        RECT  1.005000  36.015000 15.555000  36.085000 ;
        RECT  1.005000  36.085000 15.625000  36.155000 ;
        RECT  1.005000  36.155000 15.695000  36.225000 ;
        RECT  1.005000  36.225000 15.765000  36.295000 ;
        RECT  1.005000  36.295000 15.835000  36.365000 ;
        RECT  1.005000  36.365000 15.905000  36.435000 ;
        RECT  1.005000  36.435000 15.975000  36.505000 ;
        RECT  1.005000  36.505000 16.045000  36.575000 ;
        RECT  1.005000  36.575000 16.115000  36.645000 ;
        RECT  1.005000  36.645000 16.185000  36.715000 ;
        RECT  1.005000  36.715000 16.255000  36.785000 ;
        RECT  1.005000  36.785000 16.325000  36.855000 ;
        RECT  1.005000  47.100000 14.120000  54.215000 ;
        RECT  1.005000  54.215000 14.120000  54.285000 ;
        RECT  1.005000  54.285000 14.190000  54.355000 ;
        RECT  1.005000  54.355000 14.260000  54.425000 ;
        RECT  1.005000  54.425000 14.330000  54.495000 ;
        RECT  1.005000  54.495000 14.400000  54.565000 ;
        RECT  1.005000  54.565000 14.470000  54.635000 ;
        RECT  1.005000  54.635000 14.540000  54.705000 ;
        RECT  1.005000  54.705000 14.610000  54.775000 ;
        RECT  1.005000  54.775000 14.680000  54.845000 ;
        RECT  1.005000  54.845000 14.750000  54.915000 ;
        RECT  1.005000  54.915000 14.820000  54.985000 ;
        RECT  1.005000  54.985000 14.890000  55.055000 ;
        RECT  1.005000  55.055000 14.960000  55.125000 ;
        RECT  1.005000  55.125000 15.030000  55.195000 ;
        RECT  1.005000  55.195000 15.100000  55.265000 ;
        RECT  1.005000  55.265000 15.170000  55.335000 ;
        RECT  1.005000  55.335000 15.240000  55.405000 ;
        RECT  1.005000  55.405000 15.310000  55.475000 ;
        RECT  1.005000  55.475000 15.380000  55.545000 ;
        RECT  1.005000  55.545000 15.450000  55.615000 ;
        RECT  1.005000  55.615000 15.520000  55.685000 ;
        RECT  1.005000  55.685000 15.590000  55.755000 ;
        RECT  1.005000  55.755000 15.660000  55.825000 ;
        RECT  1.005000  55.825000 15.730000  55.895000 ;
        RECT  1.005000  55.895000 15.800000  55.965000 ;
        RECT  1.005000  55.965000 15.870000  56.035000 ;
        RECT  1.005000  56.035000 15.940000  56.105000 ;
        RECT  1.005000  56.105000 16.010000  56.175000 ;
        RECT  1.005000  56.175000 16.080000  56.245000 ;
        RECT  1.005000  56.245000 16.150000  56.315000 ;
        RECT  1.005000  56.315000 16.220000  56.385000 ;
        RECT  1.005000  56.385000 16.290000  56.455000 ;
        RECT  1.005000  56.455000 16.360000  56.525000 ;
        RECT  1.005000  56.525000 16.430000  56.595000 ;
        RECT  1.005000  56.595000 16.500000  56.665000 ;
        RECT  1.005000  56.665000 16.570000  56.735000 ;
        RECT  1.005000  56.735000 16.640000  56.805000 ;
        RECT  1.005000  56.805000 16.710000  56.875000 ;
        RECT  1.005000  56.875000 16.780000  56.945000 ;
        RECT  1.005000  56.945000 16.850000  57.015000 ;
        RECT  1.005000  57.015000 16.920000  57.085000 ;
        RECT  1.005000  57.085000 16.990000  57.155000 ;
        RECT  1.005000  57.155000 17.060000  57.225000 ;
        RECT  1.005000  57.225000 17.130000  57.295000 ;
        RECT  1.005000  57.295000 17.200000  57.365000 ;
        RECT  1.005000  57.365000 17.270000  57.435000 ;
        RECT  1.005000  57.435000 17.340000  57.505000 ;
        RECT  1.005000  57.505000 17.410000  57.575000 ;
        RECT  1.005000  57.575000 17.480000  57.645000 ;
        RECT  1.005000  57.645000 17.550000  57.715000 ;
        RECT  1.005000  57.715000 17.620000  57.780000 ;
        RECT  1.005000  57.780000 56.710000  66.480000 ;
        RECT  1.005000  66.480000 17.595000  66.550000 ;
        RECT  1.005000  66.550000 17.525000  66.620000 ;
        RECT  1.005000  66.620000 17.455000  66.690000 ;
        RECT  1.005000  66.690000 17.385000  66.760000 ;
        RECT  1.005000  66.760000 17.315000  66.830000 ;
        RECT  1.005000  66.830000 17.245000  66.900000 ;
        RECT  1.005000  66.900000 17.175000  66.970000 ;
        RECT  1.005000  66.970000 17.105000  67.040000 ;
        RECT  1.005000  67.040000 17.035000  67.110000 ;
        RECT  1.005000  67.110000 16.965000  67.180000 ;
        RECT  1.005000  67.180000 16.895000  67.250000 ;
        RECT  1.005000  67.250000 16.825000  67.320000 ;
        RECT  1.005000  67.320000 16.755000  67.390000 ;
        RECT  1.005000  67.390000 16.685000  67.460000 ;
        RECT  1.005000  67.460000 16.615000  67.530000 ;
        RECT  1.005000  67.530000 16.545000  67.600000 ;
        RECT  1.005000  67.600000 16.475000  67.670000 ;
        RECT  1.005000  67.670000 16.405000  67.740000 ;
        RECT  1.005000  67.740000 16.335000  67.810000 ;
        RECT  1.005000  67.810000 16.265000  67.880000 ;
        RECT  1.005000  67.880000 16.195000  67.950000 ;
        RECT  1.005000  67.950000 16.125000  68.020000 ;
        RECT  1.005000  68.020000 16.055000  68.090000 ;
        RECT  1.005000  68.090000 15.985000  68.160000 ;
        RECT  1.005000  68.160000 15.915000  68.230000 ;
        RECT  1.005000  68.230000 15.845000  68.300000 ;
        RECT  1.005000  68.300000 15.775000  68.370000 ;
        RECT  1.005000  68.370000 15.705000  68.440000 ;
        RECT  1.005000  68.440000 15.635000  68.510000 ;
        RECT  1.005000  68.510000 15.565000  68.580000 ;
        RECT  1.005000  68.580000 15.495000  68.650000 ;
        RECT  1.005000  68.650000 15.425000  68.720000 ;
        RECT  1.005000  68.720000 15.355000  68.790000 ;
        RECT  1.005000  68.790000 15.285000  68.860000 ;
        RECT  1.005000  68.860000 15.215000  68.930000 ;
        RECT  1.005000  68.930000 15.145000  69.000000 ;
        RECT  1.005000  69.000000 15.075000  69.070000 ;
        RECT  1.005000  69.070000 15.005000  69.140000 ;
        RECT  1.005000  69.140000 14.935000  69.210000 ;
        RECT  1.005000  69.210000 14.865000  69.280000 ;
        RECT  1.005000  69.280000 14.795000  69.350000 ;
        RECT  1.005000  69.350000 14.725000  69.420000 ;
        RECT  1.005000  69.420000 14.655000  69.490000 ;
        RECT  1.005000  69.490000 14.585000  69.560000 ;
        RECT  1.005000  69.560000 14.515000  69.630000 ;
        RECT  1.005000  69.630000 14.445000  69.700000 ;
        RECT  1.005000  69.700000 14.375000  69.770000 ;
        RECT  1.005000  69.770000 14.305000  69.840000 ;
        RECT  1.005000  69.840000 14.235000  69.910000 ;
        RECT  1.005000  69.910000 14.165000  69.980000 ;
        RECT  1.005000  69.980000 14.120000  70.025000 ;
        RECT  1.005000  70.025000 14.120000  77.240000 ;
        RECT  1.005000  77.240000 14.120000  77.310000 ;
        RECT  1.005000  77.310000 14.190000  77.380000 ;
        RECT  1.005000  77.380000 14.260000  77.450000 ;
        RECT  1.005000  77.450000 14.330000  77.520000 ;
        RECT  1.005000  77.520000 14.400000  77.590000 ;
        RECT  1.005000  77.590000 14.470000  77.660000 ;
        RECT  1.005000  77.660000 14.540000  77.730000 ;
        RECT  1.005000  77.730000 14.610000  77.800000 ;
        RECT  1.005000  77.800000 14.680000  77.870000 ;
        RECT  1.005000  77.870000 14.750000  77.940000 ;
        RECT  1.005000  77.940000 14.820000  78.010000 ;
        RECT  1.005000  78.010000 14.890000  78.080000 ;
        RECT  1.005000  78.080000 14.960000  78.150000 ;
        RECT  1.005000  78.150000 15.030000  78.220000 ;
        RECT  1.005000  78.220000 15.100000  78.290000 ;
        RECT  1.005000  78.290000 15.170000  78.360000 ;
        RECT  1.005000  78.360000 15.240000  78.430000 ;
        RECT  1.005000  78.430000 15.310000  78.500000 ;
        RECT  1.005000  78.500000 15.380000  78.570000 ;
        RECT  1.005000  78.570000 15.450000  78.640000 ;
        RECT  1.005000  78.640000 15.520000  78.710000 ;
        RECT  1.005000  78.710000 15.590000  78.780000 ;
        RECT  1.005000  78.780000 15.660000  78.850000 ;
        RECT  1.005000  78.850000 15.730000  78.920000 ;
        RECT  1.005000  78.920000 15.800000  78.990000 ;
        RECT  1.005000  78.990000 15.870000  79.060000 ;
        RECT  1.005000  79.060000 15.940000  79.130000 ;
        RECT  1.005000  79.130000 16.010000  79.200000 ;
        RECT  1.005000  79.200000 16.080000  79.270000 ;
        RECT  1.005000  79.270000 16.150000  79.340000 ;
        RECT  1.005000  79.340000 16.220000  79.410000 ;
        RECT  1.005000  79.410000 16.290000  79.480000 ;
        RECT  1.005000  79.480000 16.360000  79.550000 ;
        RECT  1.005000  79.550000 16.430000  79.620000 ;
        RECT  1.005000  79.620000 16.500000  79.690000 ;
        RECT  1.005000  79.690000 16.570000  79.760000 ;
        RECT  1.005000  79.760000 16.640000  79.830000 ;
        RECT  1.005000  79.830000 16.710000  79.900000 ;
        RECT  1.005000  79.900000 16.780000  79.970000 ;
        RECT  1.005000  79.970000 16.850000  80.040000 ;
        RECT  1.005000  80.040000 16.920000  80.110000 ;
        RECT  1.005000  80.110000 16.990000  80.180000 ;
        RECT  1.005000  80.180000 17.060000  80.250000 ;
        RECT  1.005000  80.250000 17.130000  80.320000 ;
        RECT  1.005000  80.320000 17.200000  80.390000 ;
        RECT  1.005000  80.390000 17.270000  80.460000 ;
        RECT  1.005000  80.460000 17.340000  80.530000 ;
        RECT  1.005000  80.530000 17.410000  80.600000 ;
        RECT  1.005000  80.600000 17.480000  80.670000 ;
        RECT  1.005000  80.670000 17.550000  80.740000 ;
        RECT  1.005000  80.740000 17.620000  80.780000 ;
        RECT  1.005000  80.780000 56.705000  89.480000 ;
        RECT  1.005000  89.480000 17.595000  89.550000 ;
        RECT  1.005000  89.550000 17.525000  89.620000 ;
        RECT  1.005000  89.620000 17.455000  89.690000 ;
        RECT  1.005000  89.690000 17.385000  89.760000 ;
        RECT  1.005000  89.760000 17.315000  89.830000 ;
        RECT  1.005000  89.830000 17.245000  89.900000 ;
        RECT  1.005000  89.900000 17.175000  89.970000 ;
        RECT  1.005000  89.970000 17.105000  90.040000 ;
        RECT  1.005000  90.040000 17.035000  90.110000 ;
        RECT  1.005000  90.110000 16.965000  90.180000 ;
        RECT  1.005000  90.180000 16.895000  90.250000 ;
        RECT  1.005000  90.250000 16.825000  90.320000 ;
        RECT  1.005000  90.320000 16.755000  90.390000 ;
        RECT  1.005000  90.390000 16.685000  90.460000 ;
        RECT  1.005000  90.460000 16.615000  90.530000 ;
        RECT  1.005000  90.530000 16.545000  90.600000 ;
        RECT  1.005000  90.600000 16.475000  90.670000 ;
        RECT  1.005000  90.670000 16.405000  90.740000 ;
        RECT  1.005000  90.740000 16.335000  90.810000 ;
        RECT  1.005000  90.810000 16.265000  90.880000 ;
        RECT  1.005000  90.880000 16.195000  90.950000 ;
        RECT  1.005000  90.950000 16.125000  91.020000 ;
        RECT  1.005000  91.020000 16.055000  91.090000 ;
        RECT  1.005000  91.090000 15.985000  91.160000 ;
        RECT  1.005000  91.160000 15.915000  91.230000 ;
        RECT  1.005000  91.230000 15.845000  91.300000 ;
        RECT  1.005000  91.300000 15.775000  91.370000 ;
        RECT  1.005000  91.370000 15.705000  91.440000 ;
        RECT  1.005000  91.440000 15.635000  91.510000 ;
        RECT  1.005000  91.510000 15.565000  91.580000 ;
        RECT  1.005000  91.580000 15.495000  91.650000 ;
        RECT  1.005000  91.650000 15.425000  91.720000 ;
        RECT  1.005000  91.720000 15.355000  91.790000 ;
        RECT  1.005000  91.790000 15.285000  91.860000 ;
        RECT  1.005000  91.860000 15.215000  91.930000 ;
        RECT  1.005000  91.930000 15.145000  92.000000 ;
        RECT  1.005000  92.000000 15.075000  92.070000 ;
        RECT  1.005000  92.070000 15.005000  92.140000 ;
        RECT  1.005000  92.140000 14.935000  92.210000 ;
        RECT  1.005000  92.210000 14.865000  92.280000 ;
        RECT  1.005000  92.280000 14.795000  92.350000 ;
        RECT  1.005000  92.350000 14.725000  92.420000 ;
        RECT  1.005000  92.420000 14.655000  92.490000 ;
        RECT  1.005000  92.490000 14.585000  92.560000 ;
        RECT  1.005000  92.560000 14.515000  92.630000 ;
        RECT  1.005000  92.630000 14.445000  92.700000 ;
        RECT  1.005000  92.700000 14.375000  92.770000 ;
        RECT  1.005000  92.770000 14.305000  92.840000 ;
        RECT  1.005000  92.840000 14.235000  92.910000 ;
        RECT  1.005000  92.910000 14.165000  92.980000 ;
        RECT  1.005000  92.980000 14.120000  93.025000 ;
        RECT  1.005000  93.025000 14.120000 100.240000 ;
        RECT  1.005000 100.240000 14.120000 100.310000 ;
        RECT  1.005000 100.310000 14.190000 100.380000 ;
        RECT  1.005000 100.380000 14.260000 100.450000 ;
        RECT  1.005000 100.450000 14.330000 100.520000 ;
        RECT  1.005000 100.520000 14.400000 100.590000 ;
        RECT  1.005000 100.590000 14.470000 100.660000 ;
        RECT  1.005000 100.660000 14.540000 100.730000 ;
        RECT  1.005000 100.730000 14.610000 100.800000 ;
        RECT  1.005000 100.800000 14.680000 100.870000 ;
        RECT  1.005000 100.870000 14.750000 100.940000 ;
        RECT  1.005000 100.940000 14.820000 101.010000 ;
        RECT  1.005000 101.010000 14.890000 101.080000 ;
        RECT  1.005000 101.080000 14.960000 101.150000 ;
        RECT  1.005000 101.150000 15.030000 101.220000 ;
        RECT  1.005000 101.220000 15.100000 101.290000 ;
        RECT  1.005000 101.290000 15.170000 101.360000 ;
        RECT  1.005000 101.360000 15.240000 101.430000 ;
        RECT  1.005000 101.430000 15.310000 101.500000 ;
        RECT  1.005000 101.500000 15.380000 101.570000 ;
        RECT  1.005000 101.570000 15.450000 101.640000 ;
        RECT  1.005000 101.640000 15.520000 101.710000 ;
        RECT  1.005000 101.710000 15.590000 101.780000 ;
        RECT  1.005000 101.780000 15.660000 101.850000 ;
        RECT  1.005000 101.850000 15.730000 101.920000 ;
        RECT  1.005000 101.920000 15.800000 101.990000 ;
        RECT  1.005000 101.990000 15.870000 102.060000 ;
        RECT  1.005000 102.060000 15.940000 102.130000 ;
        RECT  1.005000 102.130000 16.010000 102.200000 ;
        RECT  1.005000 102.200000 16.080000 102.270000 ;
        RECT  1.005000 102.270000 16.150000 102.340000 ;
        RECT  1.005000 102.340000 16.220000 102.410000 ;
        RECT  1.005000 102.410000 16.290000 102.480000 ;
        RECT  1.005000 102.480000 16.360000 102.550000 ;
        RECT  1.005000 102.550000 16.430000 102.620000 ;
        RECT  1.005000 102.620000 16.500000 102.690000 ;
        RECT  1.005000 102.690000 16.570000 102.760000 ;
        RECT  1.005000 102.760000 16.640000 102.830000 ;
        RECT  1.005000 102.830000 16.710000 102.900000 ;
        RECT  1.005000 102.900000 16.780000 102.970000 ;
        RECT  1.005000 102.970000 16.850000 103.040000 ;
        RECT  1.005000 103.040000 16.920000 103.110000 ;
        RECT  1.005000 103.110000 16.990000 103.180000 ;
        RECT  1.005000 103.180000 17.060000 103.250000 ;
        RECT  1.005000 103.250000 17.130000 103.320000 ;
        RECT  1.005000 103.320000 17.200000 103.390000 ;
        RECT  1.005000 103.390000 17.270000 103.460000 ;
        RECT  1.005000 103.460000 17.340000 103.530000 ;
        RECT  1.005000 103.530000 17.410000 103.600000 ;
        RECT  1.005000 103.600000 17.480000 103.670000 ;
        RECT  1.005000 103.670000 17.550000 103.740000 ;
        RECT  1.005000 103.740000 17.620000 103.780000 ;
        RECT  1.005000 103.780000 56.705000 112.480000 ;
        RECT  1.005000 112.480000 17.635000 112.550000 ;
        RECT  1.005000 112.550000 17.565000 112.620000 ;
        RECT  1.005000 112.620000 17.495000 112.690000 ;
        RECT  1.005000 112.690000 17.425000 112.760000 ;
        RECT  1.005000 112.760000 17.355000 112.830000 ;
        RECT  1.005000 112.830000 17.285000 112.900000 ;
        RECT  1.005000 112.900000 17.215000 112.970000 ;
        RECT  1.005000 112.970000 17.145000 113.040000 ;
        RECT  1.005000 113.040000 17.075000 113.110000 ;
        RECT  1.005000 113.110000 17.005000 113.180000 ;
        RECT  1.005000 113.180000 16.935000 113.250000 ;
        RECT  1.005000 113.250000 16.865000 113.320000 ;
        RECT  1.005000 113.320000 16.795000 113.390000 ;
        RECT  1.005000 113.390000 16.725000 113.460000 ;
        RECT  1.005000 113.460000 16.655000 113.530000 ;
        RECT  1.005000 113.530000 16.585000 113.600000 ;
        RECT  1.005000 113.600000 16.515000 113.670000 ;
        RECT  1.005000 113.670000 16.445000 113.740000 ;
        RECT  1.005000 113.740000 16.375000 113.810000 ;
        RECT  1.005000 113.810000 16.305000 113.880000 ;
        RECT  1.005000 113.880000 16.235000 113.950000 ;
        RECT  1.005000 113.950000 16.165000 114.020000 ;
        RECT  1.005000 114.020000 16.095000 114.090000 ;
        RECT  1.005000 114.090000 16.025000 114.160000 ;
        RECT  1.005000 114.160000 15.955000 114.230000 ;
        RECT  1.005000 114.230000 15.885000 114.300000 ;
        RECT  1.005000 114.300000 15.815000 114.370000 ;
        RECT  1.005000 114.370000 15.745000 114.440000 ;
        RECT  1.005000 114.440000 15.675000 114.510000 ;
        RECT  1.005000 114.510000 15.605000 114.580000 ;
        RECT  1.005000 114.580000 15.535000 114.650000 ;
        RECT  1.005000 114.650000 15.465000 114.720000 ;
        RECT  1.005000 114.720000 15.395000 114.790000 ;
        RECT  1.005000 114.790000 15.325000 114.860000 ;
        RECT  1.005000 114.860000 15.255000 114.930000 ;
        RECT  1.005000 114.930000 15.185000 115.000000 ;
        RECT  1.005000 115.000000 15.115000 115.070000 ;
        RECT  1.005000 115.070000 15.045000 115.140000 ;
        RECT  1.005000 115.140000 14.975000 115.210000 ;
        RECT  1.005000 115.210000 14.905000 115.280000 ;
        RECT  1.005000 115.280000 14.835000 115.350000 ;
        RECT  1.005000 115.350000 14.765000 115.420000 ;
        RECT  1.005000 115.420000 14.695000 115.490000 ;
        RECT  1.005000 115.490000 14.625000 115.560000 ;
        RECT  1.005000 115.560000 14.555000 115.630000 ;
        RECT  1.005000 115.630000 14.485000 115.700000 ;
        RECT  1.005000 115.700000 14.415000 115.770000 ;
        RECT  1.005000 115.770000 14.345000 115.840000 ;
        RECT  1.005000 115.840000 14.275000 115.910000 ;
        RECT  1.005000 115.910000 14.205000 115.980000 ;
        RECT  1.005000 115.980000 14.135000 116.050000 ;
        RECT  1.005000 116.050000 14.120000 116.065000 ;
        RECT  1.005000 116.065000 14.120000 123.145000 ;
        RECT  1.005000 123.145000 14.120000 123.215000 ;
        RECT  1.005000 123.215000 14.190000 123.285000 ;
        RECT  1.005000 123.285000 14.260000 123.355000 ;
        RECT  1.005000 123.355000 14.330000 123.425000 ;
        RECT  1.005000 123.425000 14.400000 123.495000 ;
        RECT  1.005000 123.495000 14.470000 123.565000 ;
        RECT  1.005000 123.565000 14.540000 123.635000 ;
        RECT  1.005000 123.635000 14.610000 123.705000 ;
        RECT  1.005000 123.705000 14.680000 123.775000 ;
        RECT  1.005000 123.775000 14.750000 123.845000 ;
        RECT  1.005000 123.845000 14.820000 123.915000 ;
        RECT  1.005000 123.915000 14.890000 123.985000 ;
        RECT  1.005000 123.985000 14.960000 124.055000 ;
        RECT  1.005000 124.055000 15.030000 124.125000 ;
        RECT  1.005000 124.125000 15.100000 124.195000 ;
        RECT  1.005000 124.195000 15.170000 124.265000 ;
        RECT  1.005000 124.265000 15.240000 124.335000 ;
        RECT  1.005000 124.335000 15.310000 124.405000 ;
        RECT  1.005000 124.405000 15.380000 124.475000 ;
        RECT  1.005000 124.475000 15.450000 124.545000 ;
        RECT  1.005000 124.545000 15.520000 124.615000 ;
        RECT  1.005000 124.615000 15.590000 124.685000 ;
        RECT  1.005000 124.685000 15.660000 124.755000 ;
        RECT  1.005000 124.755000 15.730000 124.825000 ;
        RECT  1.005000 124.825000 15.800000 124.895000 ;
        RECT  1.005000 124.895000 15.870000 124.965000 ;
        RECT  1.005000 124.965000 15.940000 125.035000 ;
        RECT  1.005000 125.035000 16.010000 125.105000 ;
        RECT  1.005000 125.105000 16.080000 125.175000 ;
        RECT  1.005000 125.175000 16.150000 125.245000 ;
        RECT  1.005000 125.245000 16.220000 125.315000 ;
        RECT  1.005000 125.315000 16.290000 125.385000 ;
        RECT  1.005000 125.385000 16.360000 125.455000 ;
        RECT  1.005000 125.455000 16.430000 125.525000 ;
        RECT  1.005000 125.525000 16.500000 125.595000 ;
        RECT  1.005000 125.595000 16.570000 125.665000 ;
        RECT  1.005000 125.665000 16.640000 125.735000 ;
        RECT  1.005000 125.735000 16.710000 125.805000 ;
        RECT  1.005000 125.805000 16.780000 125.875000 ;
        RECT  1.005000 125.875000 16.850000 125.945000 ;
        RECT  1.005000 125.945000 16.920000 126.015000 ;
        RECT  1.005000 126.015000 16.990000 126.085000 ;
        RECT  1.005000 126.085000 17.060000 126.155000 ;
        RECT  1.005000 126.155000 17.130000 126.225000 ;
        RECT  1.005000 126.225000 17.200000 126.295000 ;
        RECT  1.005000 126.295000 17.270000 126.365000 ;
        RECT  1.005000 126.365000 17.340000 126.435000 ;
        RECT  1.005000 126.435000 17.410000 126.505000 ;
        RECT  1.005000 126.505000 17.480000 126.575000 ;
        RECT  1.005000 126.575000 17.550000 126.645000 ;
        RECT  1.005000 126.645000 17.620000 126.715000 ;
        RECT  1.005000 126.715000 17.690000 126.780000 ;
        RECT  1.005000 126.780000 56.705000 135.480000 ;
        RECT  1.005000 135.480000 17.740000 135.550000 ;
        RECT  1.005000 135.550000 17.670000 135.620000 ;
        RECT  1.005000 135.620000 17.600000 135.690000 ;
        RECT  1.005000 135.690000 17.530000 135.760000 ;
        RECT  1.005000 135.760000 17.460000 135.830000 ;
        RECT  1.005000 135.830000 17.390000 135.900000 ;
        RECT  1.005000 135.900000 17.320000 135.970000 ;
        RECT  1.005000 135.970000 17.250000 136.040000 ;
        RECT  1.005000 136.040000 17.180000 136.110000 ;
        RECT  1.005000 136.110000 17.110000 136.180000 ;
        RECT  1.005000 136.180000 17.040000 136.250000 ;
        RECT  1.005000 136.250000 16.970000 136.320000 ;
        RECT  1.005000 136.320000 16.900000 136.390000 ;
        RECT  1.005000 136.390000 16.830000 136.460000 ;
        RECT  1.005000 136.460000 16.760000 136.530000 ;
        RECT  1.005000 136.530000 16.690000 136.600000 ;
        RECT  1.005000 136.600000 16.620000 136.670000 ;
        RECT  1.005000 136.670000 16.550000 136.740000 ;
        RECT  1.005000 136.740000 16.480000 136.810000 ;
        RECT  1.005000 136.810000 16.410000 136.880000 ;
        RECT  1.005000 136.880000 16.340000 136.950000 ;
        RECT  1.005000 136.950000 16.270000 137.020000 ;
        RECT  1.005000 137.020000 16.200000 137.090000 ;
        RECT  1.005000 137.090000 16.130000 137.160000 ;
        RECT  1.005000 137.160000 16.060000 137.230000 ;
        RECT  1.005000 137.230000 15.990000 137.300000 ;
        RECT  1.005000 137.300000 15.920000 137.370000 ;
        RECT  1.005000 137.370000 15.850000 137.440000 ;
        RECT  1.005000 137.440000 15.780000 137.510000 ;
        RECT  1.005000 137.510000 15.710000 137.580000 ;
        RECT  1.005000 137.580000 15.640000 137.650000 ;
        RECT  1.005000 137.650000 15.570000 137.720000 ;
        RECT  1.005000 137.720000 15.500000 137.790000 ;
        RECT  1.005000 137.790000 15.430000 137.860000 ;
        RECT  1.005000 137.860000 15.360000 137.930000 ;
        RECT  1.005000 137.930000 15.290000 138.000000 ;
        RECT  1.005000 138.000000 15.220000 138.070000 ;
        RECT  1.005000 138.070000 15.150000 138.140000 ;
        RECT  1.005000 138.140000 15.080000 138.210000 ;
        RECT  1.005000 138.210000 15.010000 138.280000 ;
        RECT  1.005000 138.280000 14.940000 138.350000 ;
        RECT  1.005000 138.350000 14.870000 138.420000 ;
        RECT  1.005000 138.420000 14.800000 138.490000 ;
        RECT  1.005000 138.490000 14.730000 138.560000 ;
        RECT  1.005000 138.560000 14.660000 138.630000 ;
        RECT  1.005000 138.630000 14.590000 138.700000 ;
        RECT  1.005000 138.700000 14.520000 138.770000 ;
        RECT  1.005000 138.770000 14.450000 138.840000 ;
        RECT  1.005000 138.840000 14.380000 138.910000 ;
        RECT  1.005000 138.910000 14.310000 138.980000 ;
        RECT  1.005000 138.980000 14.240000 139.050000 ;
        RECT  1.005000 139.050000 14.170000 139.120000 ;
        RECT  1.005000 139.120000 14.120000 139.170000 ;
        RECT  1.005000 139.170000 14.120000 146.215000 ;
        RECT  1.005000 146.215000 14.120000 146.285000 ;
        RECT  1.005000 146.285000 14.190000 146.355000 ;
        RECT  1.005000 146.355000 14.260000 146.425000 ;
        RECT  1.005000 146.425000 14.330000 146.495000 ;
        RECT  1.005000 146.495000 14.400000 146.565000 ;
        RECT  1.005000 146.565000 14.470000 146.635000 ;
        RECT  1.005000 146.635000 14.540000 146.705000 ;
        RECT  1.005000 146.705000 14.610000 146.775000 ;
        RECT  1.005000 146.775000 14.680000 146.845000 ;
        RECT  1.005000 146.845000 14.750000 146.915000 ;
        RECT  1.005000 146.915000 14.820000 146.985000 ;
        RECT  1.005000 146.985000 14.890000 147.055000 ;
        RECT  1.005000 147.055000 14.960000 147.125000 ;
        RECT  1.005000 147.125000 15.030000 147.195000 ;
        RECT  1.005000 147.195000 15.100000 147.265000 ;
        RECT  1.005000 147.265000 15.170000 147.335000 ;
        RECT  1.005000 147.335000 15.240000 147.405000 ;
        RECT  1.005000 147.405000 15.310000 147.475000 ;
        RECT  1.005000 147.475000 15.380000 147.545000 ;
        RECT  1.005000 147.545000 15.450000 147.615000 ;
        RECT  1.005000 147.615000 15.520000 147.685000 ;
        RECT  1.005000 147.685000 15.590000 147.755000 ;
        RECT  1.005000 147.755000 15.660000 147.825000 ;
        RECT  1.005000 147.825000 15.730000 147.895000 ;
        RECT  1.005000 147.895000 15.800000 147.965000 ;
        RECT  1.005000 147.965000 15.870000 148.035000 ;
        RECT  1.005000 148.035000 15.940000 148.105000 ;
        RECT  1.005000 148.105000 16.010000 148.175000 ;
        RECT  1.005000 148.175000 16.080000 148.245000 ;
        RECT  1.005000 148.245000 16.150000 148.315000 ;
        RECT  1.005000 148.315000 16.220000 148.385000 ;
        RECT  1.005000 148.385000 16.290000 148.455000 ;
        RECT  1.005000 148.455000 16.360000 148.525000 ;
        RECT  1.005000 148.525000 16.430000 148.595000 ;
        RECT  1.005000 148.595000 16.500000 148.665000 ;
        RECT  1.005000 148.665000 16.570000 148.735000 ;
        RECT  1.005000 148.735000 16.640000 148.805000 ;
        RECT  1.005000 148.805000 16.710000 148.875000 ;
        RECT  1.005000 148.875000 16.780000 148.945000 ;
        RECT  1.005000 148.945000 16.850000 149.015000 ;
        RECT  1.005000 149.015000 16.920000 149.085000 ;
        RECT  1.005000 149.085000 16.990000 149.155000 ;
        RECT  1.005000 149.155000 17.060000 149.225000 ;
        RECT  1.005000 149.225000 17.130000 149.295000 ;
        RECT  1.005000 149.295000 17.200000 149.365000 ;
        RECT  1.005000 149.365000 17.270000 149.435000 ;
        RECT  1.005000 149.435000 17.340000 149.505000 ;
        RECT  1.005000 149.505000 17.410000 149.575000 ;
        RECT  1.005000 149.575000 17.480000 149.645000 ;
        RECT  1.005000 149.645000 17.550000 149.715000 ;
        RECT  1.005000 149.715000 17.620000 149.780000 ;
        RECT  1.005000 149.780000 56.705000 158.480000 ;
        RECT  1.005000 158.480000 17.650000 158.550000 ;
        RECT  1.005000 158.550000 17.580000 158.620000 ;
        RECT  1.005000 158.620000 17.510000 158.690000 ;
        RECT  1.005000 158.690000 17.440000 158.760000 ;
        RECT  1.005000 158.760000 17.370000 158.830000 ;
        RECT  1.005000 158.830000 17.300000 158.900000 ;
        RECT  1.005000 158.900000 17.230000 158.970000 ;
        RECT  1.005000 158.970000 17.160000 159.040000 ;
        RECT  1.005000 159.040000 17.090000 159.110000 ;
        RECT  1.005000 159.110000 17.020000 159.180000 ;
        RECT  1.005000 159.180000 16.950000 159.250000 ;
        RECT  1.005000 159.250000 16.880000 159.320000 ;
        RECT  1.005000 159.320000 16.810000 159.390000 ;
        RECT  1.005000 159.390000 16.740000 159.460000 ;
        RECT  1.005000 159.460000 16.670000 159.530000 ;
        RECT  1.005000 159.530000 16.600000 159.600000 ;
        RECT  1.005000 159.600000 16.530000 159.670000 ;
        RECT  1.005000 159.670000 16.460000 159.740000 ;
        RECT  1.005000 159.740000 16.390000 159.810000 ;
        RECT  1.005000 159.810000 16.320000 159.880000 ;
        RECT  1.005000 159.880000 16.250000 159.950000 ;
        RECT  1.005000 159.950000 16.180000 160.020000 ;
        RECT  1.005000 160.020000 16.110000 160.090000 ;
        RECT  1.005000 160.090000 16.040000 160.160000 ;
        RECT  1.005000 160.160000 15.970000 160.230000 ;
        RECT  1.005000 160.230000 15.900000 160.300000 ;
        RECT  1.005000 160.300000 15.830000 160.370000 ;
        RECT  1.005000 160.370000 15.760000 160.440000 ;
        RECT  1.005000 160.440000 15.690000 160.510000 ;
        RECT  1.005000 160.510000 15.620000 160.580000 ;
        RECT  1.005000 160.580000 15.550000 160.650000 ;
        RECT  1.005000 160.650000 15.480000 160.720000 ;
        RECT  1.005000 160.720000 15.410000 160.790000 ;
        RECT  1.005000 160.790000 15.340000 160.860000 ;
        RECT  1.005000 160.860000 15.270000 160.930000 ;
        RECT  1.005000 160.930000 15.200000 161.000000 ;
        RECT  1.005000 161.000000 15.130000 161.070000 ;
        RECT  1.005000 161.070000 15.060000 161.140000 ;
        RECT  1.005000 161.140000 14.990000 161.210000 ;
        RECT  1.005000 161.210000 14.920000 161.280000 ;
        RECT  1.005000 161.280000 14.850000 161.350000 ;
        RECT  1.005000 161.350000 14.780000 161.420000 ;
        RECT  1.005000 161.420000 14.710000 161.490000 ;
        RECT  1.005000 161.490000 14.640000 161.560000 ;
        RECT  1.005000 161.560000 14.570000 161.630000 ;
        RECT  1.005000 161.630000 14.500000 161.700000 ;
        RECT  1.005000 161.700000 14.430000 161.770000 ;
        RECT  1.005000 161.770000 14.360000 161.840000 ;
        RECT  1.005000 161.840000 14.290000 161.910000 ;
        RECT  1.005000 161.910000 14.220000 161.980000 ;
        RECT  1.005000 161.980000 14.150000 162.050000 ;
        RECT  1.005000 162.050000 14.120000 162.080000 ;
        RECT  1.005000 162.080000 14.120000 169.220000 ;
        RECT  1.005000 169.220000 14.120000 169.290000 ;
        RECT  1.005000 169.290000 14.190000 169.360000 ;
        RECT  1.005000 169.360000 14.260000 169.430000 ;
        RECT  1.005000 169.430000 14.330000 169.500000 ;
        RECT  1.005000 169.500000 14.400000 169.570000 ;
        RECT  1.005000 169.570000 14.470000 169.640000 ;
        RECT  1.005000 169.640000 14.540000 169.710000 ;
        RECT  1.005000 169.710000 14.610000 169.780000 ;
        RECT  1.005000 169.780000 14.680000 169.850000 ;
        RECT  1.005000 169.850000 14.750000 169.920000 ;
        RECT  1.005000 169.920000 14.820000 169.990000 ;
        RECT  1.005000 169.990000 14.890000 170.060000 ;
        RECT  1.005000 170.060000 14.960000 170.130000 ;
        RECT  1.005000 170.130000 15.030000 170.200000 ;
        RECT  1.005000 170.200000 15.100000 170.270000 ;
        RECT  1.005000 170.270000 15.170000 170.340000 ;
        RECT  1.005000 170.340000 15.240000 170.410000 ;
        RECT  1.005000 170.410000 15.310000 170.480000 ;
        RECT  1.005000 170.480000 15.380000 170.550000 ;
        RECT  1.005000 170.550000 15.450000 170.620000 ;
        RECT  1.005000 170.620000 15.520000 170.690000 ;
        RECT  1.005000 170.690000 15.590000 170.760000 ;
        RECT  1.005000 170.760000 15.660000 170.830000 ;
        RECT  1.005000 170.830000 15.730000 170.900000 ;
        RECT  1.005000 170.900000 15.800000 170.970000 ;
        RECT  1.005000 170.970000 15.870000 171.040000 ;
        RECT  1.005000 171.040000 15.940000 171.110000 ;
        RECT  1.005000 171.110000 16.010000 171.180000 ;
        RECT  1.005000 171.180000 16.080000 171.250000 ;
        RECT  1.005000 171.250000 16.150000 171.320000 ;
        RECT  1.005000 171.320000 16.220000 171.390000 ;
        RECT  1.005000 171.390000 16.290000 171.460000 ;
        RECT  1.005000 171.460000 16.360000 171.530000 ;
        RECT  1.005000 171.530000 16.430000 171.600000 ;
        RECT  1.005000 171.600000 16.500000 171.670000 ;
        RECT  1.005000 171.670000 16.570000 171.740000 ;
        RECT  1.005000 171.740000 16.640000 171.810000 ;
        RECT  1.005000 171.810000 16.710000 171.880000 ;
        RECT  1.005000 171.880000 16.780000 171.950000 ;
        RECT  1.005000 171.950000 16.850000 172.020000 ;
        RECT  1.005000 172.020000 16.920000 172.090000 ;
        RECT  1.005000 172.090000 16.990000 172.160000 ;
        RECT  1.005000 172.160000 17.060000 172.230000 ;
        RECT  1.005000 172.230000 17.130000 172.300000 ;
        RECT  1.005000 172.300000 17.200000 172.370000 ;
        RECT  1.005000 172.370000 17.270000 172.440000 ;
        RECT  1.005000 172.440000 17.340000 172.510000 ;
        RECT  1.005000 172.510000 17.410000 172.580000 ;
        RECT  1.005000 172.580000 17.480000 172.650000 ;
        RECT  1.005000 172.650000 17.550000 172.720000 ;
        RECT  1.005000 172.720000 17.620000 172.780000 ;
        RECT  1.005000 172.780000 57.960000 181.480000 ;
        RECT  1.005000 181.480000 17.625000 181.550000 ;
        RECT  1.005000 181.550000 17.555000 181.620000 ;
        RECT  1.005000 181.620000 17.485000 181.690000 ;
        RECT  1.005000 181.690000 17.415000 181.760000 ;
        RECT  1.005000 181.760000 17.345000 181.830000 ;
        RECT  1.005000 181.830000 17.275000 181.900000 ;
        RECT  1.005000 181.900000 17.205000 181.970000 ;
        RECT  1.005000 181.970000 17.135000 182.040000 ;
        RECT  1.005000 182.040000 17.065000 182.110000 ;
        RECT  1.005000 182.110000 16.995000 182.180000 ;
        RECT  1.005000 182.180000 16.925000 182.250000 ;
        RECT  1.005000 182.250000 16.855000 182.320000 ;
        RECT  1.005000 182.320000 16.785000 182.390000 ;
        RECT  1.005000 182.390000 16.715000 182.460000 ;
        RECT  1.005000 182.460000 16.645000 182.530000 ;
        RECT  1.005000 182.530000 16.575000 182.600000 ;
        RECT  1.005000 182.600000 16.505000 182.670000 ;
        RECT  1.005000 182.670000 16.435000 182.740000 ;
        RECT  1.005000 182.740000 16.365000 182.810000 ;
        RECT  1.005000 182.810000 16.295000 182.880000 ;
        RECT  1.005000 182.880000 16.225000 182.950000 ;
        RECT  1.005000 182.950000 16.155000 183.020000 ;
        RECT  1.005000 183.020000 16.085000 183.090000 ;
        RECT  1.005000 183.090000 16.015000 183.160000 ;
        RECT  1.005000 183.160000 15.945000 183.230000 ;
        RECT  1.005000 183.230000 15.875000 183.300000 ;
        RECT  1.005000 183.300000 15.805000 183.370000 ;
        RECT  1.005000 183.370000 15.735000 183.440000 ;
        RECT  1.005000 183.440000 15.665000 183.510000 ;
        RECT  1.005000 183.510000 15.595000 183.580000 ;
        RECT  1.005000 183.580000 15.525000 183.650000 ;
        RECT  1.005000 183.650000 15.455000 183.720000 ;
        RECT  1.005000 183.720000 15.385000 183.790000 ;
        RECT  1.005000 183.790000 15.315000 183.860000 ;
        RECT  1.005000 183.860000 15.245000 183.930000 ;
        RECT  1.005000 183.930000 15.175000 184.000000 ;
        RECT  1.005000 184.000000 15.105000 184.070000 ;
        RECT  1.005000 184.070000 15.035000 184.140000 ;
        RECT  1.005000 184.140000 14.965000 184.210000 ;
        RECT  1.005000 184.210000 14.895000 184.280000 ;
        RECT  1.005000 184.280000 14.825000 184.350000 ;
        RECT  1.005000 184.350000 14.755000 184.420000 ;
        RECT  1.005000 184.420000 14.685000 184.490000 ;
        RECT  1.005000 184.490000 14.615000 184.560000 ;
        RECT  1.005000 184.560000 14.545000 184.630000 ;
        RECT  1.005000 184.630000 14.475000 184.700000 ;
        RECT  1.005000 184.700000 14.405000 184.770000 ;
        RECT  1.005000 184.770000 14.335000 184.840000 ;
        RECT  1.005000 184.840000 14.265000 184.910000 ;
        RECT  1.005000 184.910000 14.195000 184.980000 ;
        RECT  1.005000 184.980000 14.125000 185.050000 ;
        RECT  1.005000 185.050000 14.120000 185.055000 ;
        RECT  1.005000 185.055000 14.120000 189.585000 ;
        RECT  1.005000 189.585000 14.120000 189.655000 ;
        RECT  1.005000 189.655000 14.190000 189.725000 ;
        RECT  1.005000 189.725000 14.260000 189.795000 ;
        RECT  1.005000 189.795000 14.330000 189.865000 ;
        RECT  1.005000 189.865000 14.400000 189.935000 ;
        RECT  1.005000 189.935000 14.470000 190.005000 ;
        RECT  1.005000 190.005000 14.540000 190.075000 ;
        RECT  1.005000 190.075000 14.610000 190.145000 ;
        RECT  1.005000 190.145000 14.680000 190.215000 ;
        RECT  1.005000 190.215000 14.750000 190.285000 ;
        RECT  1.005000 190.285000 14.820000 190.355000 ;
        RECT  1.005000 190.355000 14.890000 190.425000 ;
        RECT  1.005000 190.425000 14.960000 190.495000 ;
        RECT  1.005000 190.495000 15.030000 190.560000 ;
        RECT  1.005000 190.560000 67.200000 195.075000 ;
        RECT  1.010000  47.095000 14.120000  47.100000 ;
        RECT  1.045000  36.855000 16.395000  36.895000 ;
        RECT  1.050000  47.055000 14.120000  47.095000 ;
        RECT  1.085000  36.895000 16.435000  36.935000 ;
        RECT  1.090000  36.935000 16.475000  36.940000 ;
        RECT  1.090000  36.940000 16.480000  37.010000 ;
        RECT  1.090000  37.010000 16.550000  37.080000 ;
        RECT  1.090000  37.080000 16.620000  37.150000 ;
        RECT  1.090000  37.150000 16.690000  37.220000 ;
        RECT  1.090000  37.220000 16.760000  37.290000 ;
        RECT  1.090000  37.290000 16.830000  37.360000 ;
        RECT  1.090000  37.360000 16.900000  37.430000 ;
        RECT  1.090000  37.430000 16.970000  37.500000 ;
        RECT  1.090000  37.500000 17.040000  37.570000 ;
        RECT  1.090000  37.570000 17.110000  37.640000 ;
        RECT  1.090000  37.640000 17.180000  37.710000 ;
        RECT  1.090000  37.710000 17.250000  37.780000 ;
        RECT  1.090000  37.780000 17.320000  37.850000 ;
        RECT  1.090000  37.850000 17.390000  37.920000 ;
        RECT  1.090000  37.920000 17.460000  37.990000 ;
        RECT  1.090000  37.990000 17.530000  38.060000 ;
        RECT  1.090000  38.060000 17.600000  38.130000 ;
        RECT  1.090000  38.130000 17.670000  38.200000 ;
        RECT  1.090000  38.200000 17.740000  38.270000 ;
        RECT  1.090000  38.270000 17.810000  38.340000 ;
        RECT  1.090000  38.340000 17.880000  38.410000 ;
        RECT  1.090000  38.410000 17.950000  38.480000 ;
        RECT  1.090000  38.480000 18.020000  38.550000 ;
        RECT  1.090000  38.550000 18.090000  38.620000 ;
        RECT  1.090000  38.620000 18.160000  38.690000 ;
        RECT  1.090000  38.690000 18.230000  38.760000 ;
        RECT  1.090000  38.760000 18.300000  38.830000 ;
        RECT  1.090000  38.830000 18.370000  38.900000 ;
        RECT  1.090000  38.900000 18.440000  38.970000 ;
        RECT  1.090000  38.970000 18.510000  39.040000 ;
        RECT  1.090000  39.040000 18.580000  39.110000 ;
        RECT  1.090000  39.110000 18.650000  39.180000 ;
        RECT  1.090000  39.180000 18.720000  39.250000 ;
        RECT  1.090000  39.250000 18.790000  39.320000 ;
        RECT  1.090000  39.320000 18.860000  39.390000 ;
        RECT  1.090000  39.390000 18.930000  39.460000 ;
        RECT  1.090000  39.460000 19.000000  39.530000 ;
        RECT  1.090000  39.530000 19.070000  39.600000 ;
        RECT  1.090000  39.600000 19.140000  39.670000 ;
        RECT  1.090000  39.670000 19.210000  39.740000 ;
        RECT  1.090000  39.740000 19.280000  39.810000 ;
        RECT  1.090000  39.810000 19.350000  39.880000 ;
        RECT  1.090000  39.880000 19.420000  39.950000 ;
        RECT  1.090000  39.950000 19.490000  40.020000 ;
        RECT  1.090000  40.020000 19.560000  40.090000 ;
        RECT  1.090000  40.090000 19.630000  40.160000 ;
        RECT  1.090000  40.160000 19.700000  40.230000 ;
        RECT  1.090000  40.230000 19.770000  40.300000 ;
        RECT  1.090000  40.300000 19.840000  40.350000 ;
        RECT  1.090000  40.350000 56.160000  40.420000 ;
        RECT  1.090000  40.420000 56.090000  40.490000 ;
        RECT  1.090000  40.490000 56.020000  40.560000 ;
        RECT  1.090000  40.560000 55.950000  40.630000 ;
        RECT  1.090000  40.630000 55.880000  40.700000 ;
        RECT  1.090000  40.700000 55.810000  40.770000 ;
        RECT  1.090000  40.770000 55.740000  40.840000 ;
        RECT  1.090000  40.840000 55.670000  40.910000 ;
        RECT  1.090000  40.910000 55.600000  40.980000 ;
        RECT  1.090000  40.980000 55.530000  41.050000 ;
        RECT  1.090000  41.050000 55.460000  41.120000 ;
        RECT  1.090000  41.120000 55.390000  41.190000 ;
        RECT  1.090000  41.190000 55.320000  41.260000 ;
        RECT  1.090000  41.260000 55.250000  41.330000 ;
        RECT  1.090000  41.330000 55.180000  41.400000 ;
        RECT  1.090000  41.400000 55.110000  41.470000 ;
        RECT  1.090000  41.470000 55.040000  41.540000 ;
        RECT  1.090000  41.540000 54.970000  41.610000 ;
        RECT  1.090000  41.610000 54.900000  41.680000 ;
        RECT  1.090000  41.680000 54.830000  41.750000 ;
        RECT  1.090000  41.750000 54.760000  41.820000 ;
        RECT  1.090000  41.820000 54.690000  41.890000 ;
        RECT  1.090000  41.890000 54.620000  41.960000 ;
        RECT  1.090000  41.960000 54.550000  42.030000 ;
        RECT  1.090000  42.030000 54.480000  42.100000 ;
        RECT  1.090000  42.100000 54.410000  42.170000 ;
        RECT  1.090000  42.170000 54.340000  42.240000 ;
        RECT  1.090000  42.240000 54.270000  42.310000 ;
        RECT  1.090000  42.310000 54.200000  42.380000 ;
        RECT  1.090000  42.380000 16.985000  42.450000 ;
        RECT  1.090000  42.450000 16.915000  42.520000 ;
        RECT  1.090000  42.520000 16.845000  42.590000 ;
        RECT  1.090000  42.590000 16.775000  42.660000 ;
        RECT  1.090000  42.660000 16.705000  42.730000 ;
        RECT  1.090000  42.730000 16.635000  42.800000 ;
        RECT  1.090000  42.800000 16.565000  42.870000 ;
        RECT  1.090000  42.870000 16.495000  42.940000 ;
        RECT  1.090000  42.940000 16.425000  43.010000 ;
        RECT  1.090000  43.010000 16.355000  43.080000 ;
        RECT  1.090000  43.080000 16.285000  43.150000 ;
        RECT  1.090000  43.150000 16.215000  43.220000 ;
        RECT  1.090000  43.220000 16.145000  43.290000 ;
        RECT  1.090000  43.290000 16.075000  43.360000 ;
        RECT  1.090000  43.360000 16.005000  43.430000 ;
        RECT  1.090000  43.430000 15.935000  43.500000 ;
        RECT  1.090000  43.500000 15.865000  43.570000 ;
        RECT  1.090000  43.570000 15.795000  43.640000 ;
        RECT  1.090000  43.640000 15.725000  43.710000 ;
        RECT  1.090000  43.710000 15.655000  43.780000 ;
        RECT  1.090000  43.780000 15.585000  43.850000 ;
        RECT  1.090000  43.850000 15.515000  43.920000 ;
        RECT  1.090000  43.920000 15.445000  43.990000 ;
        RECT  1.090000  43.990000 15.375000  44.060000 ;
        RECT  1.090000  44.060000 15.305000  44.130000 ;
        RECT  1.090000  44.130000 15.235000  44.200000 ;
        RECT  1.090000  44.200000 15.165000  44.270000 ;
        RECT  1.090000  44.270000 15.095000  44.340000 ;
        RECT  1.090000  44.340000 15.025000  44.410000 ;
        RECT  1.090000  44.410000 14.955000  44.480000 ;
        RECT  1.090000  44.480000 14.885000  44.550000 ;
        RECT  1.090000  44.550000 14.815000  44.620000 ;
        RECT  1.090000  44.620000 14.745000  44.690000 ;
        RECT  1.090000  44.690000 14.675000  44.760000 ;
        RECT  1.090000  44.760000 14.605000  44.830000 ;
        RECT  1.090000  44.830000 14.535000  44.900000 ;
        RECT  1.090000  44.900000 14.465000  44.970000 ;
        RECT  1.090000  44.970000 14.395000  45.040000 ;
        RECT  1.090000  45.040000 14.325000  45.110000 ;
        RECT  1.090000  45.110000 14.255000  45.180000 ;
        RECT  1.090000  45.180000 14.185000  45.250000 ;
        RECT  1.090000  45.250000 14.120000  45.315000 ;
        RECT  1.090000  45.315000 14.120000  47.015000 ;
        RECT  1.090000  47.015000 14.120000  47.055000 ;
        RECT 52.630000  40.295000 56.230000  40.350000 ;
        RECT 52.700000  40.225000 56.285000  40.295000 ;
        RECT 52.770000  40.155000 56.355000  40.225000 ;
        RECT 52.840000  40.085000 56.425000  40.155000 ;
        RECT 52.910000  40.015000 56.495000  40.085000 ;
        RECT 52.980000  39.945000 56.565000  40.015000 ;
        RECT 53.050000  39.875000 56.635000  39.945000 ;
        RECT 53.120000  39.805000 56.705000  39.875000 ;
        RECT 53.190000  39.735000 56.775000  39.805000 ;
        RECT 53.260000  39.665000 56.845000  39.735000 ;
        RECT 53.270000  39.655000 56.915000  39.665000 ;
        RECT 53.340000  39.585000 56.915000  39.655000 ;
        RECT 53.410000  39.515000 56.915000  39.585000 ;
        RECT 53.480000  39.445000 56.915000  39.515000 ;
        RECT 53.550000  39.375000 56.915000  39.445000 ;
        RECT 53.620000  39.305000 56.915000  39.375000 ;
        RECT 53.690000  39.235000 56.915000  39.305000 ;
        RECT 53.760000  39.165000 56.915000  39.235000 ;
        RECT 53.830000  39.095000 56.915000  39.165000 ;
        RECT 53.900000  39.025000 56.915000  39.095000 ;
        RECT 53.970000  38.955000 56.915000  39.025000 ;
        RECT 54.040000  38.885000 56.915000  38.955000 ;
        RECT 54.110000  38.815000 56.915000  38.885000 ;
        RECT 54.180000  38.745000 56.915000  38.815000 ;
        RECT 54.250000  38.675000 56.915000  38.745000 ;
        RECT 54.320000  38.605000 56.915000  38.675000 ;
        RECT 54.390000  38.535000 56.915000  38.605000 ;
        RECT 54.460000  38.465000 56.915000  38.535000 ;
        RECT 54.530000  38.395000 56.915000  38.465000 ;
        RECT 54.600000  38.325000 56.915000  38.395000 ;
        RECT 54.670000  36.115000 56.915000  38.255000 ;
        RECT 54.670000  38.255000 56.915000  38.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT  3.160000 185.360000 25.010000 200.000000 ;
        RECT  3.200000 185.320000 25.010000 185.360000 ;
        RECT  3.350000 185.170000 25.010000 185.320000 ;
        RECT  3.500000 185.020000 25.010000 185.170000 ;
        RECT  3.650000 184.870000 25.010000 185.020000 ;
        RECT  3.800000 184.720000 25.010000 184.870000 ;
        RECT  3.950000 184.570000 25.010000 184.720000 ;
        RECT  4.100000 184.420000 25.010000 184.570000 ;
        RECT  4.250000 184.270000 25.010000 184.420000 ;
        RECT  4.400000 184.120000 25.010000 184.270000 ;
        RECT  4.550000 183.970000 25.010000 184.120000 ;
        RECT  4.700000 183.820000 25.010000 183.970000 ;
        RECT  4.850000 183.670000 25.010000 183.820000 ;
        RECT  5.000000 183.520000 25.010000 183.670000 ;
        RECT  5.150000 183.370000 25.010000 183.520000 ;
        RECT  5.300000 183.220000 25.010000 183.370000 ;
        RECT  5.450000 183.070000 25.010000 183.220000 ;
        RECT  5.600000 182.920000 25.010000 183.070000 ;
        RECT  5.750000 182.770000 25.010000 182.920000 ;
        RECT  5.900000 182.620000 25.010000 182.770000 ;
        RECT  6.050000 182.470000 25.010000 182.620000 ;
        RECT  6.200000 182.320000 25.010000 182.470000 ;
        RECT  6.350000 182.170000 25.010000 182.320000 ;
        RECT  6.500000 182.020000 25.010000 182.170000 ;
        RECT  6.650000 181.870000 25.010000 182.020000 ;
        RECT  6.800000 181.720000 25.010000 181.870000 ;
        RECT  6.950000 181.570000 25.010000 181.720000 ;
        RECT  7.100000 181.420000 25.010000 181.570000 ;
        RECT  7.250000 181.270000 25.010000 181.420000 ;
        RECT  7.400000 181.120000 25.010000 181.270000 ;
        RECT  7.550000 180.970000 25.010000 181.120000 ;
        RECT  7.700000 180.820000 25.010000 180.970000 ;
        RECT  7.850000 180.670000 25.010000 180.820000 ;
        RECT  8.000000 180.520000 25.010000 180.670000 ;
        RECT  8.150000 180.370000 25.010000 180.520000 ;
        RECT  8.300000 180.220000 25.010000 180.370000 ;
        RECT  8.450000 180.070000 25.010000 180.220000 ;
        RECT  8.600000 179.920000 25.010000 180.070000 ;
        RECT  8.750000 179.770000 25.010000 179.920000 ;
        RECT  8.900000 179.620000 25.010000 179.770000 ;
        RECT  9.050000 179.470000 25.010000 179.620000 ;
        RECT  9.200000 179.320000 25.010000 179.470000 ;
        RECT  9.350000 179.170000 25.010000 179.320000 ;
        RECT  9.500000 179.020000 25.010000 179.170000 ;
        RECT  9.650000 178.870000 25.010000 179.020000 ;
        RECT  9.800000 178.720000 25.010000 178.870000 ;
        RECT  9.950000 178.570000 25.010000 178.720000 ;
        RECT 10.100000 178.420000 25.010000 178.570000 ;
        RECT 10.250000 178.270000 25.010000 178.420000 ;
        RECT 10.400000 178.120000 25.010000 178.270000 ;
        RECT 10.550000 177.970000 25.010000 178.120000 ;
        RECT 10.700000 177.820000 25.010000 177.970000 ;
        RECT 10.850000 177.670000 25.010000 177.820000 ;
        RECT 11.000000 177.520000 25.010000 177.670000 ;
        RECT 11.150000 177.370000 25.010000 177.520000 ;
        RECT 11.300000 177.220000 25.010000 177.370000 ;
        RECT 11.450000 177.070000 25.010000 177.220000 ;
        RECT 11.600000 176.920000 25.010000 177.070000 ;
        RECT 11.750000 176.770000 25.010000 176.920000 ;
        RECT 11.900000 176.620000 25.010000 176.770000 ;
        RECT 12.050000 176.470000 25.010000 176.620000 ;
        RECT 12.200000 176.320000 25.010000 176.470000 ;
        RECT 12.350000 176.170000 25.010000 176.320000 ;
        RECT 12.500000 176.020000 25.010000 176.170000 ;
        RECT 12.650000 175.870000 25.010000 176.020000 ;
        RECT 12.800000 175.720000 25.010000 175.870000 ;
        RECT 12.950000 175.570000 25.010000 175.720000 ;
        RECT 13.100000 175.420000 25.010000 175.570000 ;
        RECT 13.250000 175.270000 25.010000 175.420000 ;
        RECT 13.400000 175.120000 25.010000 175.270000 ;
        RECT 13.550000 174.970000 25.010000 175.120000 ;
        RECT 13.700000 174.820000 25.010000 174.970000 ;
        RECT 13.850000 174.670000 25.010000 174.820000 ;
        RECT 14.000000 174.520000 25.010000 174.670000 ;
        RECT 14.150000 174.370000 25.010000 174.520000 ;
        RECT 14.300000 174.220000 25.010000 174.370000 ;
        RECT 14.450000 174.070000 25.010000 174.220000 ;
        RECT 14.600000 173.920000 25.010000 174.070000 ;
        RECT 14.750000 173.770000 25.010000 173.920000 ;
        RECT 14.900000 173.620000 25.010000 173.770000 ;
        RECT 15.050000 173.470000 25.010000 173.620000 ;
        RECT 15.200000 173.320000 25.010000 173.470000 ;
        RECT 15.350000 173.170000 25.010000 173.320000 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
        RECT 15.500000 169.130000 21.500000 169.280000 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
        RECT 15.500000 171.230000 23.600000 171.380000 ;
        RECT 15.500000 171.380000 23.750000 171.530000 ;
        RECT 15.500000 171.530000 23.900000 171.680000 ;
        RECT 15.500000 171.680000 24.050000 171.830000 ;
        RECT 15.500000 171.830000 24.200000 171.980000 ;
        RECT 15.500000 171.980000 24.350000 172.130000 ;
        RECT 15.500000 172.130000 24.500000 172.280000 ;
        RECT 15.500000 172.280000 24.650000 172.430000 ;
        RECT 15.500000 172.430000 24.800000 172.580000 ;
        RECT 15.500000 172.580000 24.950000 172.640000 ;
        RECT 15.500000 172.640000 25.010000 173.020000 ;
        RECT 15.500000 173.020000 25.010000 173.170000 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
        RECT 17.595000 100.105000 25.925000 100.255000 ;
        RECT 17.745000  99.955000 26.075000 100.105000 ;
        RECT 17.895000  99.805000 26.225000  99.955000 ;
        RECT 18.045000  99.655000 26.375000  99.805000 ;
        RECT 18.195000  99.505000 26.525000  99.655000 ;
        RECT 18.345000  99.355000 26.675000  99.505000 ;
        RECT 18.495000  99.205000 26.825000  99.355000 ;
        RECT 18.645000  99.055000 26.975000  99.205000 ;
        RECT 18.795000  98.905000 27.125000  99.055000 ;
        RECT 18.945000  98.755000 27.275000  98.905000 ;
        RECT 19.095000  98.605000 27.425000  98.755000 ;
        RECT 19.245000  98.455000 27.575000  98.605000 ;
        RECT 19.395000  98.305000 27.725000  98.455000 ;
        RECT 19.545000  98.155000 27.875000  98.305000 ;
        RECT 19.695000  98.005000 28.025000  98.155000 ;
        RECT 19.845000  97.855000 28.175000  98.005000 ;
        RECT 19.995000  97.705000 28.325000  97.855000 ;
        RECT 20.145000  97.555000 28.475000  97.705000 ;
        RECT 20.295000  97.405000 28.625000  97.555000 ;
        RECT 20.445000  97.255000 28.775000  97.405000 ;
        RECT 20.595000  97.105000 28.925000  97.255000 ;
        RECT 20.745000  96.955000 29.075000  97.105000 ;
        RECT 20.895000  96.805000 29.225000  96.955000 ;
        RECT 21.045000  96.655000 29.375000  96.805000 ;
        RECT 21.195000  96.505000 29.525000  96.655000 ;
        RECT 21.345000  96.355000 29.525000  96.505000 ;
        RECT 21.495000  96.205000 29.525000  96.355000 ;
        RECT 21.645000  96.055000 29.525000  96.205000 ;
        RECT 21.795000  95.905000 29.525000  96.055000 ;
        RECT 21.945000  95.755000 29.525000  95.905000 ;
        RECT 22.095000  95.605000 29.525000  95.755000 ;
        RECT 22.245000  95.455000 29.525000  95.605000 ;
        RECT 22.395000  95.305000 29.525000  95.455000 ;
        RECT 22.545000  95.155000 29.525000  95.305000 ;
        RECT 22.695000  95.005000 29.525000  95.155000 ;
        RECT 22.845000  94.855000 29.525000  95.005000 ;
        RECT 22.995000  94.705000 29.525000  94.855000 ;
        RECT 23.145000  94.555000 29.525000  94.705000 ;
        RECT 23.295000  94.405000 29.525000  94.555000 ;
        RECT 23.445000  94.255000 29.525000  94.405000 ;
        RECT 23.595000  94.105000 29.525000  94.255000 ;
        RECT 23.745000  92.540000 29.935000  92.690000 ;
        RECT 23.745000  92.690000 29.785000  92.840000 ;
        RECT 23.745000  92.840000 29.635000  92.990000 ;
        RECT 23.745000  92.990000 29.525000  93.100000 ;
        RECT 23.745000  93.100000 29.525000  93.955000 ;
        RECT 23.745000  93.955000 29.525000  94.105000 ;
        RECT 23.820000  92.465000 30.085000  92.540000 ;
        RECT 23.895000  92.390000 30.160000  92.465000 ;
        RECT 23.945000  92.340000 36.895000  92.390000 ;
        RECT 24.095000  92.190000 36.895000  92.340000 ;
        RECT 24.245000  92.040000 36.895000  92.190000 ;
        RECT 24.395000  91.890000 36.895000  92.040000 ;
        RECT 24.545000  91.740000 36.895000  91.890000 ;
        RECT 24.695000  91.590000 36.895000  91.740000 ;
        RECT 24.845000  91.440000 36.895000  91.590000 ;
        RECT 24.995000  91.290000 36.895000  91.440000 ;
        RECT 25.145000  91.140000 36.895000  91.290000 ;
        RECT 25.295000  90.990000 36.895000  91.140000 ;
        RECT 25.445000  90.840000 36.895000  90.990000 ;
        RECT 25.595000  90.690000 36.895000  90.840000 ;
        RECT 25.745000  90.540000 36.895000  90.690000 ;
        RECT 25.895000   0.000000 36.895000  90.390000 ;
        RECT 25.895000  90.390000 36.895000  90.540000 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
        RECT 25.930000 170.460000 31.930000 170.610000 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
        RECT 25.930000 172.710000 34.180000 172.860000 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
        RECT 25.930000 173.310000 34.780000 173.460000 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
        RECT 25.930000 174.060000 35.530000 174.210000 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
        RECT 25.930000 174.660000 36.130000 174.810000 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
        RECT 25.930000 175.260000 36.730000 175.350000 ;
        RECT 25.930000 175.350000 36.820000 200.000000 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
        RECT 27.975000 100.345000 36.295000 100.495000 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
        RECT 28.425000  99.895000 36.745000 100.045000 ;
        RECT 28.495000  99.825000 36.895000  99.895000 ;
        RECT 28.645000  99.675000 36.895000  99.825000 ;
        RECT 28.795000  99.525000 36.895000  99.675000 ;
        RECT 28.945000  99.375000 36.895000  99.525000 ;
        RECT 29.095000  99.225000 36.895000  99.375000 ;
        RECT 29.245000  99.075000 36.895000  99.225000 ;
        RECT 29.395000  98.925000 36.895000  99.075000 ;
        RECT 29.545000  98.775000 36.895000  98.925000 ;
        RECT 29.695000  98.625000 36.895000  98.775000 ;
        RECT 29.845000  98.475000 36.895000  98.625000 ;
        RECT 29.995000  98.325000 36.895000  98.475000 ;
        RECT 30.145000  98.175000 36.895000  98.325000 ;
        RECT 30.295000  98.025000 36.895000  98.175000 ;
        RECT 30.445000  97.875000 36.895000  98.025000 ;
        RECT 30.595000  97.725000 36.895000  97.875000 ;
        RECT 30.745000  97.575000 36.895000  97.725000 ;
        RECT 30.895000  97.425000 36.895000  97.575000 ;
        RECT 31.045000  97.275000 36.895000  97.425000 ;
        RECT 31.195000  97.125000 36.895000  97.275000 ;
        RECT 31.345000  96.975000 36.895000  97.125000 ;
        RECT 31.385000  92.390000 36.895000  92.540000 ;
        RECT 31.495000  96.825000 36.895000  96.975000 ;
        RECT 31.535000  92.540000 36.895000  92.690000 ;
        RECT 31.645000  96.675000 36.895000  96.825000 ;
        RECT 31.685000  92.690000 36.895000  92.840000 ;
        RECT 31.795000  96.525000 36.895000  96.675000 ;
        RECT 31.835000  92.840000 36.895000  92.990000 ;
        RECT 31.945000  92.990000 36.895000  93.100000 ;
        RECT 31.945000  93.100000 36.895000  96.375000 ;
        RECT 31.945000  96.375000 36.895000  96.525000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.835000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  1.070000  43.270000  1.400000  43.440000 ;
      RECT  1.145000  43.440000  1.315000  43.810000 ;
      RECT  3.100000  27.160000 48.200000  28.030000 ;
      RECT  3.100000  28.030000  4.020000  38.695000 ;
      RECT  3.100000  38.695000 48.200000  39.565000 ;
      RECT  3.130000  27.140000 48.200000  27.160000 ;
      RECT  3.130000  39.565000 48.200000  39.585000 ;
      RECT  4.735000  29.230000 45.955000  29.430000 ;
      RECT  4.735000  29.430000  4.905000  37.425000 ;
      RECT  4.735000  37.425000 45.955000  37.595000 ;
      RECT  6.115000  29.780000  6.285000  36.570000 ;
      RECT  6.340000  36.970000 45.060000  37.230000 ;
      RECT  6.895000  29.775000  7.065000  36.570000 ;
      RECT  7.675000  29.780000  7.845000  36.570000 ;
      RECT  8.050000  43.270000  8.690000  43.440000 ;
      RECT  8.455000  29.770000  8.625000  36.570000 ;
      RECT  8.510000 162.655000 10.360000 169.150000 ;
      RECT  9.135000  43.505000 70.125000  44.755000 ;
      RECT  9.135000  44.755000 10.385000  71.570000 ;
      RECT  9.135000  71.570000 21.085000  72.820000 ;
      RECT  9.150000 169.400000 10.400000 198.445000 ;
      RECT  9.150000 198.445000 70.125000 199.695000 ;
      RECT  9.170000 133.350000 20.990000 134.540000 ;
      RECT  9.170000 134.540000 10.360000 162.655000 ;
      RECT  9.170000 169.150000 10.360000 169.400000 ;
      RECT  9.200000 133.205000 14.190000 133.350000 ;
      RECT  9.235000  29.780000  9.405000  36.570000 ;
      RECT  9.405000  74.180000  9.935000  74.350000 ;
      RECT  9.500000  74.350000  9.830000  74.355000 ;
      RECT 10.015000  29.775000 10.185000  36.570000 ;
      RECT 10.770000 162.655000 11.975000 169.905000 ;
      RECT 10.795000  29.780000 10.965000  36.570000 ;
      RECT 11.100000 170.415000 11.990000 196.835000 ;
      RECT 11.100000 196.835000 68.155000 197.725000 ;
      RECT 11.105000  45.460000 68.155000  46.350000 ;
      RECT 11.105000  46.350000 11.995000  69.975000 ;
      RECT 11.105000  69.975000 22.680000  70.865000 ;
      RECT 11.125000 135.315000 22.660000 136.165000 ;
      RECT 11.125000 136.165000 12.100000 158.915000 ;
      RECT 11.125000 158.915000 11.975000 162.655000 ;
      RECT 11.125000 169.905000 11.975000 170.415000 ;
      RECT 11.575000  29.770000 11.745000  36.570000 ;
      RECT 12.065000   1.000000 70.650000   1.890000 ;
      RECT 12.065000   1.890000 13.045000  22.230000 ;
      RECT 12.065000  22.230000 56.085000  22.350000 ;
      RECT 12.065000  22.350000 56.105000  23.240000 ;
      RECT 12.355000  29.780000 12.525000  36.570000 ;
      RECT 12.400000 159.555000 64.500000 161.990000 ;
      RECT 12.830000 182.570000 66.685000 184.990000 ;
      RECT 13.085000  46.815000 64.500000  46.990000 ;
      RECT 13.085000  46.990000 13.255000  67.965000 ;
      RECT 13.090000  46.740000 64.500000  46.815000 ;
      RECT 13.135000  29.775000 13.305000  36.570000 ;
      RECT 13.780000   4.820000 14.010000   8.825000 ;
      RECT 13.780000   8.825000 68.570000   9.055000 ;
      RECT 13.780000  11.040000 14.010000  15.045000 ;
      RECT 13.780000  15.045000 68.570000  15.275000 ;
      RECT 13.780000  17.260000 14.010000  21.265000 ;
      RECT 13.780000  21.265000 68.570000  21.495000 ;
      RECT 13.810000   2.635000 68.540000   2.835000 ;
      RECT 13.810000   2.835000 13.980000   4.820000 ;
      RECT 13.810000   9.055000 13.980000  11.040000 ;
      RECT 13.810000  15.275000 13.980000  17.260000 ;
      RECT 13.915000  29.780000 14.085000  36.570000 ;
      RECT 13.980000   2.605000 19.570000   2.635000 ;
      RECT 14.385000  47.160000 15.435000  66.930000 ;
      RECT 14.385000 139.160000 15.435000 158.930000 ;
      RECT 14.385000 162.160000 15.435000 181.930000 ;
      RECT 14.385000 185.160000 15.435000 195.185000 ;
      RECT 14.515000   4.820000 14.745000   7.770000 ;
      RECT 14.515000  11.040000 14.745000  13.990000 ;
      RECT 14.515000  17.260000 14.745000  20.210000 ;
      RECT 14.550000   3.755000 14.720000   4.820000 ;
      RECT 14.550000   7.770000 14.720000   8.505000 ;
      RECT 14.550000   9.975000 14.720000  11.040000 ;
      RECT 14.550000  13.990000 14.720000  14.725000 ;
      RECT 14.550000  16.195000 14.720000  17.260000 ;
      RECT 14.550000  20.210000 14.720000  20.945000 ;
      RECT 14.695000  29.770000 14.865000  36.570000 ;
      RECT 14.775000   3.075000 18.775000   3.305000 ;
      RECT 14.775000   9.295000 18.775000   9.525000 ;
      RECT 14.775000  15.515000 18.775000  15.745000 ;
      RECT 15.475000  29.780000 15.645000  36.570000 ;
      RECT 15.705000  67.340000 64.500000  68.995000 ;
      RECT 15.780000 136.540000 64.500000 138.990000 ;
      RECT 15.780000 159.340000 64.500000 159.555000 ;
      RECT 15.780000 182.340000 66.685000 182.570000 ;
      RECT 15.780000 195.370000 16.490000 195.540000 ;
      RECT 16.255000  29.770000 16.425000  36.570000 ;
      RECT 16.865000  47.525000 17.395000  65.695000 ;
      RECT 16.865000 139.525000 17.395000 157.695000 ;
      RECT 16.865000 162.525000 17.395000 180.695000 ;
      RECT 16.865000 185.525000 17.395000 195.055000 ;
      RECT 16.885000  47.325000 17.395000  47.525000 ;
      RECT 16.885000  65.695000 17.395000  67.035000 ;
      RECT 16.885000 139.325000 17.395000 139.525000 ;
      RECT 16.885000 157.695000 17.395000 159.035000 ;
      RECT 16.885000 162.325000 17.395000 162.525000 ;
      RECT 16.885000 180.695000 17.395000 182.035000 ;
      RECT 16.885000 185.325000 17.395000 185.525000 ;
      RECT 17.035000  29.780000 17.205000  36.570000 ;
      RECT 17.790000 195.370000 18.500000 195.540000 ;
      RECT 17.815000  29.770000 17.985000  36.570000 ;
      RECT 17.835000 133.145000 20.990000 133.350000 ;
      RECT 18.410000  74.185000 18.740000  74.200000 ;
      RECT 18.410000  74.200000 19.000000  74.370000 ;
      RECT 18.410000  74.370000 18.740000  74.385000 ;
      RECT 18.595000  29.780000 18.765000  36.570000 ;
      RECT 18.810000   4.820000 19.040000   7.770000 ;
      RECT 18.810000  11.040000 19.040000  13.990000 ;
      RECT 18.810000  17.260000 19.040000  20.210000 ;
      RECT 18.830000   3.755000 19.000000   4.820000 ;
      RECT 18.830000   7.770000 19.000000   8.505000 ;
      RECT 18.830000   9.975000 19.000000  11.040000 ;
      RECT 18.830000  13.990000 19.000000  14.725000 ;
      RECT 18.830000  16.195000 19.000000  17.260000 ;
      RECT 18.830000  20.210000 19.000000  20.945000 ;
      RECT 18.845000  47.160000 20.035000  66.870000 ;
      RECT 18.845000 139.160000 20.035000 158.870000 ;
      RECT 18.845000 162.160000 20.035000 181.870000 ;
      RECT 18.845000 185.160000 20.035000 195.010000 ;
      RECT 18.985000 195.010000 19.875000 195.075000 ;
      RECT 19.375000  29.775000 19.545000  36.570000 ;
      RECT 19.540000   4.820000 19.770000   8.825000 ;
      RECT 19.540000  11.040000 19.770000  15.045000 ;
      RECT 19.540000  17.260000 19.770000  21.265000 ;
      RECT 19.565000  97.500000 20.990000 133.145000 ;
      RECT 19.570000   2.835000 19.740000   4.820000 ;
      RECT 19.570000   9.055000 19.740000  11.040000 ;
      RECT 19.570000  15.275000 19.740000  17.260000 ;
      RECT 19.740000   2.605000 29.330000   2.635000 ;
      RECT 19.800000  72.820000 21.085000  96.895000 ;
      RECT 19.800000  96.895000 20.990000  97.500000 ;
      RECT 20.155000  29.780000 20.325000  36.570000 ;
      RECT 20.275000   4.820000 20.505000   7.770000 ;
      RECT 20.275000  11.040000 20.505000  13.990000 ;
      RECT 20.275000  17.260000 20.505000  20.210000 ;
      RECT 20.310000   3.755000 20.480000   4.820000 ;
      RECT 20.310000   7.770000 20.480000   8.505000 ;
      RECT 20.310000   9.975000 20.480000  11.040000 ;
      RECT 20.310000  13.990000 20.480000  14.725000 ;
      RECT 20.310000  16.195000 20.480000  17.260000 ;
      RECT 20.310000  20.210000 20.480000  20.945000 ;
      RECT 20.380000 195.370000 21.090000 195.540000 ;
      RECT 20.535000   3.075000 28.535000   3.305000 ;
      RECT 20.535000   9.295000 28.535000   9.525000 ;
      RECT 20.535000  15.515000 28.535000  15.745000 ;
      RECT 20.935000  29.770000 21.105000  36.570000 ;
      RECT 21.465000  47.525000 21.995000  65.695000 ;
      RECT 21.465000 139.525000 21.995000 157.695000 ;
      RECT 21.465000 162.525000 21.995000 180.695000 ;
      RECT 21.465000 185.525000 21.995000 195.055000 ;
      RECT 21.485000  47.325000 21.995000  47.525000 ;
      RECT 21.485000  65.695000 21.995000  67.035000 ;
      RECT 21.485000 139.325000 21.995000 139.525000 ;
      RECT 21.485000 157.695000 21.995000 159.035000 ;
      RECT 21.485000 162.325000 21.995000 162.525000 ;
      RECT 21.485000 180.695000 21.995000 182.035000 ;
      RECT 21.485000 185.325000 21.995000 185.525000 ;
      RECT 21.715000  29.780000 21.885000  36.570000 ;
      RECT 21.790000  70.865000 22.680000  97.450000 ;
      RECT 21.810000  97.450000 22.660000 135.315000 ;
      RECT 22.390000 195.370000 23.100000 195.540000 ;
      RECT 22.495000  29.775000 22.665000  36.570000 ;
      RECT 23.025000  90.495000 64.500000  92.990000 ;
      RECT 23.055000 113.340000 64.500000 115.990000 ;
      RECT 23.275000  29.780000 23.445000  36.570000 ;
      RECT 23.445000  47.160000 24.635000  66.870000 ;
      RECT 23.445000 139.160000 24.635000 158.870000 ;
      RECT 23.445000 162.160000 24.635000 181.870000 ;
      RECT 23.445000 185.160000 24.635000 195.010000 ;
      RECT 23.510000  68.995000 64.500000  69.990000 ;
      RECT 23.585000  70.160000 24.635000  89.930000 ;
      RECT 23.585000  93.160000 24.635000 112.930000 ;
      RECT 23.585000 116.160000 24.635000 135.930000 ;
      RECT 23.585000 195.010000 24.475000 195.030000 ;
      RECT 24.055000  29.770000 24.225000  36.570000 ;
      RECT 24.835000  29.780000 25.005000  36.570000 ;
      RECT 24.980000  90.370000 64.500000  90.495000 ;
      RECT 24.980000 136.370000 64.500000 136.540000 ;
      RECT 24.980000 195.370000 25.690000 195.540000 ;
      RECT 25.615000  29.775000 25.785000  36.570000 ;
      RECT 25.670000  90.340000 64.500000  90.370000 ;
      RECT 25.670000 136.340000 64.500000 136.370000 ;
      RECT 26.065000  47.525000 26.595000  65.695000 ;
      RECT 26.065000  70.525000 26.595000  88.695000 ;
      RECT 26.065000  93.525000 26.595000 111.695000 ;
      RECT 26.065000 116.525000 26.595000 134.695000 ;
      RECT 26.065000 139.525000 26.595000 157.695000 ;
      RECT 26.065000 162.525000 26.595000 180.695000 ;
      RECT 26.065000 185.525000 26.595000 195.055000 ;
      RECT 26.085000  47.325000 26.595000  47.525000 ;
      RECT 26.085000  65.695000 26.595000  67.035000 ;
      RECT 26.085000  70.325000 26.595000  70.525000 ;
      RECT 26.085000  88.695000 26.595000  90.035000 ;
      RECT 26.085000  93.325000 26.595000  93.525000 ;
      RECT 26.085000 111.695000 26.595000 113.035000 ;
      RECT 26.085000 116.325000 26.595000 116.525000 ;
      RECT 26.085000 134.695000 26.595000 136.035000 ;
      RECT 26.085000 139.325000 26.595000 139.525000 ;
      RECT 26.085000 157.695000 26.595000 159.035000 ;
      RECT 26.085000 162.325000 26.595000 162.525000 ;
      RECT 26.085000 180.695000 26.595000 182.035000 ;
      RECT 26.085000 185.325000 26.595000 185.525000 ;
      RECT 26.395000  29.780000 26.565000  36.570000 ;
      RECT 26.990000 195.370000 27.700000 195.540000 ;
      RECT 27.175000  29.770000 27.345000  36.570000 ;
      RECT 27.955000  29.780000 28.125000  36.570000 ;
      RECT 28.045000  47.160000 29.235000  66.870000 ;
      RECT 28.045000  70.160000 29.235000  89.870000 ;
      RECT 28.045000  93.160000 29.235000 112.870000 ;
      RECT 28.045000 116.160000 29.235000 135.870000 ;
      RECT 28.045000 139.160000 29.235000 158.870000 ;
      RECT 28.045000 162.160000 29.235000 181.870000 ;
      RECT 28.045000 185.160000 29.235000 195.010000 ;
      RECT 28.185000 195.010000 29.075000 195.030000 ;
      RECT 28.570000   4.820000 28.800000   7.770000 ;
      RECT 28.570000  11.040000 28.800000  13.990000 ;
      RECT 28.570000  17.260000 28.800000  20.210000 ;
      RECT 28.590000   3.755000 28.760000   4.820000 ;
      RECT 28.590000   7.770000 28.760000   8.505000 ;
      RECT 28.590000   9.975000 28.760000  11.040000 ;
      RECT 28.590000  13.990000 28.760000  14.725000 ;
      RECT 28.590000  16.195000 28.760000  17.260000 ;
      RECT 28.590000  20.210000 28.760000  20.945000 ;
      RECT 28.735000  29.775000 28.905000  36.570000 ;
      RECT 29.300000   4.820000 29.530000   8.825000 ;
      RECT 29.300000  11.040000 29.530000  15.045000 ;
      RECT 29.300000  17.260000 29.530000  21.265000 ;
      RECT 29.330000   2.835000 29.500000   4.820000 ;
      RECT 29.330000   9.055000 29.500000  11.040000 ;
      RECT 29.330000  15.275000 29.500000  17.260000 ;
      RECT 29.500000   2.605000 39.090000   2.635000 ;
      RECT 29.515000  29.780000 29.685000  36.570000 ;
      RECT 29.580000 195.370000 30.290000 195.540000 ;
      RECT 30.035000   4.820000 30.265000   7.770000 ;
      RECT 30.035000  11.040000 30.265000  13.990000 ;
      RECT 30.035000  17.260000 30.265000  20.210000 ;
      RECT 30.070000   3.755000 30.240000   4.820000 ;
      RECT 30.070000   7.770000 30.240000   8.505000 ;
      RECT 30.070000   9.975000 30.240000  11.040000 ;
      RECT 30.070000  13.990000 30.240000  14.725000 ;
      RECT 30.070000  16.195000 30.240000  17.260000 ;
      RECT 30.070000  20.210000 30.240000  20.945000 ;
      RECT 30.295000   3.075000 38.295000   3.305000 ;
      RECT 30.295000   9.295000 38.295000   9.525000 ;
      RECT 30.295000  15.515000 38.295000  15.745000 ;
      RECT 30.295000  29.770000 30.465000  36.570000 ;
      RECT 30.665000  47.525000 31.195000  65.695000 ;
      RECT 30.665000  70.525000 31.195000  88.695000 ;
      RECT 30.665000  93.525000 31.195000 111.695000 ;
      RECT 30.665000 116.525000 31.195000 134.695000 ;
      RECT 30.665000 139.525000 31.195000 157.695000 ;
      RECT 30.665000 162.525000 31.195000 180.695000 ;
      RECT 30.665000 185.525000 31.195000 195.055000 ;
      RECT 30.685000  47.325000 31.195000  47.525000 ;
      RECT 30.685000  65.695000 31.195000  67.035000 ;
      RECT 30.685000  70.325000 31.195000  70.525000 ;
      RECT 30.685000  88.695000 31.195000  90.035000 ;
      RECT 30.685000  93.325000 31.195000  93.525000 ;
      RECT 30.685000 111.695000 31.195000 113.035000 ;
      RECT 30.685000 116.325000 31.195000 116.525000 ;
      RECT 30.685000 134.695000 31.195000 136.035000 ;
      RECT 30.685000 139.325000 31.195000 139.525000 ;
      RECT 30.685000 157.695000 31.195000 159.035000 ;
      RECT 30.685000 162.325000 31.195000 162.525000 ;
      RECT 30.685000 180.695000 31.195000 182.035000 ;
      RECT 30.685000 185.325000 31.195000 185.525000 ;
      RECT 31.075000  29.780000 31.245000  36.570000 ;
      RECT 31.590000 195.370000 32.300000 195.540000 ;
      RECT 31.855000  29.775000 32.025000  36.570000 ;
      RECT 32.635000  29.780000 32.805000  36.570000 ;
      RECT 32.645000  47.160000 33.835000  66.870000 ;
      RECT 32.645000  70.160000 33.835000  89.870000 ;
      RECT 32.645000  93.160000 33.835000 112.870000 ;
      RECT 32.645000 116.160000 33.835000 135.870000 ;
      RECT 32.645000 139.160000 33.835000 158.870000 ;
      RECT 32.645000 162.160000 33.835000 181.870000 ;
      RECT 32.645000 185.160000 33.835000 195.010000 ;
      RECT 32.785000 195.010000 33.675000 195.030000 ;
      RECT 33.415000  29.770000 33.585000  36.570000 ;
      RECT 34.180000 195.370000 34.890000 195.540000 ;
      RECT 34.195000  29.780000 34.365000  36.570000 ;
      RECT 34.975000  29.775000 35.145000  36.570000 ;
      RECT 35.265000  47.525000 35.795000  65.695000 ;
      RECT 35.265000  70.525000 35.795000  88.695000 ;
      RECT 35.265000  93.525000 35.795000 111.695000 ;
      RECT 35.265000 116.525000 35.795000 134.695000 ;
      RECT 35.265000 139.525000 35.795000 157.695000 ;
      RECT 35.265000 162.525000 35.795000 180.695000 ;
      RECT 35.265000 185.525000 35.795000 195.055000 ;
      RECT 35.285000  47.325000 35.795000  47.525000 ;
      RECT 35.285000  65.695000 35.795000  67.035000 ;
      RECT 35.285000  70.325000 35.795000  70.525000 ;
      RECT 35.285000  88.695000 35.795000  90.035000 ;
      RECT 35.285000  93.325000 35.795000  93.525000 ;
      RECT 35.285000 111.695000 35.795000 113.035000 ;
      RECT 35.285000 116.325000 35.795000 116.525000 ;
      RECT 35.285000 134.695000 35.795000 136.035000 ;
      RECT 35.285000 139.325000 35.795000 139.525000 ;
      RECT 35.285000 157.695000 35.795000 159.035000 ;
      RECT 35.285000 162.325000 35.795000 162.525000 ;
      RECT 35.285000 180.695000 35.795000 182.035000 ;
      RECT 35.285000 185.325000 35.795000 185.525000 ;
      RECT 35.755000  29.780000 35.925000  36.570000 ;
      RECT 36.190000 195.370000 36.900000 195.540000 ;
      RECT 36.535000  29.770000 36.705000  36.570000 ;
      RECT 37.245000  47.160000 38.435000  66.870000 ;
      RECT 37.245000  70.160000 38.435000  89.870000 ;
      RECT 37.245000  93.160000 38.435000 112.870000 ;
      RECT 37.245000 116.160000 38.435000 135.870000 ;
      RECT 37.245000 139.160000 38.435000 158.870000 ;
      RECT 37.245000 162.160000 38.435000 181.870000 ;
      RECT 37.245000 185.160000 38.435000 195.010000 ;
      RECT 37.315000  29.780000 37.485000  36.570000 ;
      RECT 37.385000 195.010000 38.275000 195.030000 ;
      RECT 38.095000  29.775000 38.265000  36.570000 ;
      RECT 38.330000   4.820000 38.560000   7.770000 ;
      RECT 38.330000  11.040000 38.560000  13.990000 ;
      RECT 38.330000  17.260000 38.560000  20.210000 ;
      RECT 38.350000   3.755000 38.520000   4.820000 ;
      RECT 38.350000   7.770000 38.520000   8.505000 ;
      RECT 38.350000   9.975000 38.520000  11.040000 ;
      RECT 38.350000  13.990000 38.520000  14.725000 ;
      RECT 38.350000  16.195000 38.520000  17.260000 ;
      RECT 38.350000  20.210000 38.520000  20.945000 ;
      RECT 38.780000 195.370000 39.490000 195.540000 ;
      RECT 38.875000  29.780000 39.045000  36.570000 ;
      RECT 39.060000   4.820000 39.290000   8.825000 ;
      RECT 39.060000  11.040000 39.290000  15.045000 ;
      RECT 39.060000  17.260000 39.290000  21.265000 ;
      RECT 39.090000   2.835000 39.260000   4.820000 ;
      RECT 39.090000   9.055000 39.260000  11.040000 ;
      RECT 39.090000  15.275000 39.260000  17.260000 ;
      RECT 39.260000   2.605000 48.850000   2.635000 ;
      RECT 39.655000  29.770000 39.825000  36.570000 ;
      RECT 39.795000   4.820000 40.025000   7.770000 ;
      RECT 39.795000  11.040000 40.025000  13.990000 ;
      RECT 39.795000  17.260000 40.025000  20.210000 ;
      RECT 39.830000   3.755000 40.000000   4.820000 ;
      RECT 39.830000   7.770000 40.000000   8.505000 ;
      RECT 39.830000   9.975000 40.000000  11.040000 ;
      RECT 39.830000  13.990000 40.000000  14.725000 ;
      RECT 39.830000  16.195000 40.000000  17.260000 ;
      RECT 39.830000  20.210000 40.000000  20.945000 ;
      RECT 39.865000  47.525000 40.395000  65.695000 ;
      RECT 39.865000  70.525000 40.395000  88.695000 ;
      RECT 39.865000  93.525000 40.395000 111.695000 ;
      RECT 39.865000 116.525000 40.395000 134.695000 ;
      RECT 39.865000 139.525000 40.395000 157.695000 ;
      RECT 39.865000 162.525000 40.395000 180.695000 ;
      RECT 39.865000 185.525000 40.395000 195.055000 ;
      RECT 39.885000  47.325000 40.395000  47.525000 ;
      RECT 39.885000  65.695000 40.395000  67.035000 ;
      RECT 39.885000  70.325000 40.395000  70.525000 ;
      RECT 39.885000  88.695000 40.395000  90.035000 ;
      RECT 39.885000  93.325000 40.395000  93.525000 ;
      RECT 39.885000 111.695000 40.395000 113.035000 ;
      RECT 39.885000 116.325000 40.395000 116.525000 ;
      RECT 39.885000 134.695000 40.395000 136.035000 ;
      RECT 39.885000 139.325000 40.395000 139.525000 ;
      RECT 39.885000 157.695000 40.395000 159.035000 ;
      RECT 39.885000 162.325000 40.395000 162.525000 ;
      RECT 39.885000 180.695000 40.395000 182.035000 ;
      RECT 39.885000 185.325000 40.395000 185.525000 ;
      RECT 40.055000   3.075000 48.055000   3.305000 ;
      RECT 40.055000   9.295000 48.055000   9.525000 ;
      RECT 40.055000  15.515000 48.055000  15.745000 ;
      RECT 40.435000  29.780000 40.605000  36.570000 ;
      RECT 40.790000 195.370000 41.500000 195.540000 ;
      RECT 41.215000  29.770000 41.385000  36.570000 ;
      RECT 41.845000  47.160000 43.035000  66.870000 ;
      RECT 41.845000  70.160000 43.035000  89.870000 ;
      RECT 41.845000  93.160000 43.035000 112.870000 ;
      RECT 41.845000 116.160000 43.035000 135.870000 ;
      RECT 41.845000 139.160000 43.035000 158.870000 ;
      RECT 41.845000 162.160000 43.035000 181.870000 ;
      RECT 41.845000 185.160000 43.035000 195.010000 ;
      RECT 41.985000 195.010000 42.875000 195.030000 ;
      RECT 41.995000  29.780000 42.165000  36.570000 ;
      RECT 42.775000  29.775000 42.945000  36.570000 ;
      RECT 43.380000 195.370000 44.090000 195.540000 ;
      RECT 43.555000  29.780000 43.725000  36.570000 ;
      RECT 44.335000  29.770000 44.505000  36.570000 ;
      RECT 44.465000  47.525000 44.995000  65.695000 ;
      RECT 44.465000  70.525000 44.995000  88.695000 ;
      RECT 44.465000  93.525000 44.995000 111.695000 ;
      RECT 44.465000 116.525000 44.995000 134.695000 ;
      RECT 44.465000 139.525000 44.995000 157.695000 ;
      RECT 44.465000 162.525000 44.995000 180.695000 ;
      RECT 44.465000 185.525000 44.995000 195.055000 ;
      RECT 44.485000  47.325000 44.995000  47.525000 ;
      RECT 44.485000  65.695000 44.995000  67.035000 ;
      RECT 44.485000  70.325000 44.995000  70.525000 ;
      RECT 44.485000  88.695000 44.995000  90.035000 ;
      RECT 44.485000  93.325000 44.995000  93.525000 ;
      RECT 44.485000 111.695000 44.995000 113.035000 ;
      RECT 44.485000 116.325000 44.995000 116.525000 ;
      RECT 44.485000 134.695000 44.995000 136.035000 ;
      RECT 44.485000 139.325000 44.995000 139.525000 ;
      RECT 44.485000 157.695000 44.995000 159.035000 ;
      RECT 44.485000 162.325000 44.995000 162.525000 ;
      RECT 44.485000 180.695000 44.995000 182.035000 ;
      RECT 44.485000 185.325000 44.995000 185.525000 ;
      RECT 45.115000  29.780000 45.285000  36.570000 ;
      RECT 45.390000 195.370000 46.100000 195.540000 ;
      RECT 45.755000  29.430000 45.955000  37.425000 ;
      RECT 46.445000  47.160000 47.635000  66.870000 ;
      RECT 46.445000  70.160000 47.635000  89.870000 ;
      RECT 46.445000  93.160000 47.635000 112.870000 ;
      RECT 46.445000 116.160000 47.635000 135.870000 ;
      RECT 46.445000 139.160000 47.635000 158.870000 ;
      RECT 46.445000 162.160000 47.635000 181.870000 ;
      RECT 46.445000 185.160000 47.635000 195.010000 ;
      RECT 46.585000 195.010000 47.475000 195.030000 ;
      RECT 47.310000  28.030000 48.200000  29.215000 ;
      RECT 47.310000  29.525000 48.200000  38.695000 ;
      RECT 47.330000  29.215000 48.180000  29.525000 ;
      RECT 47.980000 195.370000 48.690000 195.540000 ;
      RECT 48.090000   4.820000 48.320000   7.770000 ;
      RECT 48.090000  11.040000 48.320000  13.990000 ;
      RECT 48.090000  17.260000 48.320000  20.210000 ;
      RECT 48.110000   3.755000 48.280000   4.820000 ;
      RECT 48.110000   7.770000 48.280000   8.505000 ;
      RECT 48.110000   9.975000 48.280000  11.040000 ;
      RECT 48.110000  13.990000 48.280000  14.725000 ;
      RECT 48.110000  16.195000 48.280000  17.260000 ;
      RECT 48.110000  20.210000 48.280000  20.945000 ;
      RECT 48.820000   4.820000 49.050000   8.825000 ;
      RECT 48.820000  11.040000 49.050000  15.045000 ;
      RECT 48.820000  17.260000 49.050000  21.265000 ;
      RECT 48.850000   2.835000 49.020000   4.820000 ;
      RECT 48.850000   9.055000 49.020000  11.040000 ;
      RECT 48.850000  15.275000 49.020000  17.260000 ;
      RECT 49.020000   2.605000 58.610000   2.635000 ;
      RECT 49.065000  47.525000 49.595000  65.695000 ;
      RECT 49.065000  70.525000 49.595000  88.695000 ;
      RECT 49.065000  93.525000 49.595000 111.695000 ;
      RECT 49.065000 116.525000 49.595000 134.695000 ;
      RECT 49.065000 139.525000 49.595000 157.695000 ;
      RECT 49.065000 162.525000 49.595000 180.695000 ;
      RECT 49.065000 185.525000 49.595000 195.055000 ;
      RECT 49.085000  47.325000 49.595000  47.525000 ;
      RECT 49.085000  65.695000 49.595000  67.035000 ;
      RECT 49.085000  70.325000 49.595000  70.525000 ;
      RECT 49.085000  88.695000 49.595000  90.035000 ;
      RECT 49.085000  93.325000 49.595000  93.525000 ;
      RECT 49.085000 111.695000 49.595000 113.035000 ;
      RECT 49.085000 116.325000 49.595000 116.525000 ;
      RECT 49.085000 134.695000 49.595000 136.035000 ;
      RECT 49.085000 139.325000 49.595000 139.525000 ;
      RECT 49.085000 157.695000 49.595000 159.035000 ;
      RECT 49.085000 162.325000 49.595000 162.525000 ;
      RECT 49.085000 180.695000 49.595000 182.035000 ;
      RECT 49.085000 185.325000 49.595000 185.525000 ;
      RECT 49.555000   4.820000 49.785000   7.770000 ;
      RECT 49.555000  11.040000 49.785000  13.990000 ;
      RECT 49.555000  17.260000 49.785000  20.210000 ;
      RECT 49.590000   3.755000 49.760000   4.820000 ;
      RECT 49.590000   7.770000 49.760000   8.505000 ;
      RECT 49.590000   9.975000 49.760000  11.040000 ;
      RECT 49.590000  13.990000 49.760000  14.725000 ;
      RECT 49.590000  16.195000 49.760000  17.260000 ;
      RECT 49.590000  20.210000 49.760000  20.945000 ;
      RECT 49.815000   3.075000 57.815000   3.305000 ;
      RECT 49.815000   9.295000 57.815000   9.525000 ;
      RECT 49.815000  15.515000 57.815000  15.745000 ;
      RECT 49.990000 195.370000 50.700000 195.540000 ;
      RECT 51.045000  47.160000 52.235000  66.870000 ;
      RECT 51.045000  70.160000 52.235000  89.870000 ;
      RECT 51.045000  93.160000 52.235000 112.870000 ;
      RECT 51.045000 116.160000 52.235000 135.870000 ;
      RECT 51.045000 139.160000 52.235000 158.870000 ;
      RECT 51.045000 162.160000 52.235000 181.870000 ;
      RECT 51.045000 185.160000 52.235000 195.010000 ;
      RECT 51.185000 195.010000 52.075000 195.030000 ;
      RECT 52.320000  29.300000 68.865000  31.060000 ;
      RECT 52.320000  31.060000 53.210000  41.455000 ;
      RECT 52.320000  41.455000 68.865000  42.495000 ;
      RECT 52.580000 195.370000 53.290000 195.540000 ;
      RECT 53.665000  47.525000 54.195000  65.695000 ;
      RECT 53.665000  70.525000 54.195000  88.695000 ;
      RECT 53.665000  93.525000 54.195000 111.695000 ;
      RECT 53.665000 116.525000 54.195000 134.695000 ;
      RECT 53.665000 139.525000 54.195000 157.695000 ;
      RECT 53.665000 162.525000 54.195000 180.695000 ;
      RECT 53.665000 185.525000 54.195000 195.055000 ;
      RECT 53.685000  47.325000 54.195000  47.525000 ;
      RECT 53.685000  65.695000 54.195000  67.035000 ;
      RECT 53.685000  70.325000 54.195000  70.525000 ;
      RECT 53.685000  88.695000 54.195000  90.035000 ;
      RECT 53.685000  93.325000 54.195000  93.525000 ;
      RECT 53.685000 111.695000 54.195000 113.035000 ;
      RECT 53.685000 116.325000 54.195000 116.525000 ;
      RECT 53.685000 134.695000 54.195000 136.035000 ;
      RECT 53.685000 139.325000 54.195000 139.525000 ;
      RECT 53.685000 157.695000 54.195000 159.035000 ;
      RECT 53.685000 162.325000 54.195000 162.525000 ;
      RECT 53.685000 180.695000 54.195000 182.035000 ;
      RECT 53.685000 185.325000 54.195000 185.525000 ;
      RECT 53.960000  31.835000 67.140000  32.005000 ;
      RECT 53.960000  32.005000 54.130000  40.410000 ;
      RECT 53.960000  40.410000 67.140000  40.580000 ;
      RECT 54.590000 195.370000 55.300000 195.540000 ;
      RECT 54.690000  32.560000 54.860000  36.190000 ;
      RECT 54.690000  36.190000 54.865000  39.290000 ;
      RECT 54.690000  39.290000 54.860000  39.350000 ;
      RECT 54.940000  39.770000 66.335000  39.940000 ;
      RECT 55.215000  23.240000 56.105000  28.345000 ;
      RECT 55.215000  28.345000 70.630000  29.300000 ;
      RECT 55.465000  32.620000 55.640000  35.770000 ;
      RECT 55.470000  32.560000 55.640000  32.620000 ;
      RECT 55.470000  35.770000 55.640000  39.350000 ;
      RECT 55.645000  47.160000 56.835000  66.870000 ;
      RECT 55.645000  70.160000 56.835000  89.870000 ;
      RECT 55.645000  93.160000 56.835000 112.870000 ;
      RECT 55.645000 116.160000 56.835000 135.870000 ;
      RECT 55.645000 139.160000 56.835000 158.870000 ;
      RECT 55.645000 162.160000 56.835000 181.870000 ;
      RECT 55.645000 185.160000 56.835000 195.010000 ;
      RECT 55.785000 195.010000 56.675000 195.140000 ;
      RECT 56.250000  32.560000 56.420000  36.190000 ;
      RECT 56.250000  36.190000 56.425000  39.290000 ;
      RECT 56.250000  39.290000 56.420000  39.350000 ;
      RECT 56.820000  23.480000 57.050000  27.485000 ;
      RECT 56.820000  27.485000 68.570000  27.715000 ;
      RECT 56.850000  21.495000 57.020000  23.480000 ;
      RECT 57.025000  32.620000 57.200000  35.770000 ;
      RECT 57.030000  32.560000 57.200000  32.620000 ;
      RECT 57.030000  35.770000 57.200000  39.350000 ;
      RECT 57.180000 195.370000 57.890000 195.540000 ;
      RECT 57.555000  23.480000 57.785000  26.430000 ;
      RECT 57.590000  22.415000 57.760000  23.480000 ;
      RECT 57.590000  26.430000 57.760000  27.165000 ;
      RECT 57.810000  32.560000 57.980000  36.190000 ;
      RECT 57.810000  36.190000 57.985000  39.290000 ;
      RECT 57.810000  39.290000 57.980000  39.350000 ;
      RECT 57.815000  21.735000 61.815000  21.965000 ;
      RECT 57.850000   4.820000 58.080000   7.770000 ;
      RECT 57.850000  11.040000 58.080000  13.990000 ;
      RECT 57.850000  17.260000 58.080000  20.210000 ;
      RECT 57.870000   3.755000 58.040000   4.820000 ;
      RECT 57.870000   7.770000 58.040000   8.505000 ;
      RECT 57.870000   9.975000 58.040000  11.040000 ;
      RECT 57.870000  13.990000 58.040000  14.725000 ;
      RECT 57.870000  16.195000 58.040000  17.260000 ;
      RECT 57.870000  20.210000 58.040000  20.945000 ;
      RECT 58.265000  47.525000 58.795000  65.695000 ;
      RECT 58.265000  70.525000 58.795000  88.695000 ;
      RECT 58.265000  93.525000 58.795000 111.695000 ;
      RECT 58.265000 116.525000 58.795000 134.695000 ;
      RECT 58.265000 139.525000 58.795000 157.695000 ;
      RECT 58.265000 162.525000 58.795000 180.695000 ;
      RECT 58.265000 185.525000 58.795000 195.055000 ;
      RECT 58.285000  47.325000 58.795000  47.525000 ;
      RECT 58.285000  65.695000 58.795000  67.035000 ;
      RECT 58.285000  70.325000 58.795000  70.525000 ;
      RECT 58.285000  88.695000 58.795000  90.035000 ;
      RECT 58.285000  93.325000 58.795000  93.525000 ;
      RECT 58.285000 111.695000 58.795000 113.035000 ;
      RECT 58.285000 116.325000 58.795000 116.525000 ;
      RECT 58.285000 134.695000 58.795000 136.035000 ;
      RECT 58.285000 139.325000 58.795000 139.525000 ;
      RECT 58.285000 157.695000 58.795000 159.035000 ;
      RECT 58.285000 162.325000 58.795000 162.525000 ;
      RECT 58.285000 180.695000 58.795000 182.035000 ;
      RECT 58.285000 185.325000 58.795000 185.525000 ;
      RECT 58.580000   4.820000 58.810000   8.825000 ;
      RECT 58.580000  11.040000 58.810000  15.045000 ;
      RECT 58.580000  17.260000 58.810000  21.265000 ;
      RECT 58.585000  32.620000 58.760000  35.770000 ;
      RECT 58.590000  32.560000 58.760000  32.620000 ;
      RECT 58.590000  35.770000 58.760000  39.350000 ;
      RECT 58.610000   2.835000 58.780000   4.820000 ;
      RECT 58.610000   9.055000 58.780000  11.040000 ;
      RECT 58.610000  15.275000 58.780000  17.260000 ;
      RECT 58.780000   2.605000 68.370000   2.635000 ;
      RECT 59.190000 195.370000 59.900000 195.540000 ;
      RECT 59.315000   4.820000 59.545000   7.770000 ;
      RECT 59.315000  11.040000 59.545000  13.990000 ;
      RECT 59.315000  17.260000 59.545000  20.210000 ;
      RECT 59.350000   3.755000 59.520000   4.820000 ;
      RECT 59.350000   7.770000 59.520000   8.505000 ;
      RECT 59.350000   9.975000 59.520000  11.040000 ;
      RECT 59.350000  13.990000 59.520000  14.725000 ;
      RECT 59.350000  16.195000 59.520000  17.260000 ;
      RECT 59.350000  20.210000 59.520000  20.945000 ;
      RECT 59.370000  32.560000 59.540000  36.190000 ;
      RECT 59.370000  36.190000 59.545000  39.290000 ;
      RECT 59.370000  39.290000 59.540000  39.350000 ;
      RECT 59.575000   3.075000 67.575000   3.305000 ;
      RECT 59.575000   9.295000 67.575000   9.525000 ;
      RECT 59.575000  15.515000 67.575000  15.745000 ;
      RECT 60.145000  32.620000 60.320000  35.770000 ;
      RECT 60.150000  32.560000 60.320000  32.620000 ;
      RECT 60.150000  35.770000 60.320000  39.350000 ;
      RECT 60.245000  47.160000 61.435000  66.870000 ;
      RECT 60.245000  70.160000 61.435000  89.870000 ;
      RECT 60.245000  93.160000 61.435000 112.870000 ;
      RECT 60.245000 116.160000 61.435000 135.870000 ;
      RECT 60.245000 139.160000 61.435000 158.870000 ;
      RECT 60.245000 162.160000 61.435000 181.870000 ;
      RECT 60.245000 185.160000 61.435000 195.010000 ;
      RECT 60.385000 195.010000 61.275000 195.140000 ;
      RECT 60.930000  32.560000 61.100000  36.190000 ;
      RECT 60.930000  36.190000 61.105000  39.290000 ;
      RECT 60.930000  39.290000 61.100000  39.350000 ;
      RECT 61.705000  32.620000 61.880000  35.770000 ;
      RECT 61.710000  32.560000 61.880000  32.620000 ;
      RECT 61.710000  35.770000 61.880000  39.350000 ;
      RECT 61.780000 195.370000 62.490000 195.540000 ;
      RECT 61.850000  23.480000 62.080000  26.430000 ;
      RECT 61.870000  22.415000 62.040000  23.480000 ;
      RECT 61.870000  26.430000 62.040000  27.165000 ;
      RECT 62.490000  32.560000 62.660000  36.190000 ;
      RECT 62.490000  36.190000 62.665000  39.290000 ;
      RECT 62.490000  39.290000 62.660000  39.350000 ;
      RECT 62.580000  23.480000 62.810000  27.485000 ;
      RECT 62.610000  21.495000 62.780000  23.480000 ;
      RECT 62.865000  47.525000 63.395000  65.695000 ;
      RECT 62.865000  70.525000 63.395000  88.695000 ;
      RECT 62.865000  93.525000 63.395000 111.695000 ;
      RECT 62.865000 116.525000 63.395000 134.695000 ;
      RECT 62.865000 139.525000 63.395000 157.695000 ;
      RECT 62.865000 162.525000 63.395000 180.695000 ;
      RECT 62.865000 185.525000 63.395000 195.055000 ;
      RECT 62.885000  47.325000 63.395000  47.525000 ;
      RECT 62.885000  65.695000 63.395000  67.035000 ;
      RECT 62.885000  70.325000 63.395000  70.525000 ;
      RECT 62.885000  88.695000 63.395000  90.035000 ;
      RECT 62.885000  93.325000 63.395000  93.525000 ;
      RECT 62.885000 111.695000 63.395000 113.035000 ;
      RECT 62.885000 116.325000 63.395000 116.525000 ;
      RECT 62.885000 134.695000 63.395000 136.035000 ;
      RECT 62.885000 139.325000 63.395000 139.525000 ;
      RECT 62.885000 157.695000 63.395000 159.035000 ;
      RECT 62.885000 162.325000 63.395000 162.525000 ;
      RECT 62.885000 180.695000 63.395000 182.035000 ;
      RECT 62.885000 185.325000 63.395000 185.525000 ;
      RECT 63.265000  32.620000 63.440000  35.770000 ;
      RECT 63.270000  32.560000 63.440000  32.620000 ;
      RECT 63.270000  35.770000 63.440000  39.350000 ;
      RECT 63.315000  23.480000 63.545000  26.430000 ;
      RECT 63.350000  22.415000 63.520000  23.480000 ;
      RECT 63.350000  26.430000 63.520000  27.165000 ;
      RECT 63.575000  21.735000 67.575000  21.965000 ;
      RECT 63.790000 195.370000 64.500000 195.540000 ;
      RECT 64.050000  32.560000 64.220000  36.190000 ;
      RECT 64.050000  36.190000 64.225000  39.290000 ;
      RECT 64.050000  39.290000 64.220000  39.350000 ;
      RECT 64.825000  32.620000 65.000000  35.770000 ;
      RECT 64.830000  32.560000 65.000000  32.620000 ;
      RECT 64.830000  35.770000 65.000000  39.350000 ;
      RECT 64.845000  47.160000 65.875000  66.930000 ;
      RECT 64.845000  70.160000 65.875000  89.930000 ;
      RECT 64.845000  93.160000 65.875000 112.935000 ;
      RECT 64.845000 116.160000 65.875000 135.930000 ;
      RECT 64.845000 139.160000 65.875000 158.930000 ;
      RECT 64.845000 162.160000 65.875000 181.930000 ;
      RECT 64.845000 185.160000 65.875000 195.180000 ;
      RECT 65.610000  32.560000 65.780000  36.190000 ;
      RECT 65.610000  36.190000 65.785000  39.290000 ;
      RECT 65.610000  39.290000 65.780000  39.350000 ;
      RECT 66.385000  32.620000 66.560000  35.770000 ;
      RECT 66.390000  32.560000 66.560000  32.620000 ;
      RECT 66.390000  35.770000 66.560000  39.350000 ;
      RECT 66.935000  32.005000 67.140000  36.065000 ;
      RECT 66.935000  36.275000 67.140000  40.410000 ;
      RECT 66.970000  36.065000 67.140000  36.275000 ;
      RECT 67.265000  46.350000 68.155000 101.315000 ;
      RECT 67.265000 166.045000 68.155000 196.835000 ;
      RECT 67.290000 101.315000 68.140000 101.710000 ;
      RECT 67.290000 101.710000 68.155000 165.645000 ;
      RECT 67.290000 165.645000 68.140000 166.045000 ;
      RECT 67.610000   4.820000 67.840000   7.770000 ;
      RECT 67.610000  11.040000 67.840000  13.990000 ;
      RECT 67.610000  17.260000 67.840000  20.210000 ;
      RECT 67.610000  23.480000 67.840000  26.430000 ;
      RECT 67.630000   3.755000 67.800000   4.820000 ;
      RECT 67.630000   7.770000 67.800000   8.505000 ;
      RECT 67.630000   9.975000 67.800000  11.040000 ;
      RECT 67.630000  13.990000 67.800000  14.725000 ;
      RECT 67.630000  16.195000 67.800000  17.260000 ;
      RECT 67.630000  20.210000 67.800000  20.945000 ;
      RECT 67.630000  22.415000 67.800000  23.480000 ;
      RECT 67.630000  26.430000 67.800000  27.165000 ;
      RECT 67.975000  31.060000 68.865000  40.480000 ;
      RECT 67.975000  41.315000 68.865000  41.455000 ;
      RECT 68.000000  40.480000 68.830000  41.315000 ;
      RECT 68.340000   4.820000 68.570000   8.825000 ;
      RECT 68.340000  11.040000 68.570000  15.045000 ;
      RECT 68.340000  17.260000 68.570000  21.265000 ;
      RECT 68.340000  23.480000 68.570000  27.485000 ;
      RECT 68.370000   2.835000 68.540000   4.820000 ;
      RECT 68.370000   9.055000 68.540000  11.040000 ;
      RECT 68.370000  15.275000 68.540000  17.260000 ;
      RECT 68.370000  21.495000 68.540000  23.480000 ;
      RECT 68.875000  44.755000 70.125000  45.995000 ;
      RECT 68.875000  46.185000 70.125000 198.445000 ;
      RECT 68.905000  45.995000 70.095000  46.185000 ;
      RECT 69.740000  22.520000 70.630000  28.345000 ;
      RECT 69.760000   1.890000 70.650000   2.770000 ;
      RECT 69.765000   3.845000 70.630000   8.915000 ;
      RECT 69.765000   9.845000 70.630000  14.915000 ;
      RECT 69.765000  16.165000 70.630000  21.235000 ;
      RECT 69.780000   2.770000 70.630000   3.845000 ;
      RECT 69.780000   8.915000 70.630000   9.845000 ;
      RECT 69.780000  14.915000 70.630000  16.165000 ;
      RECT 69.780000  21.235000 70.630000  22.520000 ;
      RECT 70.470000  42.820000 71.055000  42.990000 ;
      RECT 70.725000  42.735000 71.055000  42.820000 ;
      RECT 70.725000  42.990000 71.055000  43.015000 ;
      RECT 72.245000 199.210000 72.775000 199.380000 ;
      RECT 72.345000 199.380000 72.675000 199.420000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   2.170000  0.215000   2.240000 ;
      RECT  0.000000   2.170000  0.725000   2.680000 ;
      RECT  0.000000   2.240000  0.285000   2.310000 ;
      RECT  0.000000   2.310000  0.355000   2.380000 ;
      RECT  0.000000   2.380000  0.425000   2.450000 ;
      RECT  0.000000   2.450000  0.495000   2.520000 ;
      RECT  0.000000   2.520000  0.565000   2.590000 ;
      RECT  0.000000   2.590000  0.635000   2.660000 ;
      RECT  0.000000   2.660000  0.705000   2.680000 ;
      RECT  0.000000   2.680000  0.725000  36.970000 ;
      RECT  0.000000   2.680000  0.725000  36.970000 ;
      RECT  0.000000  36.970000  0.725000  37.015000 ;
      RECT  0.000000  36.970000  0.810000  37.055000 ;
      RECT  0.000000  37.015000  0.770000  37.055000 ;
      RECT  0.000000  37.055000  0.810000  46.900000 ;
      RECT  0.000000  37.055000  0.810000  46.900000 ;
      RECT  0.000000  46.900000  0.725000  46.985000 ;
      RECT  0.000000  46.900000  0.770000  46.940000 ;
      RECT  0.000000  46.940000  0.730000  46.980000 ;
      RECT  0.000000  46.980000  0.725000  46.985000 ;
      RECT  0.000000  46.985000  0.725000 195.355000 ;
      RECT  0.000000  46.985000  0.725000 195.355000 ;
      RECT  0.000000 195.355000 67.480000 200.000000 ;
      RECT  0.000000 195.355000 75.000000 200.000000 ;
      RECT 14.400000  45.430000 57.415000  47.315000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.175000 16.525000  54.100000 ;
      RECT 14.400000  47.315000 16.665000  54.100000 ;
      RECT 14.400000  54.100000 16.665000  54.905000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.445000  70.315000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.175000 24.540000  72.870000 ;
      RECT 14.400000  70.315000 24.680000  72.925000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.925000 23.590000  74.015000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.875000 18.130000  74.695000 ;
      RECT 14.400000  74.015000 18.270000  74.555000 ;
      RECT 14.400000  74.555000 24.680000  75.675000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.680000  77.125000 ;
      RECT 14.400000  75.730000 24.540000  77.125000 ;
      RECT 14.400000  77.125000 24.680000  79.295000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.505000  93.315000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.175000 24.540000 100.125000 ;
      RECT 14.400000  93.315000 24.680000 100.125000 ;
      RECT 14.400000 100.125000 24.680000 102.295000 ;
      RECT 14.400000 116.180000 24.540000 123.030000 ;
      RECT 14.400000 116.180000 57.415000 116.315000 ;
      RECT 14.400000 116.315000 24.680000 123.030000 ;
      RECT 14.400000 123.030000 24.680000 125.295000 ;
      RECT 14.400000 139.285000 16.525000 146.100000 ;
      RECT 14.400000 139.285000 57.450000 139.315000 ;
      RECT 14.400000 139.315000 16.665000 146.100000 ;
      RECT 14.400000 146.100000 16.665000 146.770000 ;
      RECT 14.400000 162.195000 16.525000 169.105000 ;
      RECT 14.400000 162.195000 57.465000 162.315000 ;
      RECT 14.400000 162.315000 16.665000 169.105000 ;
      RECT 14.400000 169.105000 16.665000 171.295000 ;
      RECT 14.400000 185.170000 15.340000 189.470000 ;
      RECT 14.400000 185.170000 15.480000 189.470000 ;
      RECT 14.400000 189.470000 15.480000 190.155000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.410000 162.185000 16.525000 162.195000 ;
      RECT 14.415000 185.155000 15.340000 185.170000 ;
      RECT 14.415000 185.155000 15.480000 185.170000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000 162.175000 16.525000 162.185000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000 139.230000 16.525000 139.285000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.470000  54.100000 16.525000  54.170000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 146.100000 16.525000 146.170000 ;
      RECT 14.470000 169.105000 16.525000 169.175000 ;
      RECT 14.470000 189.470000 15.340000 189.540000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.485000 185.085000 15.340000 185.155000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.510000 139.175000 16.525000 139.230000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.540000  54.170000 16.525000  54.240000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 146.170000 16.525000 146.240000 ;
      RECT 14.540000 169.175000 16.525000 169.245000 ;
      RECT 14.540000 189.540000 15.340000 189.610000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.555000 185.015000 15.340000 185.085000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 185.005000 58.580000 185.015000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.610000  54.240000 16.525000  54.310000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 146.240000 16.525000 146.310000 ;
      RECT 14.610000 169.245000 16.525000 169.315000 ;
      RECT 14.610000 189.610000 15.340000 189.680000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 184.935000 58.590000 185.005000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.680000  54.310000 16.525000  54.380000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 146.310000 16.525000 146.380000 ;
      RECT 14.680000 169.315000 16.525000 169.385000 ;
      RECT 14.680000 189.680000 15.340000 189.750000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 184.865000 58.660000 184.935000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.750000  54.380000 16.525000  54.450000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 146.380000 16.525000 146.450000 ;
      RECT 14.750000 169.385000 16.525000 169.455000 ;
      RECT 14.750000 189.750000 15.340000 189.820000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 184.795000 58.730000 184.865000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.820000  54.450000 16.525000  54.520000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 146.450000 16.525000 146.520000 ;
      RECT 14.820000 169.455000 16.525000 169.525000 ;
      RECT 14.820000 189.820000 15.340000 189.890000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 184.725000 58.800000 184.795000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.890000  54.520000 16.525000  54.590000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 146.520000 16.525000 146.590000 ;
      RECT 14.890000 169.525000 16.525000 169.595000 ;
      RECT 14.890000 189.890000 15.340000 189.960000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 184.655000 58.870000 184.725000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.960000  54.590000 16.525000  54.660000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 146.590000 16.525000 146.660000 ;
      RECT 14.960000 169.595000 16.525000 169.665000 ;
      RECT 14.960000 189.960000 15.340000 190.030000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 184.585000 58.940000 184.655000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.030000  54.660000 16.525000  54.730000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 146.660000 16.525000 146.730000 ;
      RECT 15.030000 169.665000 16.525000 169.735000 ;
      RECT 15.030000 190.030000 15.340000 190.100000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 184.515000 59.010000 184.585000 ;
      RECT 15.070000 146.770000 18.190000 148.295000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000 190.155000 75.000000 190.280000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.100000  54.730000 16.525000  54.800000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 146.730000 16.525000 146.800000 ;
      RECT 15.100000 169.735000 16.525000 169.805000 ;
      RECT 15.100000 190.100000 15.340000 190.170000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 146.800000 16.525000 146.825000 ;
      RECT 15.125000 184.445000 59.080000 184.515000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.170000  54.800000 16.525000  54.870000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 169.805000 16.525000 169.875000 ;
      RECT 15.170000 190.170000 15.340000 190.240000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 146.825000 16.525000 146.895000 ;
      RECT 15.195000 184.375000 59.150000 184.445000 ;
      RECT 15.205000  54.905000 18.790000  56.295000 ;
      RECT 15.210000 190.240000 15.340000 190.280000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.240000  54.870000 16.525000  54.940000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 169.875000 16.525000 169.945000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 146.895000 16.595000 146.965000 ;
      RECT 15.265000 184.305000 59.220000 184.375000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.310000  54.940000 16.525000  55.010000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 169.945000 16.525000 170.015000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 146.965000 16.665000 147.035000 ;
      RECT 15.335000 184.235000 59.290000 184.305000 ;
      RECT 15.345000  55.010000 16.525000  55.045000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 170.015000 16.525000 170.085000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 147.035000 16.735000 147.105000 ;
      RECT 15.405000 184.165000 59.360000 184.235000 ;
      RECT 15.415000  55.045000 17.345000  55.115000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 170.085000 16.525000 170.155000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 147.105000 16.805000 147.175000 ;
      RECT 15.475000 184.095000 59.430000 184.165000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 60.970000  31.015000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  31.015000 60.970000  35.550000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.070000 60.830000  35.550000 ;
      RECT 15.485000  35.550000 60.970000  35.975000 ;
      RECT 15.485000  55.115000 17.415000  55.185000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 170.155000 16.525000 170.225000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 147.175000 16.875000 147.245000 ;
      RECT 15.545000 184.025000 59.500000 184.095000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  55.185000 17.485000  55.255000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 170.225000 16.525000 170.295000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 147.245000 16.945000 147.315000 ;
      RECT 15.615000 183.955000 59.570000 184.025000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  55.255000 17.555000  55.325000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 170.295000 16.525000 170.365000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 147.315000 17.015000 147.385000 ;
      RECT 15.685000 183.885000 59.640000 183.955000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  55.325000 17.625000  55.395000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 170.365000 16.525000 170.435000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 147.385000 17.085000 147.455000 ;
      RECT 15.755000 183.815000 59.710000 183.885000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  55.395000 17.695000  55.465000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 170.435000 16.525000 170.505000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 147.455000 17.155000 147.525000 ;
      RECT 15.825000 183.745000 59.780000 183.815000 ;
      RECT 15.835000  55.465000 17.765000  55.535000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 170.505000 16.525000 170.575000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 147.525000 17.225000 147.595000 ;
      RECT 15.895000 183.675000 59.850000 183.745000 ;
      RECT 15.905000  55.535000 17.835000  55.605000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.975000 54.530000  38.195000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 170.575000 16.525000 170.645000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 147.595000 17.295000 147.665000 ;
      RECT 15.965000 183.605000 59.920000 183.675000 ;
      RECT 15.975000  55.605000 17.905000  55.675000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 170.645000 16.525000 170.715000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 147.665000 17.365000 147.735000 ;
      RECT 16.035000 183.535000 59.990000 183.605000 ;
      RECT 16.045000  55.675000 17.975000  55.745000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.070000  43.760000 59.300000  45.430000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 170.715000 16.525000 170.785000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 147.735000 17.435000 147.805000 ;
      RECT 16.105000 183.465000 60.060000 183.535000 ;
      RECT 16.115000  55.745000 18.045000  55.815000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 170.785000 16.525000 170.855000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 147.805000 17.505000 147.875000 ;
      RECT 16.175000 183.395000 60.130000 183.465000 ;
      RECT 16.185000  55.815000 18.115000  55.885000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 170.855000 16.525000 170.925000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 147.875000 17.575000 147.945000 ;
      RECT 16.245000 183.325000 60.200000 183.395000 ;
      RECT 16.255000  55.885000 18.185000  55.955000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 170.925000 16.525000 170.995000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 147.945000 17.645000 148.015000 ;
      RECT 16.315000 183.255000 60.270000 183.325000 ;
      RECT 16.325000  55.955000 18.255000  56.025000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 170.995000 16.525000 171.065000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 148.015000 17.715000 148.085000 ;
      RECT 16.385000 183.185000 60.340000 183.255000 ;
      RECT 16.395000  56.025000 18.325000  56.095000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 171.065000 16.525000 171.135000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 148.085000 17.785000 148.155000 ;
      RECT 16.455000 183.115000 60.410000 183.185000 ;
      RECT 16.465000  56.095000 18.395000  56.165000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 171.135000 16.525000 171.205000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 148.155000 17.855000 148.225000 ;
      RECT 16.525000 183.045000 60.480000 183.115000 ;
      RECT 16.535000  56.165000 18.465000  56.235000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.295000 58.700000  80.500000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.295000 58.700000 103.500000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000 171.295000 58.710000 172.500000 ;
      RECT 16.595000  56.295000 58.670000  57.500000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 148.225000 17.925000 148.295000 ;
      RECT 16.595000 148.295000 58.630000 149.500000 ;
      RECT 16.595000 182.975000 60.550000 183.045000 ;
      RECT 16.605000  56.235000 18.535000  56.305000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.665000 125.295000 58.700000 126.500000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 148.295000 17.995000 148.365000 ;
      RECT 16.665000 182.905000 60.620000 182.975000 ;
      RECT 16.675000  56.305000 18.605000  56.375000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.735000  56.375000 18.675000  56.435000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 148.365000 18.065000 148.435000 ;
      RECT 16.735000 182.835000 60.690000 182.905000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000 182.820000 58.635000 185.155000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 57.440000  79.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 57.440000 102.505000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000 171.435000 57.450000 171.505000 ;
      RECT 16.805000  56.435000 57.410000  56.505000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 148.435000 57.370000 148.505000 ;
      RECT 16.805000 182.765000 60.760000 182.835000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.830000 182.740000 60.830000 182.765000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 57.510000  79.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 57.510000 102.575000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000 171.505000 57.520000 171.575000 ;
      RECT 16.875000  56.505000 57.480000  56.575000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 57.440000 125.505000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 148.505000 57.440000 148.575000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.900000 182.670000 60.830000 182.740000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 57.580000  79.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 57.580000 102.645000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000 171.575000 57.590000 171.645000 ;
      RECT 16.945000  56.575000 57.550000  56.645000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 57.510000 125.575000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 148.575000 57.510000 148.645000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.970000 182.600000 60.830000 182.670000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 57.650000  79.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 57.650000 102.715000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000 171.645000 57.660000 171.715000 ;
      RECT 17.015000  56.645000 57.620000  56.715000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 57.580000 125.645000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 148.645000 57.580000 148.715000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.040000 182.530000 60.830000 182.600000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 57.720000  79.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 57.720000 102.785000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000 171.715000 57.730000 171.785000 ;
      RECT 17.085000  56.715000 57.690000  56.785000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 57.650000 125.715000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 148.715000 57.650000 148.785000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.110000 182.460000 60.830000 182.530000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 57.790000  79.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 57.790000 102.855000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000 171.785000 57.800000 171.855000 ;
      RECT 17.155000  56.785000 57.760000  56.855000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 57.720000 125.785000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 148.785000 57.720000 148.855000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.970000  43.760000 ;
      RECT 17.180000 182.390000 60.830000 182.460000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 57.860000  79.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 57.860000 102.925000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000 171.855000 57.870000 171.925000 ;
      RECT 17.225000  56.855000 57.830000  56.925000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 57.790000 125.855000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 148.855000 57.790000 148.925000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.250000 182.320000 60.830000 182.390000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 57.930000  79.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 57.930000 102.995000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000 171.925000 57.940000 171.995000 ;
      RECT 17.295000  56.925000 57.900000  56.995000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 57.860000 125.925000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 148.925000 57.860000 148.995000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.320000 182.250000 60.830000 182.320000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 58.000000  80.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 58.000000 103.065000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000 171.995000 58.010000 172.065000 ;
      RECT 17.365000  56.995000 57.970000  57.065000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 57.930000 125.995000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 148.995000 57.930000 149.065000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.390000 182.180000 60.830000 182.250000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 58.070000  80.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 58.070000 103.135000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000 172.065000 58.080000 172.135000 ;
      RECT 17.435000  57.065000 58.040000  57.135000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 58.000000 126.065000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 149.065000 58.000000 149.135000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.460000 182.110000 60.830000 182.180000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 58.140000  80.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 58.140000 103.205000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000 172.135000 58.150000 172.205000 ;
      RECT 17.505000  57.135000 58.110000  57.205000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 58.070000 126.135000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 149.135000 58.070000 149.205000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.530000 182.040000 60.830000 182.110000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 58.210000  80.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 58.210000 103.275000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000 172.205000 58.220000 172.275000 ;
      RECT 17.575000  57.205000 58.180000  57.275000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 58.140000 126.205000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 149.205000 58.140000 149.275000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.600000 181.970000 60.830000 182.040000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 58.280000  80.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 58.280000 103.345000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000 172.275000 58.290000 172.345000 ;
      RECT 17.645000  57.275000 58.250000  57.345000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 58.210000 126.275000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 149.275000 58.210000 149.345000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.670000 181.900000 60.830000 181.970000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 58.350000  80.415000 ;
      RECT 17.690000  89.850000 57.680000  93.140000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 58.350000 103.415000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000 172.345000 58.360000 172.415000 ;
      RECT 17.715000  57.345000 58.320000  57.415000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 58.280000 126.345000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 149.345000 58.280000 149.415000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.740000 181.830000 60.830000 181.900000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.750000  66.790000 57.620000  70.140000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 58.420000  80.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 58.420000 103.485000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 58.490000  80.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 58.490000 103.500000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.970000  66.790000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.970000  89.850000 ;
      RECT 17.780000 172.415000 58.430000 172.485000 ;
      RECT 17.785000  57.415000 58.390000  57.485000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 58.350000 126.415000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 149.415000 58.350000 149.485000 ;
      RECT 17.785000 158.810000 57.585000 162.195000 ;
      RECT 17.795000 172.485000 58.500000 172.500000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  57.485000 58.460000  57.500000 ;
      RECT 17.800000 149.485000 58.420000 149.500000 ;
      RECT 17.810000 181.760000 60.830000 181.830000 ;
      RECT 17.810000 181.760000 60.970000 182.820000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.820000 112.760000 57.550000 116.180000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.821000 112.760000 60.970000 112.762000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.970000 158.810000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 58.420000 126.485000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 58.490000 126.500000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.890000 135.795000 57.480000 139.285000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.970000 135.795000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.135000  38.195000 52.655000  40.070000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 59.390000  29.430000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.400000  40.070000 52.515000  40.210000 ;
      RECT 22.850000  42.520000 60.970000  42.660000 ;
      RECT 24.675000   0.000000 25.615000   0.815000 ;
      RECT 24.675000   0.000000 25.755000   0.675000 ;
      RECT 24.675000   0.675000 50.250000   8.480000 ;
      RECT 24.675000   0.815000 50.110000   8.480000 ;
      RECT 24.675000   8.480000 50.250000   8.565000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.765000   8.565000 46.695000  12.120000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 28.035000   0.000000 50.250000   0.675000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.175000   0.000000 50.110000   0.815000 ;
      RECT 28.175000   0.000000 50.110000   8.480000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 37.175000  12.120000 37.610000  25.940000 ;
      RECT 37.175000  12.120000 46.660000  12.155000 ;
      RECT 37.175000  12.155000 37.750000  25.800000 ;
      RECT 37.175000  25.800000 55.935000  25.980000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 60.970000  82.770000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.770000 60.970000  89.760000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.825000 60.830000  89.760000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 60.970000 105.770000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.770000 60.970000 112.760000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.825000 60.830000 112.705000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 60.970000 128.770000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.770000 60.970000 135.760000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.825000 60.830000 135.740000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 60.970000 151.840000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.840000 60.970000 158.760000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.895000 60.830000 158.755000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 60.970000  59.800000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.800000 60.970000  66.760000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.855000 60.830000  66.735000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 57.055000  35.975000 60.970000  39.725000 ;
      RECT 57.055000  39.725000 60.970000  42.520000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.195000  35.835000 60.830000  39.780000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 58.240000 172.500000 58.515000 172.570000 ;
      RECT 58.240000 172.500000 60.970000 174.760000 ;
      RECT 58.240000 172.570000 58.585000 172.640000 ;
      RECT 58.240000 172.640000 58.655000 172.710000 ;
      RECT 58.240000 172.710000 58.725000 172.780000 ;
      RECT 58.240000 172.780000 58.795000 172.850000 ;
      RECT 58.240000 172.850000 58.865000 172.920000 ;
      RECT 58.240000 172.920000 58.935000 172.990000 ;
      RECT 58.240000 172.990000 59.005000 173.060000 ;
      RECT 58.240000 173.060000 59.075000 173.130000 ;
      RECT 58.240000 173.130000 59.145000 173.200000 ;
      RECT 58.240000 173.200000 59.215000 173.270000 ;
      RECT 58.240000 173.270000 59.285000 173.340000 ;
      RECT 58.240000 173.340000 59.355000 173.410000 ;
      RECT 58.240000 173.410000 59.425000 173.480000 ;
      RECT 58.240000 173.480000 59.495000 173.550000 ;
      RECT 58.240000 173.550000 59.565000 173.620000 ;
      RECT 58.240000 173.620000 59.635000 173.690000 ;
      RECT 58.240000 173.690000 59.705000 173.760000 ;
      RECT 58.240000 173.760000 59.775000 173.830000 ;
      RECT 58.240000 173.830000 59.845000 173.900000 ;
      RECT 58.240000 173.900000 59.915000 173.970000 ;
      RECT 58.240000 173.970000 59.985000 174.040000 ;
      RECT 58.240000 174.040000 60.055000 174.110000 ;
      RECT 58.240000 174.110000 60.125000 174.180000 ;
      RECT 58.240000 174.180000 60.195000 174.250000 ;
      RECT 58.240000 174.250000 60.265000 174.320000 ;
      RECT 58.240000 174.320000 60.335000 174.390000 ;
      RECT 58.240000 174.390000 60.405000 174.460000 ;
      RECT 58.240000 174.460000 60.475000 174.530000 ;
      RECT 58.240000 174.530000 60.545000 174.600000 ;
      RECT 58.240000 174.600000 60.615000 174.670000 ;
      RECT 58.240000 174.670000 60.685000 174.740000 ;
      RECT 58.240000 174.740000 60.755000 174.810000 ;
      RECT 58.240000 174.760000 60.970000 181.760000 ;
      RECT 58.240000 174.810000 60.825000 174.815000 ;
      RECT 58.240000 174.815000 60.830000 181.760000 ;
      RECT 67.480000 190.280000 75.000000 195.355000 ;
      RECT 67.480000 190.295000 75.000000 200.000000 ;
      RECT 70.480000 193.295000 72.000000 197.000000 ;
      RECT 74.430000   0.000000 75.000000 190.155000 ;
      RECT 74.570000   0.000000 75.000000 190.295000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.195000  36.635000 ;
      RECT  0.000000  36.635000  0.810000  37.250000 ;
      RECT  0.000000  36.730000  0.150000  36.880000 ;
      RECT  0.000000  36.880000  0.300000  37.030000 ;
      RECT  0.000000  37.030000  0.450000  37.180000 ;
      RECT  0.000000  37.180000  0.600000  37.290000 ;
      RECT  0.000000  37.250000  0.810000  46.220000 ;
      RECT  0.000000  37.290000  0.710000  46.180000 ;
      RECT  0.000000  46.180000  0.560000  46.330000 ;
      RECT  0.000000  46.220000  0.195000  46.835000 ;
      RECT  0.000000  46.330000  0.410000  46.480000 ;
      RECT  0.000000  46.480000  0.260000  46.630000 ;
      RECT  0.000000  46.630000  0.110000  46.780000 ;
      RECT  0.000000  46.835000  0.195000 173.455000 ;
      RECT  0.000000 173.455000  2.760000 185.195000 ;
      RECT  0.000000 173.555000 14.250000 173.705000 ;
      RECT  0.000000 173.705000 14.100000 173.855000 ;
      RECT  0.000000 173.855000 13.950000 174.005000 ;
      RECT  0.000000 174.005000 13.800000 174.155000 ;
      RECT  0.000000 174.155000 13.650000 174.305000 ;
      RECT  0.000000 174.305000 13.500000 174.455000 ;
      RECT  0.000000 174.455000 13.350000 174.605000 ;
      RECT  0.000000 174.605000 13.200000 174.755000 ;
      RECT  0.000000 174.755000 13.050000 174.905000 ;
      RECT  0.000000 174.905000 12.900000 175.055000 ;
      RECT  0.000000 175.055000 12.750000 175.205000 ;
      RECT  0.000000 175.205000 12.600000 175.355000 ;
      RECT  0.000000 175.355000 12.450000 175.505000 ;
      RECT  0.000000 175.505000 12.300000 175.655000 ;
      RECT  0.000000 175.655000 12.150000 175.805000 ;
      RECT  0.000000 175.805000 12.000000 175.955000 ;
      RECT  0.000000 175.955000 11.850000 176.105000 ;
      RECT  0.000000 176.105000 11.700000 176.255000 ;
      RECT  0.000000 176.255000 11.550000 176.405000 ;
      RECT  0.000000 176.405000 11.400000 176.555000 ;
      RECT  0.000000 176.555000 11.250000 176.705000 ;
      RECT  0.000000 176.705000 11.100000 176.855000 ;
      RECT  0.000000 176.855000 10.950000 177.005000 ;
      RECT  0.000000 177.005000 10.800000 177.155000 ;
      RECT  0.000000 177.155000 10.650000 177.305000 ;
      RECT  0.000000 177.305000 10.500000 177.455000 ;
      RECT  0.000000 177.455000 10.350000 177.605000 ;
      RECT  0.000000 177.605000 10.200000 177.755000 ;
      RECT  0.000000 177.755000 10.050000 177.905000 ;
      RECT  0.000000 177.905000  9.900000 178.055000 ;
      RECT  0.000000 178.055000  9.750000 178.205000 ;
      RECT  0.000000 178.205000  9.600000 178.355000 ;
      RECT  0.000000 178.355000  9.450000 178.505000 ;
      RECT  0.000000 178.505000  9.300000 178.655000 ;
      RECT  0.000000 178.655000  9.150000 178.805000 ;
      RECT  0.000000 178.805000  9.000000 178.955000 ;
      RECT  0.000000 178.955000  8.850000 179.105000 ;
      RECT  0.000000 179.105000  8.700000 179.255000 ;
      RECT  0.000000 179.255000  8.550000 179.405000 ;
      RECT  0.000000 179.405000  8.400000 179.555000 ;
      RECT  0.000000 179.555000  8.250000 179.705000 ;
      RECT  0.000000 179.705000  8.100000 179.855000 ;
      RECT  0.000000 179.855000  7.950000 180.005000 ;
      RECT  0.000000 180.005000  7.800000 180.155000 ;
      RECT  0.000000 180.155000  7.650000 180.305000 ;
      RECT  0.000000 180.305000  7.500000 180.455000 ;
      RECT  0.000000 180.455000  7.350000 180.605000 ;
      RECT  0.000000 180.605000  7.200000 180.755000 ;
      RECT  0.000000 180.755000  7.050000 180.905000 ;
      RECT  0.000000 180.905000  6.900000 181.055000 ;
      RECT  0.000000 181.055000  6.750000 181.205000 ;
      RECT  0.000000 181.205000  6.600000 181.355000 ;
      RECT  0.000000 181.355000  6.450000 181.505000 ;
      RECT  0.000000 181.505000  6.300000 181.655000 ;
      RECT  0.000000 181.655000  6.150000 181.805000 ;
      RECT  0.000000 181.805000  6.000000 181.955000 ;
      RECT  0.000000 181.955000  5.850000 182.105000 ;
      RECT  0.000000 182.105000  5.700000 182.255000 ;
      RECT  0.000000 182.255000  5.550000 182.405000 ;
      RECT  0.000000 182.405000  5.400000 182.555000 ;
      RECT  0.000000 182.555000  5.250000 182.705000 ;
      RECT  0.000000 182.705000  5.100000 182.855000 ;
      RECT  0.000000 182.855000  4.950000 183.005000 ;
      RECT  0.000000 183.005000  4.800000 183.155000 ;
      RECT  0.000000 183.155000  4.650000 183.305000 ;
      RECT  0.000000 183.305000  4.500000 183.455000 ;
      RECT  0.000000 183.455000  4.350000 183.605000 ;
      RECT  0.000000 183.605000  4.200000 183.755000 ;
      RECT  0.000000 183.755000  4.050000 183.905000 ;
      RECT  0.000000 183.905000  3.900000 184.055000 ;
      RECT  0.000000 184.055000  3.750000 184.205000 ;
      RECT  0.000000 184.205000  3.600000 184.355000 ;
      RECT  0.000000 184.355000  3.450000 184.505000 ;
      RECT  0.000000 184.505000  3.300000 184.655000 ;
      RECT  0.000000 184.655000  3.150000 184.805000 ;
      RECT  0.000000 184.805000  3.000000 184.955000 ;
      RECT  0.000000 184.955000  2.850000 185.105000 ;
      RECT  0.000000 185.105000  2.760000 185.195000 ;
      RECT  0.000000 185.195000  2.760000 200.000000 ;
      RECT  0.000000 185.195000  2.760000 200.000000 ;
      RECT  3.000000 176.555000  7.005000 176.705000 ;
      RECT  3.000000 176.555000  7.005000 176.705000 ;
      RECT  3.000000 176.705000  6.855000 176.855000 ;
      RECT  3.000000 176.705000  6.855000 176.855000 ;
      RECT  3.000000 176.855000  6.705000 177.005000 ;
      RECT  3.000000 176.855000  6.705000 177.005000 ;
      RECT  3.000000 177.005000  6.555000 177.155000 ;
      RECT  3.000000 177.005000  6.555000 177.155000 ;
      RECT  3.000000 177.155000  6.405000 177.305000 ;
      RECT  3.000000 177.155000  6.405000 177.305000 ;
      RECT  3.000000 177.305000  6.255000 177.455000 ;
      RECT  3.000000 177.305000  6.255000 177.455000 ;
      RECT  3.000000 177.455000  6.105000 177.605000 ;
      RECT  3.000000 177.455000  6.105000 177.605000 ;
      RECT  3.000000 177.605000  5.955000 177.755000 ;
      RECT  3.000000 177.605000  5.955000 177.755000 ;
      RECT  3.000000 177.755000  5.805000 177.905000 ;
      RECT  3.000000 177.755000  5.805000 177.905000 ;
      RECT  3.000000 177.905000  5.655000 178.055000 ;
      RECT  3.000000 177.905000  5.655000 178.055000 ;
      RECT  3.000000 178.055000  5.505000 178.205000 ;
      RECT  3.000000 178.055000  5.505000 178.205000 ;
      RECT  3.000000 178.205000  5.355000 178.355000 ;
      RECT  3.000000 178.205000  5.355000 178.355000 ;
      RECT  3.000000 178.355000  5.205000 178.505000 ;
      RECT  3.000000 178.355000  5.205000 178.505000 ;
      RECT  3.000000 178.505000  5.055000 178.655000 ;
      RECT  3.000000 178.505000  5.055000 178.655000 ;
      RECT  3.000000 178.655000  4.905000 178.805000 ;
      RECT  3.000000 178.655000  4.905000 178.805000 ;
      RECT  3.000000 178.805000  4.755000 178.955000 ;
      RECT  3.000000 178.805000  4.755000 178.955000 ;
      RECT  3.000000 178.955000  4.605000 179.105000 ;
      RECT  3.000000 178.955000  4.605000 179.105000 ;
      RECT  3.000000 179.105000  4.455000 179.255000 ;
      RECT  3.000000 179.105000  4.455000 179.255000 ;
      RECT  3.000000 179.255000  4.305000 179.405000 ;
      RECT  3.000000 179.255000  4.305000 179.405000 ;
      RECT  3.000000 179.405000  4.155000 179.555000 ;
      RECT  3.000000 179.405000  4.155000 179.555000 ;
      RECT  3.000000 179.555000  4.005000 179.705000 ;
      RECT  3.000000 179.555000  4.005000 179.705000 ;
      RECT  3.000000 179.705000  3.855000 179.855000 ;
      RECT  3.000000 179.705000  3.855000 179.855000 ;
      RECT  3.000000 179.855000  3.705000 180.005000 ;
      RECT  3.000000 179.855000  3.705000 180.005000 ;
      RECT  3.000000 180.005000  3.555000 180.155000 ;
      RECT  3.000000 180.005000  3.555000 180.155000 ;
      RECT  3.000000 180.155000  3.405000 180.305000 ;
      RECT  3.000000 180.155000  3.405000 180.305000 ;
      RECT  3.000000 180.305000  3.255000 180.455000 ;
      RECT  3.000000 180.305000  3.255000 180.455000 ;
      RECT  3.000000 180.455000  3.105000 180.605000 ;
      RECT  3.000000 180.455000  3.105000 180.605000 ;
      RECT  3.000000 180.605000  3.005000 180.705000 ;
      RECT  3.000000 180.605000  3.005000 180.705000 ;
      RECT 13.800000 101.520000 15.100000 102.035000 ;
      RECT 13.800000 102.035000 15.100000 172.855000 ;
      RECT 13.800000 172.855000 14.500000 173.455000 ;
      RECT 13.900000 101.560000 15.425000 101.710000 ;
      RECT 13.900000 101.710000 15.275000 101.860000 ;
      RECT 13.900000 101.860000 15.125000 102.010000 ;
      RECT 13.900000 102.010000 15.100000 102.035000 ;
      RECT 13.900000 102.035000 15.100000 172.855000 ;
      RECT 13.900000 172.855000 14.950000 173.005000 ;
      RECT 13.900000 173.005000 14.800000 173.155000 ;
      RECT 13.900000 173.155000 14.650000 173.305000 ;
      RECT 13.900000 173.305000 14.500000 173.455000 ;
      RECT 13.900000 173.455000 14.400000 173.555000 ;
      RECT 14.020000 101.440000 15.575000 101.560000 ;
      RECT 14.170000 101.290000 15.695000 101.440000 ;
      RECT 14.320000 101.140000 15.845000 101.290000 ;
      RECT 14.470000 100.990000 15.995000 101.140000 ;
      RECT 14.620000 100.840000 16.145000 100.990000 ;
      RECT 14.770000 100.690000 16.295000 100.840000 ;
      RECT 14.920000 100.540000 16.445000 100.690000 ;
      RECT 15.070000 100.390000 16.595000 100.540000 ;
      RECT 15.220000 100.240000 16.745000 100.390000 ;
      RECT 15.370000 100.090000 16.895000 100.240000 ;
      RECT 15.520000  99.940000 17.045000 100.090000 ;
      RECT 15.670000  99.790000 17.195000  99.940000 ;
      RECT 15.820000  99.640000 17.345000  99.790000 ;
      RECT 15.970000  99.490000 17.495000  99.640000 ;
      RECT 16.120000  99.340000 17.645000  99.490000 ;
      RECT 16.270000  99.190000 17.795000  99.340000 ;
      RECT 16.420000  99.040000 17.945000  99.190000 ;
      RECT 16.570000  98.890000 18.095000  99.040000 ;
      RECT 16.720000  98.740000 18.245000  98.890000 ;
      RECT 16.870000  98.590000 18.395000  98.740000 ;
      RECT 17.020000  98.440000 18.545000  98.590000 ;
      RECT 17.170000  98.290000 18.695000  98.440000 ;
      RECT 17.320000  98.140000 18.845000  98.290000 ;
      RECT 17.470000  97.990000 18.995000  98.140000 ;
      RECT 17.620000  97.840000 19.145000  97.990000 ;
      RECT 17.770000  97.690000 19.295000  97.840000 ;
      RECT 17.920000  97.540000 19.445000  97.690000 ;
      RECT 18.070000  97.390000 19.595000  97.540000 ;
      RECT 18.220000  97.240000 19.745000  97.390000 ;
      RECT 18.370000  97.090000 19.895000  97.240000 ;
      RECT 18.520000  96.940000 20.045000  97.090000 ;
      RECT 18.670000  96.790000 20.195000  96.940000 ;
      RECT 18.820000  96.640000 20.345000  96.790000 ;
      RECT 18.970000  96.490000 20.495000  96.640000 ;
      RECT 19.120000  96.340000 20.645000  96.490000 ;
      RECT 19.270000  96.190000 20.795000  96.340000 ;
      RECT 19.420000  96.040000 20.945000  96.190000 ;
      RECT 19.570000  95.890000 21.095000  96.040000 ;
      RECT 19.720000  95.740000 21.245000  95.890000 ;
      RECT 19.870000  95.590000 21.395000  95.740000 ;
      RECT 20.020000  95.440000 21.545000  95.590000 ;
      RECT 20.170000  95.290000 21.695000  95.440000 ;
      RECT 20.320000  95.140000 21.845000  95.290000 ;
      RECT 20.470000  94.990000 21.995000  95.140000 ;
      RECT 20.620000  94.840000 22.145000  94.990000 ;
      RECT 20.770000  94.690000 22.295000  94.840000 ;
      RECT 20.920000  94.540000 22.445000  94.690000 ;
      RECT 21.070000  94.390000 22.595000  94.540000 ;
      RECT 21.220000  94.240000 22.745000  94.390000 ;
      RECT 21.370000  94.090000 22.895000  94.240000 ;
      RECT 21.520000  93.940000 23.045000  94.090000 ;
      RECT 21.670000  93.790000 23.195000  93.940000 ;
      RECT 21.695000  93.765000 23.345000  93.790000 ;
      RECT 21.845000  93.615000 23.345000  93.765000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 168.965000 25.530000 172.475000 ;
      RECT 21.970000 104.775000 25.530000 104.845000 ;
      RECT 21.995000  93.465000 23.345000  93.615000 ;
      RECT 22.050000 168.965000 25.530000 169.115000 ;
      RECT 22.120000 104.625000 25.530000 104.775000 ;
      RECT 22.145000  93.315000 23.345000  93.465000 ;
      RECT 22.200000 169.115000 25.530000 169.265000 ;
      RECT 22.270000 104.475000 25.530000 104.625000 ;
      RECT 22.295000  93.165000 23.345000  93.315000 ;
      RECT 22.350000 169.265000 25.530000 169.415000 ;
      RECT 22.420000 104.325000 25.530000 104.475000 ;
      RECT 22.445000  93.015000 23.345000  93.165000 ;
      RECT 22.500000 169.415000 25.530000 169.565000 ;
      RECT 22.570000 104.175000 25.530000 104.325000 ;
      RECT 22.595000  92.865000 23.345000  93.015000 ;
      RECT 22.650000 169.565000 25.530000 169.715000 ;
      RECT 22.720000 104.025000 25.530000 104.175000 ;
      RECT 22.745000  92.715000 23.345000  92.865000 ;
      RECT 22.800000 169.715000 25.530000 169.865000 ;
      RECT 22.870000 103.875000 25.530000 104.025000 ;
      RECT 22.895000  92.565000 23.345000  92.715000 ;
      RECT 22.945000  92.375000 23.345000  93.790000 ;
      RECT 22.950000 169.865000 25.530000 170.015000 ;
      RECT 23.020000 103.725000 25.530000 103.875000 ;
      RECT 23.045000  92.415000 23.345000  92.565000 ;
      RECT 23.100000 170.015000 25.530000 170.165000 ;
      RECT 23.170000 103.575000 25.530000 103.725000 ;
      RECT 23.195000  92.265000 23.345000  92.415000 ;
      RECT 23.250000 170.165000 25.530000 170.315000 ;
      RECT 23.320000 103.425000 25.530000 103.575000 ;
      RECT 23.400000 170.315000 25.530000 170.465000 ;
      RECT 23.470000 103.275000 25.530000 103.425000 ;
      RECT 23.550000 170.465000 25.530000 170.615000 ;
      RECT 23.620000 103.125000 25.530000 103.275000 ;
      RECT 23.700000 170.615000 25.530000 170.765000 ;
      RECT 23.770000 102.975000 25.530000 103.125000 ;
      RECT 23.850000 170.765000 25.530000 170.915000 ;
      RECT 23.920000 102.825000 25.530000 102.975000 ;
      RECT 24.000000 170.915000 25.530000 171.065000 ;
      RECT 24.070000 102.675000 25.530000 102.825000 ;
      RECT 24.150000 171.065000 25.530000 171.215000 ;
      RECT 24.220000 102.525000 25.530000 102.675000 ;
      RECT 24.300000 171.215000 25.530000 171.365000 ;
      RECT 24.370000 102.375000 25.530000 102.525000 ;
      RECT 24.450000 171.365000 25.530000 171.515000 ;
      RECT 24.520000 102.225000 25.530000 102.375000 ;
      RECT 24.520000 102.225000 25.530000 104.845000 ;
      RECT 24.525000 102.220000 25.530000 102.225000 ;
      RECT 24.600000 171.515000 25.530000 171.665000 ;
      RECT 24.675000 102.070000 25.535000 102.220000 ;
      RECT 24.695000   0.000000 25.495000  90.225000 ;
      RECT 24.695000  90.225000 25.095000  90.625000 ;
      RECT 24.750000 171.665000 25.530000 171.815000 ;
      RECT 24.795000   0.000000 25.495000  90.225000 ;
      RECT 24.795000  90.225000 25.345000  90.375000 ;
      RECT 24.795000  90.375000 25.195000  90.525000 ;
      RECT 24.795000  90.525000 25.045000  90.675000 ;
      RECT 24.795000  90.675000 24.895000  90.825000 ;
      RECT 24.825000 101.920000 25.685000 102.070000 ;
      RECT 24.900000 171.815000 25.530000 171.965000 ;
      RECT 24.975000 101.770000 25.835000 101.920000 ;
      RECT 25.050000 171.965000 25.530000 172.115000 ;
      RECT 25.125000 101.620000 25.985000 101.770000 ;
      RECT 25.200000 172.115000 25.530000 172.265000 ;
      RECT 25.275000 101.470000 26.135000 101.620000 ;
      RECT 25.350000 172.265000 25.530000 172.415000 ;
      RECT 25.410000 172.475000 25.530000 200.000000 ;
      RECT 25.425000 101.320000 26.285000 101.470000 ;
      RECT 25.500000 172.415000 25.530000 172.565000 ;
      RECT 25.575000 101.170000 26.435000 101.320000 ;
      RECT 25.725000 101.020000 26.585000 101.170000 ;
      RECT 25.875000 100.870000 26.735000 101.020000 ;
      RECT 26.025000 100.720000 26.885000 100.870000 ;
      RECT 26.175000 100.570000 27.035000 100.720000 ;
      RECT 26.325000 100.420000 27.185000 100.570000 ;
      RECT 26.475000 100.270000 27.335000 100.420000 ;
      RECT 26.625000 100.120000 27.485000 100.270000 ;
      RECT 26.775000  99.970000 27.635000 100.120000 ;
      RECT 26.925000  99.820000 27.785000  99.970000 ;
      RECT 27.075000  99.670000 27.935000  99.820000 ;
      RECT 27.225000  99.520000 28.085000  99.670000 ;
      RECT 27.375000  99.370000 28.235000  99.520000 ;
      RECT 27.525000  99.220000 28.385000  99.370000 ;
      RECT 27.675000  99.070000 28.535000  99.220000 ;
      RECT 27.825000  98.920000 28.685000  99.070000 ;
      RECT 27.975000  98.770000 28.835000  98.920000 ;
      RECT 28.125000  98.620000 28.985000  98.770000 ;
      RECT 28.275000  98.470000 29.135000  98.620000 ;
      RECT 28.425000  98.320000 29.285000  98.470000 ;
      RECT 28.575000  98.170000 29.435000  98.320000 ;
      RECT 28.725000  98.020000 29.585000  98.170000 ;
      RECT 28.875000  97.870000 29.735000  98.020000 ;
      RECT 29.025000  97.720000 29.885000  97.870000 ;
      RECT 29.175000  97.570000 30.035000  97.720000 ;
      RECT 29.325000  97.420000 30.185000  97.570000 ;
      RECT 29.475000  97.270000 30.335000  97.420000 ;
      RECT 29.625000  97.120000 30.485000  97.270000 ;
      RECT 29.775000  96.970000 30.635000  97.120000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  96.210000 30.935000  96.820000 ;
      RECT 29.925000  96.210000 31.395000  96.360000 ;
      RECT 29.925000  96.360000 31.245000  96.510000 ;
      RECT 29.925000  96.510000 31.095000  96.660000 ;
      RECT 29.925000  96.660000 30.945000  96.810000 ;
      RECT 29.925000  96.810000 30.935000  96.820000 ;
      RECT 29.925000  96.820000 30.785000  96.970000 ;
      RECT 29.950000  93.240000 31.520000  93.265000 ;
      RECT 30.100000  93.090000 31.370000  93.240000 ;
      RECT 30.250000  92.940000 31.220000  93.090000 ;
      RECT 30.400000  92.790000 31.070000  92.940000 ;
      RECT 30.400000  92.790000 31.545000  93.265000 ;
      RECT 32.330000  99.865000 37.490000 110.785000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 42.455000 110.785000 ;
      RECT 32.330000 105.820000 42.455000 175.185000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 170.295000 37.565000 175.185000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.220000 175.185000 37.565000 190.420000 ;
      RECT 37.220000 175.270000 37.305000 175.355000 ;
      RECT 37.220000 175.355000 37.565000 190.420000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.295000   0.000000 37.490000 100.060000 ;
      RECT 37.295000 100.060000 37.490000 105.025000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.480000 175.270000 37.565000 175.355000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 101.970000 44.860000 102.580000 ;
      RECT 43.265000 100.355000 44.835000 100.380000 ;
      RECT 43.390000 101.970000 44.860000 102.120000 ;
      RECT 43.415000 100.205000 44.685000 100.355000 ;
      RECT 43.540000 102.120000 44.860000 102.270000 ;
      RECT 43.565000 100.055000 44.535000 100.205000 ;
      RECT 43.690000 102.270000 44.860000 102.420000 ;
      RECT 43.715000  99.905000 44.385000 100.055000 ;
      RECT 43.715000  99.905000 44.860000 100.380000 ;
      RECT 43.840000 102.420000 44.860000 102.570000 ;
      RECT 43.850000 102.570000 44.860000 102.580000 ;
      RECT 43.850000 102.580000 50.265000 107.985000 ;
      RECT 44.000000 102.580000 44.860000 102.730000 ;
      RECT 44.150000 102.730000 45.010000 102.880000 ;
      RECT 44.300000 102.880000 45.160000 103.030000 ;
      RECT 44.450000 103.030000 45.310000 103.180000 ;
      RECT 44.600000 103.180000 45.460000 103.330000 ;
      RECT 44.750000 103.330000 45.610000 103.480000 ;
      RECT 44.900000 103.480000 45.760000 103.630000 ;
      RECT 45.050000 103.630000 45.910000 103.780000 ;
      RECT 45.200000 103.780000 46.060000 103.930000 ;
      RECT 45.350000 103.930000 46.210000 104.080000 ;
      RECT 45.500000 104.080000 46.360000 104.230000 ;
      RECT 45.650000 104.230000 46.510000 104.380000 ;
      RECT 45.800000 104.380000 46.660000 104.530000 ;
      RECT 45.950000 104.530000 46.810000 104.680000 ;
      RECT 46.100000 104.680000 46.960000 104.830000 ;
      RECT 46.250000 104.830000 47.110000 104.980000 ;
      RECT 46.400000 104.980000 47.260000 105.130000 ;
      RECT 46.550000 105.130000 47.410000 105.280000 ;
      RECT 46.700000 105.280000 47.560000 105.430000 ;
      RECT 46.850000 105.430000 47.710000 105.580000 ;
      RECT 47.000000 105.580000 47.860000 105.730000 ;
      RECT 47.150000 105.730000 48.010000 105.880000 ;
      RECT 47.300000 105.880000 48.160000 106.030000 ;
      RECT 47.450000 106.030000 48.310000 106.180000 ;
      RECT 47.600000 106.180000 48.460000 106.330000 ;
      RECT 47.750000 106.330000 48.610000 106.480000 ;
      RECT 47.900000 106.480000 48.760000 106.630000 ;
      RECT 48.050000 106.630000 48.910000 106.780000 ;
      RECT 48.200000 106.780000 49.060000 106.930000 ;
      RECT 48.350000 106.930000 49.210000 107.080000 ;
      RECT 48.500000 107.080000 49.360000 107.230000 ;
      RECT 48.650000 107.230000 49.510000 107.380000 ;
      RECT 48.800000 107.380000 49.660000 107.530000 ;
      RECT 48.950000 107.530000 49.810000 107.680000 ;
      RECT 49.100000 107.680000 49.960000 107.830000 ;
      RECT 49.250000 107.830000 50.110000 107.980000 ;
      RECT 49.255000 107.980000 50.260000 107.985000 ;
      RECT 49.255000 107.985000 50.265000 108.135000 ;
      RECT 49.255000 107.985000 52.885000 110.605000 ;
      RECT 49.255000 108.135000 50.415000 108.285000 ;
      RECT 49.255000 108.285000 50.565000 108.435000 ;
      RECT 49.255000 108.435000 50.715000 108.585000 ;
      RECT 49.255000 108.585000 50.865000 108.735000 ;
      RECT 49.255000 108.735000 51.015000 108.885000 ;
      RECT 49.255000 108.885000 51.165000 109.035000 ;
      RECT 49.255000 109.035000 51.315000 109.185000 ;
      RECT 49.255000 109.185000 51.465000 109.335000 ;
      RECT 49.255000 109.335000 51.615000 109.485000 ;
      RECT 49.255000 109.485000 51.765000 109.635000 ;
      RECT 49.255000 109.635000 51.915000 109.785000 ;
      RECT 49.255000 109.785000 52.065000 109.935000 ;
      RECT 49.255000 109.935000 52.215000 110.085000 ;
      RECT 49.255000 110.085000 52.365000 110.235000 ;
      RECT 49.255000 110.235000 52.515000 110.385000 ;
      RECT 49.255000 110.385000 52.665000 110.535000 ;
      RECT 49.255000 110.535000 52.815000 110.605000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 168.970000 49.375000 172.480000 ;
      RECT 49.255000 168.970000 52.735000 169.120000 ;
      RECT 49.255000 169.120000 52.585000 169.270000 ;
      RECT 49.255000 169.270000 52.435000 169.420000 ;
      RECT 49.255000 169.420000 52.285000 169.570000 ;
      RECT 49.255000 169.570000 52.135000 169.720000 ;
      RECT 49.255000 169.720000 51.985000 169.870000 ;
      RECT 49.255000 169.870000 51.835000 170.020000 ;
      RECT 49.255000 170.020000 51.685000 170.170000 ;
      RECT 49.255000 170.170000 51.535000 170.320000 ;
      RECT 49.255000 170.320000 51.385000 170.470000 ;
      RECT 49.255000 170.470000 51.235000 170.620000 ;
      RECT 49.255000 170.620000 51.085000 170.770000 ;
      RECT 49.255000 170.770000 50.935000 170.920000 ;
      RECT 49.255000 170.920000 50.785000 171.070000 ;
      RECT 49.255000 171.070000 50.635000 171.220000 ;
      RECT 49.255000 171.220000 50.485000 171.370000 ;
      RECT 49.255000 171.370000 50.335000 171.520000 ;
      RECT 49.255000 171.520000 50.185000 171.670000 ;
      RECT 49.255000 171.670000 50.035000 171.820000 ;
      RECT 49.255000 171.820000 49.885000 171.970000 ;
      RECT 49.255000 171.970000 49.735000 172.120000 ;
      RECT 49.255000 172.120000 49.585000 172.270000 ;
      RECT 49.255000 172.270000 49.435000 172.420000 ;
      RECT 49.255000 172.420000 49.285000 172.570000 ;
      RECT 49.255000 172.480000 49.375000 190.420000 ;
      RECT 49.290000   0.000000 49.990000  89.650000 ;
      RECT 49.290000   0.000000 50.090000  90.310000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.310000 55.765000  95.985000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.985000 57.915000  98.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 59.330000  99.550000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.550000 61.200000 101.420000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.310000 101.420000 61.200000 107.795000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.685000 107.795000 61.200000 172.855000 ;
      RECT 59.685000 107.945000 59.835000 108.095000 ;
      RECT 59.685000 108.095000 59.985000 108.245000 ;
      RECT 59.685000 108.245000 60.135000 108.395000 ;
      RECT 59.685000 108.395000 60.285000 108.545000 ;
      RECT 59.685000 108.545000 60.435000 108.695000 ;
      RECT 59.685000 108.695000 60.585000 108.845000 ;
      RECT 59.685000 108.845000 60.735000 108.995000 ;
      RECT 59.685000 108.995000 60.885000 109.145000 ;
      RECT 59.685000 109.145000 61.035000 109.210000 ;
      RECT 59.685000 109.210000 61.100000 172.855000 ;
      RECT 59.685000 172.855000 61.200000 173.620000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.835000 172.855000 61.100000 173.005000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.985000 173.005000 61.100000 173.155000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.135000 173.155000 61.100000 173.305000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.285000 173.305000 61.100000 173.455000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.435000 173.455000 61.100000 173.605000 ;
      RECT 60.450000 173.620000 75.000000 185.195000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 173.605000 61.100000 173.720000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.450000 174.470000 75.000000 174.620000 ;
      RECT 61.450000 174.470000 75.000000 174.620000 ;
      RECT 61.600000 174.620000 75.000000 174.770000 ;
      RECT 61.600000 174.620000 75.000000 174.770000 ;
      RECT 61.750000 174.770000 75.000000 174.920000 ;
      RECT 61.750000 174.770000 75.000000 174.920000 ;
      RECT 61.900000 174.920000 75.000000 175.070000 ;
      RECT 61.900000 174.920000 75.000000 175.070000 ;
      RECT 62.050000 175.070000 75.000000 175.220000 ;
      RECT 62.050000 175.070000 75.000000 175.220000 ;
      RECT 62.200000 175.220000 75.000000 175.370000 ;
      RECT 62.200000 175.220000 75.000000 175.370000 ;
      RECT 62.350000 175.370000 75.000000 175.520000 ;
      RECT 62.350000 175.370000 75.000000 175.520000 ;
      RECT 62.500000 175.520000 75.000000 175.670000 ;
      RECT 62.500000 175.520000 75.000000 175.670000 ;
      RECT 62.650000 175.670000 75.000000 175.820000 ;
      RECT 62.650000 175.670000 75.000000 175.820000 ;
      RECT 62.800000 175.820000 75.000000 175.970000 ;
      RECT 62.800000 175.820000 75.000000 175.970000 ;
      RECT 62.950000 175.970000 75.000000 176.120000 ;
      RECT 62.950000 175.970000 75.000000 176.120000 ;
      RECT 63.100000 176.120000 75.000000 176.270000 ;
      RECT 63.100000 176.120000 75.000000 176.270000 ;
      RECT 63.250000 176.270000 75.000000 176.420000 ;
      RECT 63.250000 176.270000 75.000000 176.420000 ;
      RECT 63.400000 176.420000 75.000000 176.570000 ;
      RECT 63.400000 176.420000 75.000000 176.570000 ;
      RECT 63.550000 176.570000 75.000000 176.720000 ;
      RECT 63.550000 176.570000 75.000000 176.720000 ;
      RECT 63.700000 176.720000 75.000000 176.870000 ;
      RECT 63.700000 176.720000 75.000000 176.870000 ;
      RECT 63.850000 176.870000 75.000000 177.020000 ;
      RECT 63.850000 176.870000 75.000000 177.020000 ;
      RECT 64.000000 177.020000 75.000000 177.170000 ;
      RECT 64.000000 177.020000 75.000000 177.170000 ;
      RECT 64.150000 177.170000 75.000000 177.320000 ;
      RECT 64.150000 177.170000 75.000000 177.320000 ;
      RECT 64.300000 177.320000 75.000000 177.470000 ;
      RECT 64.300000 177.320000 75.000000 177.470000 ;
      RECT 64.450000 177.470000 75.000000 177.620000 ;
      RECT 64.450000 177.470000 75.000000 177.620000 ;
      RECT 64.600000 177.620000 75.000000 177.770000 ;
      RECT 64.600000 177.620000 75.000000 177.770000 ;
      RECT 64.750000 177.770000 75.000000 177.920000 ;
      RECT 64.750000 177.770000 75.000000 177.920000 ;
      RECT 64.900000 177.920000 75.000000 178.070000 ;
      RECT 64.900000 177.920000 75.000000 178.070000 ;
      RECT 65.050000 178.070000 75.000000 178.220000 ;
      RECT 65.050000 178.070000 75.000000 178.220000 ;
      RECT 65.200000 178.220000 75.000000 178.370000 ;
      RECT 65.200000 178.220000 75.000000 178.370000 ;
      RECT 65.350000 178.370000 75.000000 178.520000 ;
      RECT 65.350000 178.370000 75.000000 178.520000 ;
      RECT 65.500000 178.520000 75.000000 178.670000 ;
      RECT 65.500000 178.520000 75.000000 178.670000 ;
      RECT 65.650000 178.670000 75.000000 178.820000 ;
      RECT 65.650000 178.670000 75.000000 178.820000 ;
      RECT 65.800000 178.820000 75.000000 178.970000 ;
      RECT 65.800000 178.820000 75.000000 178.970000 ;
      RECT 65.950000 178.970000 75.000000 179.120000 ;
      RECT 65.950000 178.970000 75.000000 179.120000 ;
      RECT 66.100000 179.120000 75.000000 179.270000 ;
      RECT 66.100000 179.120000 75.000000 179.270000 ;
      RECT 66.250000 179.270000 75.000000 179.420000 ;
      RECT 66.250000 179.270000 75.000000 179.420000 ;
      RECT 66.400000 179.420000 75.000000 179.570000 ;
      RECT 66.400000 179.420000 75.000000 179.570000 ;
      RECT 66.550000 179.570000 75.000000 179.720000 ;
      RECT 66.550000 179.570000 75.000000 179.720000 ;
      RECT 66.700000 179.720000 75.000000 179.870000 ;
      RECT 66.700000 179.720000 75.000000 179.870000 ;
      RECT 66.850000 179.870000 75.000000 180.020000 ;
      RECT 66.850000 179.870000 75.000000 180.020000 ;
      RECT 67.000000 180.020000 75.000000 180.170000 ;
      RECT 67.000000 180.020000 75.000000 180.170000 ;
      RECT 67.150000 180.170000 75.000000 180.320000 ;
      RECT 67.150000 180.170000 75.000000 180.320000 ;
      RECT 67.300000 180.320000 75.000000 180.470000 ;
      RECT 67.300000 180.320000 75.000000 180.470000 ;
      RECT 67.450000 180.470000 75.000000 180.620000 ;
      RECT 67.450000 180.470000 75.000000 180.620000 ;
      RECT 67.600000 180.620000 75.000000 180.770000 ;
      RECT 67.600000 180.620000 75.000000 180.770000 ;
      RECT 67.750000 180.770000 75.000000 180.920000 ;
      RECT 67.750000 180.770000 75.000000 180.920000 ;
      RECT 67.900000 180.920000 75.000000 181.070000 ;
      RECT 67.900000 180.920000 75.000000 181.070000 ;
      RECT 68.050000 181.070000 75.000000 181.220000 ;
      RECT 68.050000 181.070000 75.000000 181.220000 ;
      RECT 68.200000 181.220000 75.000000 181.370000 ;
      RECT 68.200000 181.220000 75.000000 181.370000 ;
      RECT 68.350000 181.370000 75.000000 181.520000 ;
      RECT 68.350000 181.370000 75.000000 181.520000 ;
      RECT 68.500000 181.520000 75.000000 181.670000 ;
      RECT 68.500000 181.520000 75.000000 181.670000 ;
      RECT 68.650000 181.670000 75.000000 181.820000 ;
      RECT 68.650000 181.670000 75.000000 181.820000 ;
      RECT 68.800000 181.820000 75.000000 181.970000 ;
      RECT 68.800000 181.820000 75.000000 181.970000 ;
      RECT 68.950000 181.970000 75.000000 182.120000 ;
      RECT 68.950000 181.970000 75.000000 182.120000 ;
      RECT 69.100000 182.120000 75.000000 182.270000 ;
      RECT 69.100000 182.120000 75.000000 182.270000 ;
      RECT 69.250000 182.270000 75.000000 182.420000 ;
      RECT 69.250000 182.270000 75.000000 182.420000 ;
      RECT 69.400000 182.420000 75.000000 182.570000 ;
      RECT 69.400000 182.420000 75.000000 182.570000 ;
      RECT 69.550000 182.570000 75.000000 182.720000 ;
      RECT 69.550000 182.570000 75.000000 182.720000 ;
      RECT 69.700000 182.720000 75.000000 182.870000 ;
      RECT 69.700000 182.720000 75.000000 182.870000 ;
      RECT 69.850000 182.870000 75.000000 183.020000 ;
      RECT 69.850000 182.870000 75.000000 183.020000 ;
      RECT 70.000000 183.020000 75.000000 183.170000 ;
      RECT 70.000000 183.020000 75.000000 183.170000 ;
      RECT 70.150000 183.170000 75.000000 183.320000 ;
      RECT 70.150000 183.170000 75.000000 183.320000 ;
      RECT 70.300000 183.320000 75.000000 183.470000 ;
      RECT 70.300000 183.320000 75.000000 183.470000 ;
      RECT 70.450000 183.470000 75.000000 183.620000 ;
      RECT 70.450000 183.470000 75.000000 183.620000 ;
      RECT 70.600000 183.620000 75.000000 183.770000 ;
      RECT 70.600000 183.620000 75.000000 183.770000 ;
      RECT 70.750000 183.770000 75.000000 183.920000 ;
      RECT 70.750000 183.770000 75.000000 183.920000 ;
      RECT 70.900000 183.920000 75.000000 184.070000 ;
      RECT 70.900000 183.920000 75.000000 184.070000 ;
      RECT 71.050000 184.070000 75.000000 184.220000 ;
      RECT 71.050000 184.070000 75.000000 184.220000 ;
      RECT 71.200000 184.220000 75.000000 184.370000 ;
      RECT 71.200000 184.220000 75.000000 184.370000 ;
      RECT 71.350000 184.370000 75.000000 184.520000 ;
      RECT 71.350000 184.370000 75.000000 184.520000 ;
      RECT 71.500000 184.520000 75.000000 184.670000 ;
      RECT 71.500000 184.520000 75.000000 184.670000 ;
      RECT 71.650000 184.670000 75.000000 184.820000 ;
      RECT 71.650000 184.670000 75.000000 184.820000 ;
      RECT 71.800000 184.820000 75.000000 184.970000 ;
      RECT 71.800000 184.820000 75.000000 184.970000 ;
      RECT 71.950000 184.970000 75.000000 185.120000 ;
      RECT 71.950000 184.970000 75.000000 185.120000 ;
      RECT 72.025000 185.195000 75.000000 190.440000 ;
      RECT 72.025000 185.345000 72.175000 185.495000 ;
      RECT 72.025000 185.495000 72.325000 185.645000 ;
      RECT 72.025000 185.645000 72.475000 185.795000 ;
      RECT 72.025000 185.795000 72.625000 185.945000 ;
      RECT 72.025000 185.945000 72.775000 186.095000 ;
      RECT 72.025000 186.095000 72.925000 186.245000 ;
      RECT 72.025000 186.245000 73.075000 186.395000 ;
      RECT 72.025000 186.395000 73.225000 186.545000 ;
      RECT 72.025000 186.545000 73.375000 186.695000 ;
      RECT 72.025000 186.695000 73.525000 186.845000 ;
      RECT 72.025000 186.845000 73.675000 186.995000 ;
      RECT 72.025000 186.995000 73.825000 187.145000 ;
      RECT 72.025000 187.145000 73.975000 187.295000 ;
      RECT 72.025000 187.295000 74.125000 187.445000 ;
      RECT 72.025000 187.445000 74.275000 187.595000 ;
      RECT 72.025000 187.595000 74.425000 187.745000 ;
      RECT 72.025000 187.745000 74.575000 187.895000 ;
      RECT 72.025000 187.895000 74.725000 188.045000 ;
      RECT 72.025000 188.045000 74.875000 188.170000 ;
      RECT 72.025000 188.170000 75.000000 190.440000 ;
      RECT 72.100000 185.120000 75.000000 185.270000 ;
      RECT 72.100000 185.120000 75.000000 185.270000 ;
      RECT 72.250000 185.270000 75.000000 185.420000 ;
      RECT 72.250000 185.270000 75.000000 185.420000 ;
      RECT 72.400000 185.420000 75.000000 185.570000 ;
      RECT 72.400000 185.420000 75.000000 185.570000 ;
      RECT 72.550000 185.570000 75.000000 185.720000 ;
      RECT 72.550000 185.570000 75.000000 185.720000 ;
      RECT 72.700000 185.720000 75.000000 185.870000 ;
      RECT 72.700000 185.720000 75.000000 185.870000 ;
      RECT 72.850000 185.870000 75.000000 186.020000 ;
      RECT 72.850000 185.870000 75.000000 186.020000 ;
      RECT 73.000000 186.020000 75.000000 186.170000 ;
      RECT 73.000000 186.020000 75.000000 186.170000 ;
      RECT 73.150000 186.170000 75.000000 186.320000 ;
      RECT 73.150000 186.170000 75.000000 186.320000 ;
      RECT 73.300000 186.320000 75.000000 186.470000 ;
      RECT 73.300000 186.320000 75.000000 186.470000 ;
      RECT 73.450000 186.470000 75.000000 186.620000 ;
      RECT 73.450000 186.470000 75.000000 186.620000 ;
      RECT 73.600000 186.620000 75.000000 186.770000 ;
      RECT 73.600000 186.620000 75.000000 186.770000 ;
      RECT 73.750000 186.770000 75.000000 186.920000 ;
      RECT 73.750000 186.770000 75.000000 186.920000 ;
      RECT 73.900000 186.920000 75.000000 187.070000 ;
      RECT 73.900000 186.920000 75.000000 187.070000 ;
      RECT 74.050000 187.070000 75.000000 187.220000 ;
      RECT 74.050000 187.070000 75.000000 187.220000 ;
      RECT 74.200000 187.220000 75.000000 187.370000 ;
      RECT 74.200000 187.220000 75.000000 187.370000 ;
      RECT 74.350000 187.370000 75.000000 187.520000 ;
      RECT 74.350000 187.370000 75.000000 187.520000 ;
      RECT 74.500000 187.520000 75.000000 187.670000 ;
      RECT 74.500000 187.520000 75.000000 187.670000 ;
      RECT 74.590000   0.000000 75.000000 173.620000 ;
      RECT 74.650000 187.670000 75.000000 187.820000 ;
      RECT 74.650000 187.670000 75.000000 187.820000 ;
      RECT 74.690000   0.000000 75.000000 173.720000 ;
      RECT 74.800000 187.820000 75.000000 187.970000 ;
      RECT 74.800000 187.820000 75.000000 187.970000 ;
      RECT 74.950000 187.970000 75.000000 188.120000 ;
      RECT 74.950000 187.970000 75.000000 188.120000 ;
    LAYER met4 ;
      RECT  4.800000 104.380000  5.160000 104.530000 ;
      RECT  4.800000 104.530000  5.525000 104.680000 ;
      RECT  4.800000 104.680000  5.885000 104.830000 ;
      RECT  4.800000 104.830000  6.245000 104.980000 ;
      RECT  4.800000 104.980000  6.610000 105.130000 ;
      RECT  4.800000 105.130000  6.970000 105.280000 ;
      RECT  4.800000 105.280000  7.330000 105.350000 ;
      RECT  4.800000 105.350000  7.500000 165.450000 ;
      RECT  4.800000 165.450000  7.500000 165.600000 ;
      RECT  4.800000 165.600000  7.650000 165.750000 ;
      RECT  4.800000 165.750000  7.800000 165.900000 ;
      RECT  4.800000 165.900000  7.950000 166.050000 ;
      RECT  4.800000 166.050000  8.100000 166.200000 ;
      RECT  4.800000 166.200000  8.250000 166.350000 ;
      RECT  4.800000 166.350000  8.400000 166.500000 ;
      RECT  4.800000 166.500000  8.550000 166.570000 ;
      RECT  4.840000 104.265000  7.460000 165.545000 ;
      RECT  4.880000 104.150000  8.620000 104.230000 ;
      RECT  4.950000 166.570000  8.620000 166.720000 ;
      RECT  5.030000 104.000000  8.700000 104.150000 ;
      RECT  5.100000 166.720000  8.770000 166.870000 ;
      RECT  5.160000 104.230000  8.470000 104.380000 ;
      RECT  5.180000 103.850000  8.850000 104.000000 ;
      RECT  5.250000 166.870000  8.920000 167.020000 ;
      RECT  5.330000 103.700000  9.000000 103.850000 ;
      RECT  5.400000 167.020000  9.070000 167.170000 ;
      RECT  5.470000 165.675000  7.595000 167.175000 ;
      RECT  5.480000 103.550000  9.150000 103.700000 ;
      RECT  5.525000 104.380000  8.320000 104.530000 ;
      RECT  5.550000 167.170000  9.220000 167.320000 ;
      RECT  5.630000 103.400000  9.300000 103.550000 ;
      RECT  5.655000 103.425000  6.280000 104.075000 ;
      RECT  5.700000 167.320000  9.370000 167.470000 ;
      RECT  5.780000 103.250000  9.450000 103.400000 ;
      RECT  5.850000 167.470000  9.520000 167.620000 ;
      RECT  5.885000 104.530000  8.170000 104.680000 ;
      RECT  5.930000 103.100000  9.600000 103.250000 ;
      RECT  6.000000 167.620000  9.670000 167.770000 ;
      RECT  6.080000 102.950000  9.750000 103.100000 ;
      RECT  6.150000 167.770000  9.820000 167.920000 ;
      RECT  6.230000 102.800000  9.900000 102.950000 ;
      RECT  6.235000 167.300000  6.860000 167.950000 ;
      RECT  6.245000 104.680000  8.020000 104.830000 ;
      RECT  6.300000 167.920000  9.970000 168.070000 ;
      RECT  6.380000 102.650000 10.050000 102.800000 ;
      RECT  6.450000 168.070000 10.120000 168.220000 ;
      RECT  6.510000 102.630000  8.635000 104.130000 ;
      RECT  6.530000 102.500000 10.200000 102.650000 ;
      RECT  6.600000 168.220000 10.270000 168.370000 ;
      RECT  6.610000 104.830000  7.870000 104.980000 ;
      RECT  6.680000 102.350000 10.350000 102.500000 ;
      RECT  6.750000 168.370000 10.420000 168.520000 ;
      RECT  6.830000 102.200000 10.500000 102.350000 ;
      RECT  6.900000 168.520000 10.570000 168.670000 ;
      RECT  6.970000 104.980000  7.720000 105.130000 ;
      RECT  6.980000 102.050000 10.650000 102.200000 ;
      RECT  7.050000 168.670000 10.720000 168.820000 ;
      RECT  7.070000 167.275000  9.195000 168.775000 ;
      RECT  7.130000 101.900000 10.800000 102.050000 ;
      RECT  7.200000 168.820000 10.870000 168.970000 ;
      RECT  7.275000 101.855000  7.900000 102.505000 ;
      RECT  7.280000 101.750000 10.950000 101.900000 ;
      RECT  7.310000 104.205000  7.935000 104.855000 ;
      RECT  7.330000 105.130000  7.570000 105.280000 ;
      RECT  7.350000 168.970000 11.020000 169.120000 ;
      RECT  7.430000 101.600000 11.100000 101.750000 ;
      RECT  7.500000 169.120000 11.170000 169.270000 ;
      RECT  7.580000 101.450000 11.250000 101.600000 ;
      RECT  7.650000 169.270000 11.320000 169.420000 ;
      RECT  7.675000 166.490000  8.300000 167.140000 ;
      RECT  7.730000 101.300000 11.400000 101.450000 ;
      RECT  7.800000 169.420000 11.470000 169.570000 ;
      RECT  7.875000 168.940000  8.500000 169.590000 ;
      RECT  7.880000 101.150000 11.550000 101.300000 ;
      RECT  7.950000 169.570000 11.620000 169.720000 ;
      RECT  8.030000 101.000000 11.700000 101.150000 ;
      RECT  8.100000 169.720000 11.770000 169.870000 ;
      RECT  8.110000 101.030000 10.235000 102.530000 ;
      RECT  8.180000 100.850000 11.850000 101.000000 ;
      RECT  8.250000 169.870000 11.920000 170.020000 ;
      RECT  8.330000 100.700000 12.000000 100.850000 ;
      RECT  8.400000 170.020000 12.070000 170.170000 ;
      RECT  8.480000 100.550000 12.150000 100.700000 ;
      RECT  8.550000 170.170000 12.220000 170.320000 ;
      RECT  8.630000 100.400000 12.300000 100.550000 ;
      RECT  8.630000 170.320000 12.370000 170.400000 ;
      RECT  8.690000 168.895000 10.815000 170.395000 ;
      RECT  8.715000 102.665000  9.340000 103.315000 ;
      RECT  8.780000 100.250000 62.550000 100.400000 ;
      RECT  8.780000 170.400000 12.390000 170.550000 ;
      RECT  8.915000 100.215000  9.540000 100.865000 ;
      RECT  8.930000 100.100000 62.610000 100.250000 ;
      RECT  8.930000 170.550000 12.325000 170.700000 ;
      RECT  9.080000  99.950000 62.675000 100.100000 ;
      RECT  9.080000 170.700000 12.265000 170.850000 ;
      RECT  9.230000  99.800000 62.735000  99.950000 ;
      RECT  9.230000 170.850000 12.200000 171.000000 ;
      RECT  9.300000 168.115000  9.925000 168.765000 ;
      RECT  9.320000 170.425000  9.730000 171.075000 ;
      RECT  9.380000  99.650000 62.800000  99.800000 ;
      RECT  9.380000 171.000000 12.140000 171.150000 ;
      RECT  9.530000  99.500000 62.860000  99.650000 ;
      RECT  9.530000 171.150000 12.075000 171.300000 ;
      RECT  9.680000  99.350000 62.925000  99.500000 ;
      RECT  9.680000 171.300000 12.015000 171.450000 ;
      RECT  9.730000  99.410000 11.855000 100.910000 ;
      RECT  9.830000  99.200000 62.985000  99.350000 ;
      RECT  9.830000 171.450000 11.950000 171.600000 ;
      RECT  9.965000 170.770000 11.105000 171.580000 ;
      RECT  9.980000  99.050000 63.050000  99.200000 ;
      RECT  9.980000 171.600000 11.890000 171.750000 ;
      RECT 10.130000  98.900000 63.110000  99.050000 ;
      RECT 10.130000 171.750000 11.830000 171.900000 ;
      RECT 10.280000  98.750000 63.170000  98.900000 ;
      RECT 10.280000 171.900000 11.765000 172.050000 ;
      RECT 10.340000 101.040000 10.965000 101.690000 ;
      RECT 10.430000  98.600000 63.235000  98.750000 ;
      RECT 10.430000 172.050000 11.705000 172.200000 ;
      RECT 10.580000  98.450000 63.295000  98.600000 ;
      RECT 10.580000 172.200000 11.640000 172.350000 ;
      RECT 10.610000 171.715000 11.020000 172.365000 ;
      RECT 10.620000  98.510000 11.245000  99.160000 ;
      RECT 10.730000  98.300000 63.360000  98.450000 ;
      RECT 10.730000 172.350000 11.580000 172.500000 ;
      RECT 10.880000  98.150000 63.420000  98.300000 ;
      RECT 10.880000 172.500000 11.515000 172.650000 ;
      RECT 10.890000 169.555000 11.515000 170.205000 ;
      RECT 11.030000  98.000000 63.485000  98.150000 ;
      RECT 11.030000 172.650000 11.455000 172.800000 ;
      RECT 11.180000  97.850000 63.545000  98.000000 ;
      RECT 11.180000 172.800000 11.390000 172.950000 ;
      RECT 11.330000  97.700000 63.610000  97.850000 ;
      RECT 11.330000 170.400000 13.335000 173.100000 ;
      RECT 11.390000 172.950000 63.670000 173.100000 ;
      RECT 11.455000 172.800000 63.820000 172.950000 ;
      RECT 11.515000 172.650000 63.970000 172.800000 ;
      RECT 11.580000 172.500000 64.120000 172.650000 ;
      RECT 11.640000 172.350000 64.270000 172.500000 ;
      RECT 11.705000 172.200000 64.420000 172.350000 ;
      RECT 11.765000 172.050000 64.570000 172.200000 ;
      RECT 11.830000 171.900000 64.720000 172.050000 ;
      RECT 11.890000 171.750000 64.870000 171.900000 ;
      RECT 11.950000 171.600000 65.020000 171.750000 ;
      RECT 12.015000 171.450000 65.170000 171.600000 ;
      RECT 12.075000 171.300000 65.320000 171.450000 ;
      RECT 12.140000 171.150000 65.470000 171.300000 ;
      RECT 12.200000 171.000000 65.620000 171.150000 ;
      RECT 12.265000 170.850000 65.770000 171.000000 ;
      RECT 12.325000 170.700000 65.920000 170.850000 ;
      RECT 12.390000 170.550000 66.070000 170.700000 ;
      RECT 12.450000 170.400000 66.220000 170.550000 ;
      RECT 58.800000  97.740000 59.420000  98.535000 ;
      RECT 59.465000  97.725000 63.575000  99.225000 ;
      RECT 60.180000  99.285000 60.630000  99.935000 ;
      RECT 60.700000  99.420000 62.760000 100.350000 ;
      RECT 61.655000 170.400000 63.665000 173.100000 ;
      RECT 62.610000 100.250000 66.220000 100.400000 ;
      RECT 62.630000 170.320000 66.370000 170.400000 ;
      RECT 62.675000 100.100000 66.070000 100.250000 ;
      RECT 62.700000 100.400000 66.370000 100.550000 ;
      RECT 62.735000  99.950000 65.920000 100.100000 ;
      RECT 62.780000 170.170000 66.450000 170.320000 ;
      RECT 62.800000  99.800000 65.770000  99.950000 ;
      RECT 62.850000 100.550000 66.520000 100.700000 ;
      RECT 62.860000  99.650000 65.620000  99.800000 ;
      RECT 62.925000  99.500000 65.470000  99.650000 ;
      RECT 62.930000 170.020000 66.600000 170.170000 ;
      RECT 62.985000  99.350000 65.320000  99.500000 ;
      RECT 63.000000 100.700000 66.670000 100.850000 ;
      RECT 63.050000  99.200000 65.170000  99.350000 ;
      RECT 63.080000 169.870000 66.750000 170.020000 ;
      RECT 63.110000  99.050000 65.020000  99.200000 ;
      RECT 63.135000  99.410000 65.260000 100.910000 ;
      RECT 63.150000 100.850000 66.820000 101.000000 ;
      RECT 63.170000  98.900000 64.870000  99.050000 ;
      RECT 63.230000 169.720000 66.900000 169.870000 ;
      RECT 63.235000  98.750000 64.720000  98.900000 ;
      RECT 63.295000  98.600000 64.570000  98.750000 ;
      RECT 63.300000 101.000000 66.970000 101.150000 ;
      RECT 63.360000  98.450000 64.420000  98.600000 ;
      RECT 63.380000 169.570000 67.050000 169.720000 ;
      RECT 63.420000  98.300000 64.270000  98.450000 ;
      RECT 63.450000 101.150000 67.120000 101.300000 ;
      RECT 63.475000 169.555000 64.100000 170.205000 ;
      RECT 63.485000  98.150000 64.120000  98.300000 ;
      RECT 63.530000 169.420000 67.200000 169.570000 ;
      RECT 63.545000  98.000000 63.970000  98.150000 ;
      RECT 63.600000 101.300000 67.270000 101.450000 ;
      RECT 63.610000  97.850000 63.820000  98.000000 ;
      RECT 63.680000 169.270000 67.350000 169.420000 ;
      RECT 63.745000  98.510000 64.370000  99.160000 ;
      RECT 63.750000 101.450000 67.420000 101.600000 ;
      RECT 63.830000 169.120000 67.500000 169.270000 ;
      RECT 63.885000 170.770000 65.025000 171.580000 ;
      RECT 63.900000 101.600000 67.570000 101.750000 ;
      RECT 63.970000 171.715000 64.380000 172.365000 ;
      RECT 63.980000 168.970000 67.650000 169.120000 ;
      RECT 64.025000 101.040000 64.650000 101.690000 ;
      RECT 64.050000 101.750000 67.720000 101.900000 ;
      RECT 64.130000 168.820000 67.800000 168.970000 ;
      RECT 64.175000 168.895000 66.300000 170.395000 ;
      RECT 64.200000 101.900000 67.870000 102.050000 ;
      RECT 64.280000 168.670000 67.950000 168.820000 ;
      RECT 64.350000 102.050000 68.020000 102.200000 ;
      RECT 64.430000 168.520000 68.100000 168.670000 ;
      RECT 64.500000 102.200000 68.170000 102.350000 ;
      RECT 64.580000 168.370000 68.250000 168.520000 ;
      RECT 64.650000 102.350000 68.320000 102.500000 ;
      RECT 64.730000 168.220000 68.400000 168.370000 ;
      RECT 64.755000 101.030000 66.880000 102.530000 ;
      RECT 64.800000 102.500000 68.470000 102.650000 ;
      RECT 64.880000 168.070000 68.550000 168.220000 ;
      RECT 64.950000 102.650000 68.620000 102.800000 ;
      RECT 65.030000 167.920000 68.700000 168.070000 ;
      RECT 65.065000 168.115000 65.690000 168.765000 ;
      RECT 65.100000 102.800000 68.770000 102.950000 ;
      RECT 65.180000 167.770000 68.850000 167.920000 ;
      RECT 65.250000 102.950000 68.920000 103.100000 ;
      RECT 65.260000 170.425000 65.670000 171.075000 ;
      RECT 65.330000 167.620000 69.000000 167.770000 ;
      RECT 65.400000 103.100000 69.070000 103.250000 ;
      RECT 65.450000 100.215000 66.075000 100.865000 ;
      RECT 65.480000 167.470000 69.150000 167.620000 ;
      RECT 65.550000 103.250000 69.220000 103.400000 ;
      RECT 65.630000 167.320000 69.300000 167.470000 ;
      RECT 65.650000 102.665000 66.275000 103.315000 ;
      RECT 65.700000 103.400000 69.370000 103.550000 ;
      RECT 65.780000 167.170000 69.450000 167.320000 ;
      RECT 65.795000 167.275000 67.920000 168.775000 ;
      RECT 65.850000 103.550000 69.520000 103.700000 ;
      RECT 65.930000 167.020000 69.600000 167.170000 ;
      RECT 66.000000 103.700000 69.670000 103.850000 ;
      RECT 66.080000 166.870000 69.750000 167.020000 ;
      RECT 66.150000 103.850000 69.820000 104.000000 ;
      RECT 66.230000 166.720000 69.900000 166.870000 ;
      RECT 66.300000 104.000000 69.970000 104.150000 ;
      RECT 66.355000 102.630000 68.480000 104.130000 ;
      RECT 66.380000 104.150000 70.120000 104.230000 ;
      RECT 66.380000 166.570000 70.050000 166.720000 ;
      RECT 66.450000 166.500000 70.030000 166.570000 ;
      RECT 66.490000 168.940000 67.115000 169.590000 ;
      RECT 66.530000 104.230000 70.200000 104.380000 ;
      RECT 66.600000 166.350000 69.670000 166.500000 ;
      RECT 66.680000 104.380000 70.200000 104.530000 ;
      RECT 66.690000 166.490000 67.315000 167.140000 ;
      RECT 66.750000 166.200000 69.310000 166.350000 ;
      RECT 66.830000 104.530000 70.200000 104.680000 ;
      RECT 66.900000 166.050000 68.945000 166.200000 ;
      RECT 66.980000 104.680000 70.200000 104.830000 ;
      RECT 67.050000 165.900000 68.585000 166.050000 ;
      RECT 67.055000 104.205000 67.680000 104.855000 ;
      RECT 67.090000 101.855000 67.715000 102.505000 ;
      RECT 67.130000 104.830000 70.200000 104.980000 ;
      RECT 67.200000 165.750000 68.225000 165.900000 ;
      RECT 67.280000 104.980000 70.200000 105.130000 ;
      RECT 67.350000 165.600000 67.860000 165.750000 ;
      RECT 67.395000 165.675000 69.520000 167.175000 ;
      RECT 67.430000 105.130000 70.200000 105.280000 ;
      RECT 67.500000 105.280000 70.200000 105.350000 ;
      RECT 67.500000 105.350000 70.200000 165.450000 ;
      RECT 67.530000 104.265000 70.150000 165.545000 ;
      RECT 67.860000 165.450000 70.200000 165.600000 ;
      RECT 68.130000 167.300000 68.755000 167.950000 ;
      RECT 68.225000 165.600000 70.200000 165.750000 ;
      RECT 68.550000 103.230000 69.170000 104.115000 ;
      RECT 68.585000 165.750000 70.200000 165.900000 ;
      RECT 68.945000 165.900000 70.200000 166.050000 ;
      RECT 69.200000 103.590000 69.535000 104.240000 ;
      RECT 69.310000 166.050000 70.200000 166.200000 ;
      RECT 69.670000 166.200000 70.200000 166.350000 ;
      RECT 70.030000 166.350000 70.200000 166.500000 ;
  END
END sky130_fd_io__top_power_hvc_wpad
MACRO sky130_fd_io__top_gpiov2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430000 0.000000 62.690000 1.915000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865000  0.000000 46.195000 36.665000 ;
        RECT 45.865000 36.665000 46.195000 36.735000 ;
        RECT 45.865000 36.735000 46.265000 36.805000 ;
        RECT 45.965000 36.805000 46.335000 36.905000 ;
        RECT 46.065000 36.905000 46.435000 37.005000 ;
        RECT 46.070000 37.005000 46.535000 37.010000 ;
        RECT 46.220000 37.010000 48.225000 37.160000 ;
        RECT 46.370000 37.160000 48.075000 37.310000 ;
        RECT 46.400000 37.310000 48.045000 37.340000 ;
        RECT 47.910000 37.005000 48.375000 37.010000 ;
        RECT 47.960000 35.870000 48.740000 36.190000 ;
        RECT 47.975000 36.940000 48.380000 37.005000 ;
        RECT 48.040000 36.875000 48.445000 36.940000 ;
        RECT 48.070000 36.190000 48.630000 36.300000 ;
        RECT 48.110000 36.805000 48.510000 36.875000 ;
        RECT 48.180000 36.300000 48.520000 36.410000 ;
        RECT 48.180000 36.410000 48.515000 36.415000 ;
        RECT 48.180000 36.415000 48.510000 36.420000 ;
        RECT 48.180000 36.420000 48.510000 36.735000 ;
        RECT 48.180000 36.735000 48.510000 36.805000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.080000 57.360000 24.590000 57.430000 ;
        RECT 23.080000 57.430000 24.520000 57.500000 ;
        RECT 23.080000 57.500000 24.450000 57.570000 ;
        RECT 23.080000 57.570000 24.380000 57.640000 ;
        RECT 24.285000 57.345000 24.660000 57.360000 ;
        RECT 24.355000 57.275000 24.675000 57.345000 ;
        RECT 24.425000 57.205000 24.745000 57.275000 ;
        RECT 24.495000 57.135000 24.815000 57.205000 ;
        RECT 24.565000 57.065000 24.885000 57.135000 ;
        RECT 24.620000 57.010000 24.955000 57.065000 ;
        RECT 24.675000 53.255000 25.010000 53.310000 ;
        RECT 24.675000 53.310000 24.955000 53.365000 ;
        RECT 24.675000 53.365000 24.955000 56.955000 ;
        RECT 24.675000 56.955000 24.955000 57.010000 ;
        RECT 24.740000 53.190000 25.065000 53.255000 ;
        RECT 24.810000 53.120000 25.130000 53.190000 ;
        RECT 24.880000 53.050000 25.200000 53.120000 ;
        RECT 24.950000 52.980000 25.270000 53.050000 ;
        RECT 25.020000 52.910000 25.340000 52.980000 ;
        RECT 25.090000 52.840000 25.410000 52.910000 ;
        RECT 25.160000 52.770000 25.480000 52.840000 ;
        RECT 25.230000 52.700000 25.550000 52.770000 ;
        RECT 25.300000 52.630000 25.620000 52.700000 ;
        RECT 25.370000 52.560000 25.690000 52.630000 ;
        RECT 25.440000 52.490000 25.760000 52.560000 ;
        RECT 25.510000 52.420000 25.830000 52.490000 ;
        RECT 25.580000 52.350000 25.900000 52.420000 ;
        RECT 25.650000 52.280000 25.970000 52.350000 ;
        RECT 25.720000 52.210000 26.040000 52.280000 ;
        RECT 25.790000 52.140000 29.735000 52.210000 ;
        RECT 25.860000 52.070000 29.805000 52.140000 ;
        RECT 25.930000 52.000000 29.875000 52.070000 ;
        RECT 26.000000 51.930000 29.945000 52.000000 ;
        RECT 29.645000 51.910000 30.015000 51.930000 ;
        RECT 29.715000 51.840000 30.035000 51.910000 ;
        RECT 29.785000 51.770000 30.105000 51.840000 ;
        RECT 29.855000 51.700000 30.175000 51.770000 ;
        RECT 29.925000 51.630000 30.245000 51.700000 ;
        RECT 29.995000 51.560000 30.315000 51.630000 ;
        RECT 30.060000 51.495000 30.385000 51.560000 ;
        RECT 30.125000 17.630000 30.440000 17.685000 ;
        RECT 30.125000 17.685000 30.385000 17.740000 ;
        RECT 30.125000 17.740000 30.385000 36.345000 ;
        RECT 30.125000 36.345000 30.385000 36.400000 ;
        RECT 30.125000 36.400000 30.440000 36.455000 ;
        RECT 30.125000 38.010000 30.440000 38.065000 ;
        RECT 30.125000 38.065000 30.385000 38.120000 ;
        RECT 30.125000 38.120000 30.385000 51.430000 ;
        RECT 30.125000 51.430000 30.385000 51.495000 ;
        RECT 30.140000 37.995000 30.495000 38.010000 ;
        RECT 30.180000 17.575000 30.495000 17.630000 ;
        RECT 30.195000 36.455000 30.495000 36.525000 ;
        RECT 30.210000 37.925000 30.510000 37.995000 ;
        RECT 30.250000 17.505000 30.550000 17.575000 ;
        RECT 30.265000 36.525000 30.565000 36.595000 ;
        RECT 30.280000 36.595000 30.635000 36.610000 ;
        RECT 30.280000 37.855000 30.580000 37.925000 ;
        RECT 30.320000 17.435000 30.620000 17.505000 ;
        RECT 30.335000 36.610000 30.650000 36.665000 ;
        RECT 30.335000 37.800000 30.650000 37.855000 ;
        RECT 30.390000 17.365000 30.690000 17.435000 ;
        RECT 30.390000 36.665000 30.650000 36.720000 ;
        RECT 30.390000 36.720000 30.650000 37.745000 ;
        RECT 30.390000 37.745000 30.650000 37.800000 ;
        RECT 30.460000 17.295000 30.760000 17.365000 ;
        RECT 30.530000 17.225000 30.830000 17.295000 ;
        RECT 30.600000 17.155000 30.900000 17.225000 ;
        RECT 30.670000 17.085000 30.970000 17.155000 ;
        RECT 30.740000 17.015000 31.040000 17.085000 ;
        RECT 30.750000  0.000000 31.010000  2.155000 ;
        RECT 30.750000  2.155000 31.010000  2.210000 ;
        RECT 30.750000  2.210000 31.065000  2.265000 ;
        RECT 30.810000 16.945000 31.110000 17.015000 ;
        RECT 30.820000  2.265000 31.120000  2.335000 ;
        RECT 30.880000 16.875000 31.180000 16.945000 ;
        RECT 30.890000  2.335000 31.190000  2.405000 ;
        RECT 30.950000 16.805000 31.250000 16.875000 ;
        RECT 30.960000  2.405000 31.260000  2.475000 ;
        RECT 31.020000 16.735000 31.320000 16.805000 ;
        RECT 31.030000  2.475000 31.330000  2.545000 ;
        RECT 31.090000 16.665000 31.390000 16.735000 ;
        RECT 31.100000  2.545000 31.400000  2.615000 ;
        RECT 31.160000 16.595000 31.460000 16.665000 ;
        RECT 31.170000  2.615000 31.470000  2.685000 ;
        RECT 31.195000  2.685000 31.540000  2.710000 ;
        RECT 31.230000 16.525000 31.530000 16.595000 ;
        RECT 31.250000  2.710000 31.565000  2.765000 ;
        RECT 31.300000 16.455000 31.600000 16.525000 ;
        RECT 31.305000  2.765000 31.565000  2.820000 ;
        RECT 31.305000  2.820000 31.565000  4.335000 ;
        RECT 31.305000  4.335000 31.565000  4.390000 ;
        RECT 31.305000  4.390000 31.620000  4.445000 ;
        RECT 31.370000 16.385000 31.670000 16.455000 ;
        RECT 31.375000  4.445000 31.675000  4.515000 ;
        RECT 31.440000 16.315000 31.740000 16.385000 ;
        RECT 31.445000  4.515000 31.745000  4.585000 ;
        RECT 31.510000 16.245000 31.810000 16.315000 ;
        RECT 31.515000  4.585000 31.815000  4.655000 ;
        RECT 31.580000  4.655000 31.885000  4.720000 ;
        RECT 31.580000 16.175000 31.880000 16.245000 ;
        RECT 31.635000  4.720000 31.950000  4.775000 ;
        RECT 31.635000 16.120000 31.950000 16.175000 ;
        RECT 31.690000  4.775000 31.950000  4.830000 ;
        RECT 31.690000  4.830000 31.950000 16.065000 ;
        RECT 31.690000 16.065000 31.950000 16.120000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.590000 0.545000 50.360000 0.825000 ;
        RECT 49.625000 0.510000 50.325000 0.545000 ;
        RECT 49.695000 0.440000 50.255000 0.510000 ;
        RECT 49.765000 0.370000 50.185000 0.440000 ;
        RECT 49.835000 0.300000 50.115000 0.370000 ;
        RECT 49.845000 0.290000 50.115000 0.300000 ;
        RECT 49.855000 0.000000 50.115000 0.280000 ;
        RECT 49.855000 0.280000 50.115000 0.290000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.540000 1.195000 67.360000 1.475000 ;
        RECT 66.595000 1.140000 67.305000 1.195000 ;
        RECT 66.665000 1.070000 67.235000 1.140000 ;
        RECT 66.735000 1.000000 67.165000 1.070000 ;
        RECT 66.805000 0.930000 67.095000 1.000000 ;
        RECT 66.820000 0.915000 67.095000 0.930000 ;
        RECT 66.835000 0.000000 67.095000 0.900000 ;
        RECT 66.835000 0.900000 67.095000 0.915000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490000 0.000000 28.750000 3.960000 ;
        RECT 28.490000 3.960000 28.750000 4.015000 ;
        RECT 28.490000 4.015000 28.805000 4.070000 ;
        RECT 28.560000 4.070000 28.860000 4.140000 ;
        RECT 28.630000 4.140000 28.930000 4.210000 ;
        RECT 28.700000 4.210000 29.000000 4.280000 ;
        RECT 28.770000 4.280000 29.070000 4.350000 ;
        RECT 28.840000 4.350000 29.140000 4.420000 ;
        RECT 28.910000 4.420000 29.210000 4.490000 ;
        RECT 28.980000 4.490000 29.280000 4.560000 ;
        RECT 29.050000 4.560000 29.350000 4.630000 ;
        RECT 29.100000 4.630000 29.420000 4.680000 ;
        RECT 29.155000 4.680000 29.470000 4.735000 ;
        RECT 29.210000 4.735000 29.470000 4.790000 ;
        RECT 29.210000 4.790000 29.470000 6.780000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  4.860000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.135000 2.225000 35.450000 2.280000 ;
        RECT 35.135000 2.280000 35.395000 2.335000 ;
        RECT 35.135000 2.335000 35.395000 3.885000 ;
        RECT 35.140000 2.220000 35.505000 2.225000 ;
        RECT 35.210000 2.150000 35.510000 2.220000 ;
        RECT 35.280000 2.080000 35.580000 2.150000 ;
        RECT 35.350000 2.010000 35.650000 2.080000 ;
        RECT 35.405000 1.955000 35.720000 2.010000 ;
        RECT 35.460000 0.000000 35.720000 1.900000 ;
        RECT 35.460000 1.900000 35.720000 1.955000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390000 0.000000 38.650000 3.715000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.315000 56.460000  7.630000 56.515000 ;
        RECT  7.315000 56.515000  7.575000 56.570000 ;
        RECT  7.315000 56.570000  7.575000 73.615000 ;
        RECT  7.315000 73.615000  7.575000 73.670000 ;
        RECT  7.315000 73.670000  7.630000 73.725000 ;
        RECT  7.375000 56.400000  7.685000 56.460000 ;
        RECT  7.385000 73.725000  7.685000 73.795000 ;
        RECT  7.445000 56.330000  7.745000 56.400000 ;
        RECT  7.455000 73.795000  7.755000 73.865000 ;
        RECT  7.515000 56.260000  7.815000 56.330000 ;
        RECT  7.525000 73.865000  7.825000 73.935000 ;
        RECT  7.585000 56.190000  7.885000 56.260000 ;
        RECT  7.595000 73.935000  7.895000 74.005000 ;
        RECT  7.655000 56.120000  7.955000 56.190000 ;
        RECT  7.665000 74.005000  7.965000 74.075000 ;
        RECT  7.695000 74.075000  8.035000 74.105000 ;
        RECT  7.725000 56.050000  8.025000 56.120000 ;
        RECT  7.750000 74.105000  8.065000 74.160000 ;
        RECT  7.795000 55.980000  8.095000 56.050000 ;
        RECT  7.805000 74.160000  8.065000 74.215000 ;
        RECT  7.805000 74.215000  8.065000 74.680000 ;
        RECT  7.805000 74.680000  8.065000 74.735000 ;
        RECT  7.805000 74.735000  8.120000 74.790000 ;
        RECT  7.865000 55.910000  8.165000 55.980000 ;
        RECT  7.875000 74.790000  8.175000 74.860000 ;
        RECT  7.920000 55.855000  8.235000 55.910000 ;
        RECT  7.920000 77.285000  8.560000 77.545000 ;
        RECT  7.945000 74.860000  8.245000 74.930000 ;
        RECT  7.975000 53.960000  8.290000 54.015000 ;
        RECT  7.975000 54.015000  8.235000 54.070000 ;
        RECT  7.975000 54.070000  8.235000 55.800000 ;
        RECT  7.975000 55.800000  8.235000 55.855000 ;
        RECT  8.015000 74.930000  8.315000 75.000000 ;
        RECT  8.030000 53.905000  8.345000 53.960000 ;
        RECT  8.085000 53.850000  8.400000 53.905000 ;
        RECT  8.085000 75.000000  8.385000 75.070000 ;
        RECT  8.085000 77.240000  8.515000 77.285000 ;
        RECT  8.100000 75.070000  8.455000 75.085000 ;
        RECT  8.130000 77.195000  8.470000 77.240000 ;
        RECT  8.140000 53.795000  8.455000 53.850000 ;
        RECT  8.155000 75.085000  8.470000 75.140000 ;
        RECT  8.170000 77.155000  8.470000 77.195000 ;
        RECT  8.195000 44.075000  8.510000 44.130000 ;
        RECT  8.195000 44.130000  8.455000 44.185000 ;
        RECT  8.195000 44.185000  8.455000 53.740000 ;
        RECT  8.195000 53.740000  8.455000 53.795000 ;
        RECT  8.210000 44.060000  8.565000 44.075000 ;
        RECT  8.210000 75.140000  8.470000 75.195000 ;
        RECT  8.210000 75.195000  8.470000 77.115000 ;
        RECT  8.210000 77.115000  8.470000 77.155000 ;
        RECT  8.280000 43.990000  8.580000 44.060000 ;
        RECT  8.350000 43.920000  8.650000 43.990000 ;
        RECT  8.420000 43.850000  8.720000 43.920000 ;
        RECT  8.490000 43.780000  8.790000 43.850000 ;
        RECT  8.560000 43.710000  8.860000 43.780000 ;
        RECT  8.630000 43.640000  8.930000 43.710000 ;
        RECT  8.700000 43.570000  9.000000 43.640000 ;
        RECT  8.770000 43.500000  9.070000 43.570000 ;
        RECT  8.840000 43.430000  9.140000 43.500000 ;
        RECT  8.910000 43.360000  9.210000 43.430000 ;
        RECT  8.980000 43.290000  9.280000 43.360000 ;
        RECT  9.050000 43.220000  9.350000 43.290000 ;
        RECT  9.120000 43.150000  9.420000 43.220000 ;
        RECT  9.190000 43.080000  9.490000 43.150000 ;
        RECT  9.260000 43.010000  9.560000 43.080000 ;
        RECT  9.330000 42.940000  9.630000 43.010000 ;
        RECT  9.400000 42.870000  9.700000 42.940000 ;
        RECT  9.470000 42.800000  9.770000 42.870000 ;
        RECT  9.540000 42.730000  9.840000 42.800000 ;
        RECT  9.610000 42.660000  9.910000 42.730000 ;
        RECT  9.680000 42.590000  9.980000 42.660000 ;
        RECT  9.750000 42.520000 10.050000 42.590000 ;
        RECT  9.820000 42.450000 10.120000 42.520000 ;
        RECT  9.890000 42.380000 10.190000 42.450000 ;
        RECT  9.960000 42.310000 10.260000 42.380000 ;
        RECT 10.030000 42.240000 10.330000 42.310000 ;
        RECT 10.100000 42.170000 10.400000 42.240000 ;
        RECT 10.170000 42.100000 10.470000 42.170000 ;
        RECT 10.240000 42.030000 10.540000 42.100000 ;
        RECT 10.310000 41.960000 10.610000 42.030000 ;
        RECT 10.380000 41.890000 10.680000 41.960000 ;
        RECT 10.450000 41.820000 10.750000 41.890000 ;
        RECT 10.520000 41.750000 10.820000 41.820000 ;
        RECT 10.590000 41.680000 10.890000 41.750000 ;
        RECT 10.660000 41.610000 10.960000 41.680000 ;
        RECT 10.730000 41.540000 11.030000 41.610000 ;
        RECT 10.800000 41.470000 11.100000 41.540000 ;
        RECT 10.870000 41.400000 11.170000 41.470000 ;
        RECT 10.940000 41.330000 11.240000 41.400000 ;
        RECT 11.010000 41.260000 11.310000 41.330000 ;
        RECT 11.080000 41.190000 11.380000 41.260000 ;
        RECT 11.150000 41.120000 11.450000 41.190000 ;
        RECT 11.220000 41.050000 11.520000 41.120000 ;
        RECT 11.290000 40.980000 11.590000 41.050000 ;
        RECT 11.360000 40.910000 11.660000 40.980000 ;
        RECT 11.430000 40.840000 11.730000 40.910000 ;
        RECT 11.500000 40.770000 11.800000 40.840000 ;
        RECT 11.570000 40.700000 11.870000 40.770000 ;
        RECT 11.640000 40.630000 11.940000 40.700000 ;
        RECT 11.710000 40.560000 12.010000 40.630000 ;
        RECT 11.780000 40.490000 12.080000 40.560000 ;
        RECT 11.850000 40.420000 12.150000 40.490000 ;
        RECT 11.920000 40.350000 12.220000 40.420000 ;
        RECT 11.990000 40.280000 12.290000 40.350000 ;
        RECT 12.060000 40.210000 12.360000 40.280000 ;
        RECT 12.130000 40.140000 12.430000 40.210000 ;
        RECT 12.200000 40.070000 12.500000 40.140000 ;
        RECT 12.270000 40.000000 12.570000 40.070000 ;
        RECT 12.340000 39.930000 12.640000 40.000000 ;
        RECT 12.410000 39.860000 12.710000 39.930000 ;
        RECT 12.480000 39.790000 12.780000 39.860000 ;
        RECT 12.550000 39.720000 12.850000 39.790000 ;
        RECT 12.620000 39.650000 12.920000 39.720000 ;
        RECT 12.690000 39.580000 12.990000 39.650000 ;
        RECT 12.755000  0.000000 13.015000  5.240000 ;
        RECT 12.755000  5.240000 13.015000  5.295000 ;
        RECT 12.755000  5.295000 13.070000  5.350000 ;
        RECT 12.760000 39.510000 13.060000 39.580000 ;
        RECT 12.825000  5.350000 13.125000  5.420000 ;
        RECT 12.830000 39.440000 13.130000 39.510000 ;
        RECT 12.895000  5.420000 13.195000  5.490000 ;
        RECT 12.900000 39.370000 13.200000 39.440000 ;
        RECT 12.965000  5.490000 13.265000  5.560000 ;
        RECT 12.970000 39.300000 13.270000 39.370000 ;
        RECT 13.035000  5.560000 13.335000  5.630000 ;
        RECT 13.040000 39.230000 13.340000 39.300000 ;
        RECT 13.105000  5.630000 13.405000  5.700000 ;
        RECT 13.110000 39.160000 13.410000 39.230000 ;
        RECT 13.175000  5.700000 13.475000  5.770000 ;
        RECT 13.180000 39.090000 13.480000 39.160000 ;
        RECT 13.245000  5.770000 13.545000  5.840000 ;
        RECT 13.250000 39.020000 13.550000 39.090000 ;
        RECT 13.315000  5.840000 13.615000  5.910000 ;
        RECT 13.320000 38.950000 13.620000 39.020000 ;
        RECT 13.385000  5.910000 13.685000  5.980000 ;
        RECT 13.390000 38.880000 13.690000 38.950000 ;
        RECT 13.455000  5.980000 13.755000  6.050000 ;
        RECT 13.460000 38.810000 13.760000 38.880000 ;
        RECT 13.525000  6.050000 13.825000  6.120000 ;
        RECT 13.530000 38.740000 13.830000 38.810000 ;
        RECT 13.595000  6.120000 13.895000  6.190000 ;
        RECT 13.600000 38.670000 13.900000 38.740000 ;
        RECT 13.665000  6.190000 13.965000  6.260000 ;
        RECT 13.670000 38.600000 13.970000 38.670000 ;
        RECT 13.735000  6.260000 14.035000  6.330000 ;
        RECT 13.740000 38.530000 14.040000 38.600000 ;
        RECT 13.805000  6.330000 14.105000  6.400000 ;
        RECT 13.810000 38.460000 14.110000 38.530000 ;
        RECT 13.860000  6.400000 14.175000  6.455000 ;
        RECT 13.880000 38.390000 14.180000 38.460000 ;
        RECT 13.915000  6.455000 14.230000  6.510000 ;
        RECT 13.950000 38.320000 14.250000 38.390000 ;
        RECT 13.970000  6.510000 14.230000  6.565000 ;
        RECT 13.970000  6.565000 14.230000 18.115000 ;
        RECT 13.970000 18.115000 14.230000 18.170000 ;
        RECT 13.970000 18.170000 14.285000 18.225000 ;
        RECT 14.020000 38.250000 14.320000 38.320000 ;
        RECT 14.040000 18.225000 14.340000 18.295000 ;
        RECT 14.090000 38.180000 14.390000 38.250000 ;
        RECT 14.110000 18.295000 14.410000 18.365000 ;
        RECT 14.160000 38.110000 14.460000 38.180000 ;
        RECT 14.180000 18.365000 14.480000 18.435000 ;
        RECT 14.230000 38.040000 14.530000 38.110000 ;
        RECT 14.250000 18.435000 14.550000 18.505000 ;
        RECT 14.300000 37.970000 14.600000 38.040000 ;
        RECT 14.320000 18.505000 14.620000 18.575000 ;
        RECT 14.370000 37.900000 14.670000 37.970000 ;
        RECT 14.390000 18.575000 14.690000 18.645000 ;
        RECT 14.440000 37.830000 14.740000 37.900000 ;
        RECT 14.460000 18.645000 14.760000 18.715000 ;
        RECT 14.510000 37.760000 14.810000 37.830000 ;
        RECT 14.530000 18.715000 14.830000 18.785000 ;
        RECT 14.580000 37.690000 14.880000 37.760000 ;
        RECT 14.600000 18.785000 14.900000 18.855000 ;
        RECT 14.650000 37.620000 14.950000 37.690000 ;
        RECT 14.670000 18.855000 14.970000 18.925000 ;
        RECT 14.720000 37.550000 15.020000 37.620000 ;
        RECT 14.740000 18.925000 15.040000 18.995000 ;
        RECT 14.790000 37.480000 15.090000 37.550000 ;
        RECT 14.810000 18.995000 15.110000 19.065000 ;
        RECT 14.860000 37.410000 15.160000 37.480000 ;
        RECT 14.880000 19.065000 15.180000 19.135000 ;
        RECT 14.915000 37.355000 15.230000 37.410000 ;
        RECT 14.950000 19.135000 15.250000 19.205000 ;
        RECT 14.970000 31.960000 15.285000 32.015000 ;
        RECT 14.970000 32.015000 15.230000 32.070000 ;
        RECT 14.970000 32.070000 15.230000 37.300000 ;
        RECT 14.970000 37.300000 15.230000 37.355000 ;
        RECT 14.995000 31.935000 15.340000 31.960000 ;
        RECT 15.020000 19.205000 15.320000 19.275000 ;
        RECT 15.065000 31.865000 15.365000 31.935000 ;
        RECT 15.090000 19.275000 15.390000 19.345000 ;
        RECT 15.135000 31.795000 15.435000 31.865000 ;
        RECT 15.160000 19.345000 15.460000 19.415000 ;
        RECT 15.205000 31.725000 15.505000 31.795000 ;
        RECT 15.230000 19.415000 15.530000 19.485000 ;
        RECT 15.275000 19.485000 15.600000 19.530000 ;
        RECT 15.275000 31.655000 15.575000 31.725000 ;
        RECT 15.330000 19.530000 15.645000 19.585000 ;
        RECT 15.330000 31.600000 15.645000 31.655000 ;
        RECT 15.385000 19.585000 15.645000 19.640000 ;
        RECT 15.385000 19.640000 15.645000 31.545000 ;
        RECT 15.385000 31.545000 15.645000 31.600000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580000 0.000000 78.910000 176.480000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.250000 43.835000 11.565000 43.890000 ;
        RECT 11.250000 43.890000 11.510000 43.945000 ;
        RECT 11.250000 43.945000 11.510000 47.275000 ;
        RECT 11.250000 47.275000 11.510000 47.330000 ;
        RECT 11.250000 47.330000 11.565000 47.385000 ;
        RECT 11.270000 43.815000 11.620000 43.835000 ;
        RECT 11.320000 47.385000 11.620000 47.455000 ;
        RECT 11.340000 43.745000 11.640000 43.815000 ;
        RECT 11.390000 47.455000 11.690000 47.525000 ;
        RECT 11.410000 43.675000 11.710000 43.745000 ;
        RECT 11.460000 47.525000 11.760000 47.595000 ;
        RECT 11.480000 43.605000 11.780000 43.675000 ;
        RECT 11.530000 47.595000 11.830000 47.665000 ;
        RECT 11.550000 43.535000 11.850000 43.605000 ;
        RECT 11.600000 47.665000 11.900000 47.735000 ;
        RECT 11.620000 43.465000 11.920000 43.535000 ;
        RECT 11.670000 47.735000 11.970000 47.805000 ;
        RECT 11.680000 47.805000 12.040000 47.815000 ;
        RECT 11.690000 43.395000 11.990000 43.465000 ;
        RECT 11.750000 47.815000 13.850000 47.885000 ;
        RECT 11.760000 43.325000 12.060000 43.395000 ;
        RECT 11.820000 47.885000 13.920000 47.955000 ;
        RECT 11.830000 43.255000 12.130000 43.325000 ;
        RECT 11.890000 47.955000 13.990000 48.025000 ;
        RECT 11.900000 43.185000 12.200000 43.255000 ;
        RECT 11.940000 48.025000 14.060000 48.075000 ;
        RECT 11.970000 43.115000 12.270000 43.185000 ;
        RECT 12.040000 43.045000 12.340000 43.115000 ;
        RECT 12.110000 42.975000 12.410000 43.045000 ;
        RECT 12.180000 42.905000 12.480000 42.975000 ;
        RECT 12.250000 42.835000 12.550000 42.905000 ;
        RECT 12.320000 42.765000 12.620000 42.835000 ;
        RECT 12.390000 42.695000 12.690000 42.765000 ;
        RECT 12.460000 42.625000 12.760000 42.695000 ;
        RECT 12.530000 42.555000 12.830000 42.625000 ;
        RECT 12.600000 42.485000 12.900000 42.555000 ;
        RECT 12.670000 42.415000 12.970000 42.485000 ;
        RECT 12.740000 42.345000 13.040000 42.415000 ;
        RECT 12.810000 42.275000 13.110000 42.345000 ;
        RECT 12.880000 42.205000 13.180000 42.275000 ;
        RECT 12.950000 42.135000 13.250000 42.205000 ;
        RECT 13.020000 42.065000 13.320000 42.135000 ;
        RECT 13.090000 41.995000 13.390000 42.065000 ;
        RECT 13.160000 41.925000 13.460000 41.995000 ;
        RECT 13.230000 41.855000 13.530000 41.925000 ;
        RECT 13.300000 41.785000 13.600000 41.855000 ;
        RECT 13.370000 41.715000 13.670000 41.785000 ;
        RECT 13.440000 41.645000 13.740000 41.715000 ;
        RECT 13.510000 41.575000 13.810000 41.645000 ;
        RECT 13.565000 41.520000 13.880000 41.575000 ;
        RECT 13.620000 40.430000 13.935000 40.485000 ;
        RECT 13.620000 40.485000 13.880000 40.540000 ;
        RECT 13.620000 40.540000 13.880000 41.465000 ;
        RECT 13.620000 41.465000 13.880000 41.520000 ;
        RECT 13.640000 40.410000 13.990000 40.430000 ;
        RECT 13.710000 40.340000 14.010000 40.410000 ;
        RECT 13.780000 40.270000 14.080000 40.340000 ;
        RECT 13.810000 48.075000 14.110000 48.145000 ;
        RECT 13.850000 40.200000 14.150000 40.270000 ;
        RECT 13.880000 48.145000 14.180000 48.215000 ;
        RECT 13.920000 40.130000 14.220000 40.200000 ;
        RECT 13.950000 48.215000 14.250000 48.285000 ;
        RECT 13.990000 40.060000 14.290000 40.130000 ;
        RECT 14.020000 48.285000 14.320000 48.355000 ;
        RECT 14.060000 39.990000 14.360000 40.060000 ;
        RECT 14.090000 48.355000 14.390000 48.425000 ;
        RECT 14.130000 39.920000 14.430000 39.990000 ;
        RECT 14.160000 48.425000 14.460000 48.495000 ;
        RECT 14.180000 39.870000 15.420000 39.920000 ;
        RECT 14.195000 58.050000 14.835000 58.310000 ;
        RECT 14.210000 58.035000 14.820000 58.050000 ;
        RECT 14.230000 48.495000 14.530000 48.565000 ;
        RECT 14.240000 48.565000 14.600000 48.575000 ;
        RECT 14.250000 39.800000 15.470000 39.870000 ;
        RECT 14.280000 57.965000 14.750000 58.035000 ;
        RECT 14.295000 48.575000 14.610000 48.630000 ;
        RECT 14.320000 39.730000 15.540000 39.800000 ;
        RECT 14.350000 48.630000 14.610000 48.685000 ;
        RECT 14.350000 48.685000 14.610000 57.825000 ;
        RECT 14.350000 57.825000 14.610000 57.860000 ;
        RECT 14.350000 57.860000 14.645000 57.895000 ;
        RECT 14.350000 57.895000 14.680000 57.965000 ;
        RECT 14.390000 39.660000 15.610000 39.730000 ;
        RECT 15.365000 39.605000 15.680000 39.660000 ;
        RECT 15.435000 39.535000 15.735000 39.605000 ;
        RECT 15.505000 39.465000 15.805000 39.535000 ;
        RECT 15.575000 39.395000 15.875000 39.465000 ;
        RECT 15.645000 39.325000 15.945000 39.395000 ;
        RECT 15.715000 39.255000 16.015000 39.325000 ;
        RECT 15.785000 39.185000 16.085000 39.255000 ;
        RECT 15.855000 39.115000 16.155000 39.185000 ;
        RECT 15.925000 39.045000 16.225000 39.115000 ;
        RECT 15.995000 38.975000 16.295000 39.045000 ;
        RECT 16.065000 38.905000 16.365000 38.975000 ;
        RECT 16.135000 38.835000 16.435000 38.905000 ;
        RECT 16.205000 38.765000 16.505000 38.835000 ;
        RECT 16.275000 38.695000 16.575000 38.765000 ;
        RECT 16.310000  0.000000 16.570000  2.210000 ;
        RECT 16.310000  2.210000 16.570000  2.265000 ;
        RECT 16.310000  2.265000 16.625000  2.320000 ;
        RECT 16.345000 38.625000 16.645000 38.695000 ;
        RECT 16.365000 31.560000 16.680000 31.615000 ;
        RECT 16.365000 31.615000 16.625000 31.670000 ;
        RECT 16.365000 31.670000 16.625000 34.210000 ;
        RECT 16.365000 34.210000 16.625000 34.265000 ;
        RECT 16.365000 34.265000 16.680000 34.320000 ;
        RECT 16.370000 31.555000 16.735000 31.560000 ;
        RECT 16.380000  2.320000 16.680000  2.390000 ;
        RECT 16.415000 38.555000 16.715000 38.625000 ;
        RECT 16.435000 31.490000 16.740000 31.555000 ;
        RECT 16.435000 34.320000 16.735000 34.390000 ;
        RECT 16.450000  2.390000 16.750000  2.460000 ;
        RECT 16.485000 38.485000 16.785000 38.555000 ;
        RECT 16.500000 31.425000 16.805000 31.490000 ;
        RECT 16.505000 34.390000 16.805000 34.460000 ;
        RECT 16.520000  2.460000 16.820000  2.530000 ;
        RECT 16.555000 31.370000 16.870000 31.425000 ;
        RECT 16.555000 38.415000 16.855000 38.485000 ;
        RECT 16.575000 34.460000 16.875000 34.530000 ;
        RECT 16.590000  2.530000 16.890000  2.600000 ;
        RECT 16.610000  7.160000 16.925000  7.215000 ;
        RECT 16.610000  7.215000 16.870000  7.270000 ;
        RECT 16.610000  7.270000 16.870000 11.540000 ;
        RECT 16.610000 12.475000 16.870000 31.315000 ;
        RECT 16.610000 31.315000 16.870000 31.370000 ;
        RECT 16.615000 12.470000 16.870000 12.475000 ;
        RECT 16.625000 38.345000 16.925000 38.415000 ;
        RECT 16.635000  7.135000 16.980000  7.160000 ;
        RECT 16.645000 34.530000 16.945000 34.600000 ;
        RECT 16.655000 11.540000 16.870000 11.585000 ;
        RECT 16.660000  2.600000 16.960000  2.670000 ;
        RECT 16.660000 12.425000 16.870000 12.470000 ;
        RECT 16.695000 38.275000 16.995000 38.345000 ;
        RECT 16.700000 11.585000 16.870000 11.630000 ;
        RECT 16.705000  7.065000 17.005000  7.135000 ;
        RECT 16.705000 11.630000 16.870000 11.635000 ;
        RECT 16.705000 11.635000 16.870000 12.380000 ;
        RECT 16.705000 12.380000 16.870000 12.425000 ;
        RECT 16.715000 34.600000 17.015000 34.670000 ;
        RECT 16.730000  2.670000 17.030000  2.740000 ;
        RECT 16.765000 38.205000 17.065000 38.275000 ;
        RECT 16.775000  6.995000 17.075000  7.065000 ;
        RECT 16.785000 34.670000 17.085000 34.740000 ;
        RECT 16.800000  2.740000 17.100000  2.810000 ;
        RECT 16.835000 38.135000 17.135000 38.205000 ;
        RECT 16.845000  6.925000 17.145000  6.995000 ;
        RECT 16.855000 34.740000 17.155000 34.810000 ;
        RECT 16.870000  2.810000 17.170000  2.880000 ;
        RECT 16.905000 38.065000 17.205000 38.135000 ;
        RECT 16.915000  6.855000 17.215000  6.925000 ;
        RECT 16.925000 34.810000 17.225000 34.880000 ;
        RECT 16.940000  2.880000 17.240000  2.950000 ;
        RECT 16.975000 37.995000 17.275000 38.065000 ;
        RECT 16.985000  2.950000 17.310000  2.995000 ;
        RECT 16.985000  6.785000 17.285000  6.855000 ;
        RECT 16.995000 34.880000 17.295000 34.950000 ;
        RECT 17.040000  2.995000 17.355000  3.050000 ;
        RECT 17.040000  6.730000 17.355000  6.785000 ;
        RECT 17.045000 37.925000 17.345000 37.995000 ;
        RECT 17.065000 34.950000 17.365000 35.020000 ;
        RECT 17.095000  3.050000 17.355000  3.105000 ;
        RECT 17.095000  3.105000 17.355000  6.675000 ;
        RECT 17.095000  6.675000 17.355000  6.730000 ;
        RECT 17.115000 37.855000 17.415000 37.925000 ;
        RECT 17.135000 35.020000 17.435000 35.090000 ;
        RECT 17.185000 37.785000 17.485000 37.855000 ;
        RECT 17.205000 35.090000 17.505000 35.160000 ;
        RECT 17.255000 37.715000 17.555000 37.785000 ;
        RECT 17.275000 35.160000 17.575000 35.230000 ;
        RECT 17.325000 37.645000 17.625000 37.715000 ;
        RECT 17.345000 35.230000 17.645000 35.300000 ;
        RECT 17.395000 37.575000 17.695000 37.645000 ;
        RECT 17.415000 35.300000 17.715000 35.370000 ;
        RECT 17.465000 35.370000 17.785000 35.420000 ;
        RECT 17.465000 37.505000 17.765000 37.575000 ;
        RECT 17.520000 35.420000 17.835000 35.475000 ;
        RECT 17.520000 37.450000 17.835000 37.505000 ;
        RECT 17.575000 35.475000 17.835000 35.530000 ;
        RECT 17.575000 35.530000 17.835000 37.395000 ;
        RECT 17.575000 37.395000 17.835000 37.450000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815000 0.000000 32.075000 3.965000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600000 0.000000 26.860000 1.695000 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420000 0.000000 5.650000 4.375000 ;
        RECT 5.420000 4.375000 5.650000 4.425000 ;
        RECT 5.420000 4.425000 5.700000 4.475000 ;
        RECT 5.490000 4.475000 5.750000 4.545000 ;
        RECT 5.560000 4.545000 5.820000 4.615000 ;
        RECT 5.630000 4.615000 5.890000 4.685000 ;
        RECT 5.700000 4.685000 5.960000 4.755000 ;
        RECT 5.770000 4.755000 6.030000 4.825000 ;
        RECT 5.840000 4.825000 6.100000 4.895000 ;
        RECT 5.910000 4.895000 6.170000 4.965000 ;
        RECT 5.910000 6.425000 6.550000 6.685000 ;
        RECT 5.980000 4.965000 6.240000 5.035000 ;
        RECT 6.050000 5.035000 6.310000 5.105000 ;
        RECT 6.120000 5.105000 6.380000 5.175000 ;
        RECT 6.180000 6.390000 6.550000 6.425000 ;
        RECT 6.190000 5.175000 6.450000 5.245000 ;
        RECT 6.220000 5.245000 6.520000 5.275000 ;
        RECT 6.250000 6.320000 6.550000 6.390000 ;
        RECT 6.270000 5.275000 6.550000 5.325000 ;
        RECT 6.320000 5.325000 6.550000 5.375000 ;
        RECT 6.320000 5.375000 6.550000 6.250000 ;
        RECT 6.320000 6.250000 6.550000 6.320000 ;
    END
  END IB_MODE_SEL
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  303.1200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240000 0.000000 79.570000 176.480000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245000 0.000000 45.505000 4.980000 ;
        RECT 45.245000 4.980000 45.505000 5.035000 ;
        RECT 45.245000 5.035000 45.560000 5.090000 ;
        RECT 45.315000 5.090000 45.615000 5.160000 ;
        RECT 45.385000 5.160000 45.685000 5.230000 ;
        RECT 45.455000 5.230000 45.755000 5.300000 ;
        RECT 45.525000 5.300000 45.825000 5.370000 ;
        RECT 45.595000 5.370000 45.895000 5.440000 ;
        RECT 45.665000 5.440000 45.965000 5.510000 ;
        RECT 45.735000 5.510000 46.035000 5.580000 ;
        RECT 45.745000 5.580000 46.105000 5.590000 ;
        RECT 45.800000 5.590000 46.115000 5.645000 ;
        RECT 45.855000 5.645000 46.115000 5.700000 ;
        RECT 45.855000 5.700000 46.115000 6.780000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  291.9480 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400000   0.000000 1.020000 178.235000 ;
        RECT 0.400000 178.235000 1.020000 178.360000 ;
        RECT 0.400000 178.360000 1.145000 178.485000 ;
        RECT 0.550000 178.485000 1.270000 178.635000 ;
        RECT 0.700000 178.635000 1.420000 178.785000 ;
        RECT 0.850000 178.785000 1.570000 178.935000 ;
        RECT 1.000000 178.935000 1.720000 179.085000 ;
        RECT 1.150000 179.085000 1.870000 179.235000 ;
        RECT 1.300000 179.235000 2.020000 179.385000 ;
        RECT 1.450000 179.385000 2.170000 179.535000 ;
        RECT 1.600000 179.535000 2.320000 179.685000 ;
        RECT 1.750000 179.685000 2.470000 179.835000 ;
        RECT 1.900000 179.835000 2.620000 179.985000 ;
        RECT 2.050000 179.985000 2.770000 180.135000 ;
        RECT 2.200000 180.135000 2.920000 180.285000 ;
        RECT 2.350000 180.285000 3.070000 180.435000 ;
        RECT 2.355000 180.435000 3.220000 180.440000 ;
        RECT 2.505000 180.440000 4.565000 180.590000 ;
        RECT 2.655000 180.590000 4.565000 180.740000 ;
        RECT 2.805000 180.740000 4.565000 180.890000 ;
        RECT 2.955000 180.890000 4.565000 181.040000 ;
        RECT 3.085000 181.040000 4.565000 181.170000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAGATEAREA  1.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375000  0.000000 3.605000  4.375000 ;
        RECT 3.375000  4.375000 3.605000  4.425000 ;
        RECT 3.375000  4.425000 3.655000  4.475000 ;
        RECT 3.445000  4.475000 3.705000  4.545000 ;
        RECT 3.515000  4.545000 3.775000  4.615000 ;
        RECT 3.585000  4.615000 3.845000  4.685000 ;
        RECT 3.655000  4.685000 3.915000  4.755000 ;
        RECT 3.725000  4.755000 3.985000  4.825000 ;
        RECT 3.770000  4.825000 4.055000  4.870000 ;
        RECT 3.840000  4.870000 5.225000  4.940000 ;
        RECT 3.910000  4.940000 5.295000  5.010000 ;
        RECT 3.980000  5.010000 5.365000  5.080000 ;
        RECT 4.000000  5.080000 5.435000  5.100000 ;
        RECT 5.195000  5.100000 5.455000  5.170000 ;
        RECT 5.265000  5.170000 5.525000  5.240000 ;
        RECT 5.300000  5.240000 5.595000  5.275000 ;
        RECT 5.350000  5.275000 5.630000  5.325000 ;
        RECT 5.400000  5.325000 5.630000  5.375000 ;
        RECT 5.400000  5.375000 5.630000  8.250000 ;
        RECT 5.400000  8.250000 5.630000  8.300000 ;
        RECT 5.400000  8.300000 5.680000  8.350000 ;
        RECT 5.470000  8.350000 5.730000  8.420000 ;
        RECT 5.540000  8.420000 5.800000  8.490000 ;
        RECT 5.610000  8.490000 5.870000  8.560000 ;
        RECT 5.680000  8.560000 5.940000  8.630000 ;
        RECT 5.750000  8.630000 6.010000  8.700000 ;
        RECT 5.820000  8.700000 6.080000  8.770000 ;
        RECT 5.890000  8.770000 6.150000  8.840000 ;
        RECT 5.960000  8.840000 6.220000  8.910000 ;
        RECT 5.965000 42.985000 6.225000 43.625000 ;
        RECT 5.970000 42.980000 6.220000 42.985000 ;
        RECT 5.975000 39.420000 6.255000 39.470000 ;
        RECT 5.975000 39.470000 6.205000 39.520000 ;
        RECT 5.975000 39.520000 6.205000 42.965000 ;
        RECT 5.975000 42.965000 6.205000 42.970000 ;
        RECT 5.975000 42.970000 6.210000 42.975000 ;
        RECT 5.975000 42.975000 6.215000 42.980000 ;
        RECT 5.985000 39.410000 6.305000 39.420000 ;
        RECT 6.030000  8.910000 6.290000  8.980000 ;
        RECT 6.055000 39.340000 6.315000 39.410000 ;
        RECT 6.100000  8.980000 6.360000  9.050000 ;
        RECT 6.125000 39.270000 6.385000 39.340000 ;
        RECT 6.170000  9.050000 6.430000  9.120000 ;
        RECT 6.195000 39.200000 6.455000 39.270000 ;
        RECT 6.240000  9.120000 6.500000  9.190000 ;
        RECT 6.265000 39.130000 6.525000 39.200000 ;
        RECT 6.310000  9.190000 6.570000  9.260000 ;
        RECT 6.335000 39.060000 6.595000 39.130000 ;
        RECT 6.380000  9.260000 6.640000  9.330000 ;
        RECT 6.405000 38.990000 6.665000 39.060000 ;
        RECT 6.450000  9.330000 6.710000  9.400000 ;
        RECT 6.475000  9.400000 6.780000  9.425000 ;
        RECT 6.475000 38.920000 6.735000 38.990000 ;
        RECT 6.525000  9.425000 6.805000  9.475000 ;
        RECT 6.525000 38.870000 6.805000 38.920000 ;
        RECT 6.575000  9.475000 6.805000  9.525000 ;
        RECT 6.575000  9.525000 6.805000 38.820000 ;
        RECT 6.575000 38.820000 6.805000 38.870000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355000  0.000000 22.615000  6.315000 ;
        RECT 22.355000  6.315000 22.615000  6.370000 ;
        RECT 22.355000  6.370000 22.670000  6.425000 ;
        RECT 22.425000  6.425000 22.725000  6.495000 ;
        RECT 22.495000  6.495000 22.795000  6.565000 ;
        RECT 22.565000  6.565000 22.865000  6.635000 ;
        RECT 22.635000  6.635000 22.935000  6.705000 ;
        RECT 22.655000  6.705000 23.005000  6.725000 ;
        RECT 22.710000  6.725000 23.025000  6.780000 ;
        RECT 22.765000  6.780000 23.025000  6.835000 ;
        RECT 22.765000  6.835000 23.025000 14.375000 ;
        RECT 22.765000 14.375000 23.025000 14.430000 ;
        RECT 22.765000 14.430000 23.080000 14.485000 ;
        RECT 22.835000 14.485000 23.135000 14.555000 ;
        RECT 22.905000 14.555000 23.205000 14.625000 ;
        RECT 22.975000 14.625000 23.275000 14.695000 ;
        RECT 23.045000 14.695000 23.345000 14.765000 ;
        RECT 23.095000 38.695000 23.735000 38.955000 ;
        RECT 23.115000 14.765000 23.415000 14.835000 ;
        RECT 23.185000 14.835000 23.485000 14.905000 ;
        RECT 23.255000 14.905000 23.555000 14.975000 ;
        RECT 23.265000 38.625000 23.735000 38.695000 ;
        RECT 23.325000 14.975000 23.625000 15.045000 ;
        RECT 23.335000 38.555000 23.735000 38.625000 ;
        RECT 23.395000 15.045000 23.695000 15.115000 ;
        RECT 23.405000 38.485000 23.735000 38.555000 ;
        RECT 23.465000 15.115000 23.765000 15.185000 ;
        RECT 23.475000 25.180000 23.790000 25.235000 ;
        RECT 23.475000 25.235000 23.735000 25.290000 ;
        RECT 23.475000 25.290000 23.735000 38.415000 ;
        RECT 23.475000 38.415000 23.735000 38.485000 ;
        RECT 23.510000 25.145000 23.845000 25.180000 ;
        RECT 23.535000 15.185000 23.835000 15.255000 ;
        RECT 23.545000 15.255000 23.905000 15.265000 ;
        RECT 23.545000 25.110000 23.880000 25.145000 ;
        RECT 23.600000 15.265000 23.915000 15.320000 ;
        RECT 23.600000 25.055000 23.915000 25.110000 ;
        RECT 23.655000 15.320000 23.915000 15.375000 ;
        RECT 23.655000 15.375000 23.915000 25.000000 ;
        RECT 23.655000 25.000000 23.915000 25.055000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  216.1550 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.115000 125.470000 53.655000 147.015000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  3.812250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280000 0.000000 76.920000 1.625000 ;
        RECT 76.280000 1.625000 76.920000 1.695000 ;
        RECT 76.280000 1.695000 76.990000 1.765000 ;
        RECT 76.280000 1.765000 77.060000 1.835000 ;
        RECT 76.280000 1.835000 77.130000 1.905000 ;
        RECT 76.280000 1.905000 77.200000 1.975000 ;
        RECT 76.280000 1.975000 77.270000 2.045000 ;
        RECT 76.280000 2.045000 77.340000 2.055000 ;
        RECT 76.350000 2.055000 77.350000 2.125000 ;
        RECT 76.420000 2.125000 77.420000 2.195000 ;
        RECT 76.490000 2.195000 77.490000 2.265000 ;
        RECT 76.560000 2.265000 77.560000 2.335000 ;
        RECT 76.630000 2.335000 77.630000 2.405000 ;
        RECT 76.700000 2.405000 77.700000 2.475000 ;
        RECT 76.770000 2.475000 77.770000 2.545000 ;
        RECT 76.820000 2.545000 77.840000 2.595000 ;
        RECT 76.890000 2.595000 77.890000 2.665000 ;
        RECT 76.960000 2.665000 77.890000 2.735000 ;
        RECT 77.030000 2.735000 77.890000 2.805000 ;
        RECT 77.100000 2.805000 77.890000 2.875000 ;
        RECT 77.150000 2.875000 77.890000 2.925000 ;
        RECT 77.150000 2.925000 77.890000 5.235000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  2.618000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275000 0.000000 68.925000 3.960000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  4.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.600000  7.425000 60.560000   7.575000 ;
        RECT 59.600000  7.575000 60.410000   7.725000 ;
        RECT 59.600000  7.725000 60.385000   7.750000 ;
        RECT 59.600000  7.750000 60.385000  10.610000 ;
        RECT 59.600000 10.610000 60.385000  10.760000 ;
        RECT 59.600000 10.760000 60.535000  10.910000 ;
        RECT 59.600000 10.910000 60.685000  10.935000 ;
        RECT 59.655000  7.370000 60.710000   7.425000 ;
        RECT 59.750000 10.935000 60.710000  11.085000 ;
        RECT 59.805000  7.220000 60.765000   7.370000 ;
        RECT 59.900000 11.085000 60.860000  11.235000 ;
        RECT 59.955000  7.070000 60.915000   7.220000 ;
        RECT 59.985000  7.040000 63.890000   7.070000 ;
        RECT 60.050000 11.235000 61.010000  11.385000 ;
        RECT 60.135000  6.890000 63.890000   7.040000 ;
        RECT 60.200000 11.385000 61.160000  11.535000 ;
        RECT 60.285000  6.740000 63.890000   6.890000 ;
        RECT 60.350000 11.535000 61.310000  11.685000 ;
        RECT 60.435000  6.590000 63.890000   6.740000 ;
        RECT 60.500000 11.685000 61.460000  11.835000 ;
        RECT 60.585000  6.440000 63.890000   6.590000 ;
        RECT 60.610000 19.065000 61.570000  19.215000 ;
        RECT 60.610000 19.215000 61.420000  19.365000 ;
        RECT 60.610000 19.365000 61.395000  19.390000 ;
        RECT 60.610000 19.390000 61.395000  47.360000 ;
        RECT 60.650000 11.835000 61.610000  11.985000 ;
        RECT 60.690000 18.985000 61.720000  19.065000 ;
        RECT 60.735000  6.290000 63.890000   6.440000 ;
        RECT 60.800000 11.985000 61.760000  12.135000 ;
        RECT 60.840000 18.835000 61.800000  18.985000 ;
        RECT 60.950000 12.135000 61.910000  12.285000 ;
        RECT 60.990000 18.685000 61.950000  18.835000 ;
        RECT 61.100000 12.285000 62.060000  12.435000 ;
        RECT 61.140000 12.435000 62.210000  12.475000 ;
        RECT 61.140000 18.535000 62.100000  18.685000 ;
        RECT 61.170000 18.505000 62.250000  18.535000 ;
        RECT 61.290000 12.475000 62.250000  12.625000 ;
        RECT 61.320000 18.355000 62.250000  18.505000 ;
        RECT 61.440000 12.625000 62.250000  12.775000 ;
        RECT 61.470000 12.775000 62.250000  12.805000 ;
        RECT 61.470000 12.805000 62.250000  18.205000 ;
        RECT 61.470000 18.205000 62.250000  18.355000 ;
        RECT 61.710000 35.760000 63.070000  35.910000 ;
        RECT 61.710000 35.910000 62.920000  36.060000 ;
        RECT 61.710000 36.060000 62.780000  36.200000 ;
        RECT 61.710000 36.200000 62.780000  73.005000 ;
        RECT 61.710000 73.005000 62.780000  73.155000 ;
        RECT 61.710000 73.155000 62.930000  73.305000 ;
        RECT 61.710000 73.305000 63.080000  73.455000 ;
        RECT 61.710000 73.455000 63.230000  73.605000 ;
        RECT 61.710000 73.605000 63.380000  73.755000 ;
        RECT 61.710000 73.755000 63.530000  73.905000 ;
        RECT 61.710000 73.905000 63.680000  74.055000 ;
        RECT 61.710000 74.055000 63.830000  74.185000 ;
        RECT 61.735000 35.735000 63.220000  35.760000 ;
        RECT 61.750000 74.185000 63.960000  74.225000 ;
        RECT 61.790000 74.225000 64.000000  74.265000 ;
        RECT 61.885000 35.585000 63.245000  35.735000 ;
        RECT 61.940000 74.265000 68.555000  74.415000 ;
        RECT 62.035000 35.435000 63.395000  35.585000 ;
        RECT 62.090000 74.415000 68.705000  74.565000 ;
        RECT 62.185000 35.285000 63.545000  35.435000 ;
        RECT 62.220000  6.155000 63.890000   6.290000 ;
        RECT 62.235000  7.070000 63.890000   7.220000 ;
        RECT 62.240000 74.565000 68.855000  74.715000 ;
        RECT 62.325000 35.145000 63.695000  35.285000 ;
        RECT 62.370000  6.005000 63.890000   6.155000 ;
        RECT 62.385000  7.220000 63.890000   7.370000 ;
        RECT 62.390000 74.715000 69.005000  74.865000 ;
        RECT 62.475000 34.995000 63.695000  35.145000 ;
        RECT 62.520000  5.855000 63.890000   6.005000 ;
        RECT 62.535000  7.370000 63.890000   7.520000 ;
        RECT 62.540000 74.865000 69.155000  75.015000 ;
        RECT 62.625000 17.825000 63.890000  18.070000 ;
        RECT 62.625000 18.070000 63.795000  18.165000 ;
        RECT 62.625000 18.165000 63.700000  18.260000 ;
        RECT 62.625000 18.260000 63.695000  18.265000 ;
        RECT 62.625000 18.265000 63.695000  34.845000 ;
        RECT 62.625000 34.845000 63.695000  34.995000 ;
        RECT 62.630000 17.820000 63.890000  17.825000 ;
        RECT 62.670000  5.705000 63.890000   5.855000 ;
        RECT 62.685000  7.520000 63.890000   7.670000 ;
        RECT 62.690000 75.015000 69.305000  75.165000 ;
        RECT 62.725000 17.725000 63.890000  17.820000 ;
        RECT 62.820000  0.000000 63.890000   5.555000 ;
        RECT 62.820000  5.555000 63.890000   5.705000 ;
        RECT 62.820000  7.670000 63.890000   7.805000 ;
        RECT 62.820000  7.805000 63.890000  17.630000 ;
        RECT 62.820000 17.630000 63.890000  17.725000 ;
        RECT 62.840000 75.165000 69.455000  75.315000 ;
        RECT 62.860000 75.315000 69.605000  75.335000 ;
        RECT 67.870000 75.335000 69.625000  75.400000 ;
        RECT 67.935000 75.400000 69.690000  75.465000 ;
        RECT 67.940000 75.465000 69.755000  75.470000 ;
        RECT 68.090000 75.470000 69.760000  75.620000 ;
        RECT 68.240000 75.620000 69.760000  75.770000 ;
        RECT 68.390000 75.770000 69.760000  75.920000 ;
        RECT 68.540000 75.920000 69.760000  76.070000 ;
        RECT 68.690000 76.070000 69.760000  76.220000 ;
        RECT 68.690000 76.220000 69.760000 101.910000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.000000 106.585000 12.500000 118.955000 ;
        RECT 7.665000 118.955000 12.500000 119.105000 ;
        RECT 7.815000 119.105000 12.500000 119.255000 ;
        RECT 7.850000 106.565000 12.500000 106.585000 ;
        RECT 7.965000 119.255000 12.500000 119.405000 ;
        RECT 8.000000 106.415000 12.500000 106.565000 ;
        RECT 8.115000 119.405000 12.500000 119.555000 ;
        RECT 8.150000 106.265000 12.500000 106.415000 ;
        RECT 8.265000 119.555000 12.500000 119.705000 ;
        RECT 8.300000 106.115000 12.500000 106.265000 ;
        RECT 8.415000 119.705000 12.500000 119.855000 ;
        RECT 8.450000 105.965000 12.500000 106.115000 ;
        RECT 8.565000 119.855000 12.500000 120.005000 ;
        RECT 8.600000 105.815000 12.500000 105.965000 ;
        RECT 8.715000 120.005000 12.500000 120.155000 ;
        RECT 8.750000 105.665000 12.500000 105.815000 ;
        RECT 8.865000 120.155000 12.500000 120.305000 ;
        RECT 8.900000 105.515000 12.500000 105.665000 ;
        RECT 9.015000 120.305000 12.500000 120.455000 ;
        RECT 9.050000 105.365000 12.500000 105.515000 ;
        RECT 9.165000 120.455000 12.500000 120.605000 ;
        RECT 9.200000 105.215000 12.500000 105.365000 ;
        RECT 9.315000 120.605000 12.500000 120.755000 ;
        RECT 9.350000 105.065000 12.500000 105.215000 ;
        RECT 9.465000 120.755000 12.500000 120.905000 ;
        RECT 9.500000 104.915000 12.500000 105.065000 ;
        RECT 9.615000 120.905000 12.500000 121.055000 ;
        RECT 9.650000 104.765000 12.500000 104.915000 ;
        RECT 9.765000 121.055000 12.500000 121.205000 ;
        RECT 9.800000 104.615000 12.500000 104.765000 ;
        RECT 9.810000 121.205000 12.500000 121.250000 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.390000 1.185000 78.210000 1.465000 ;
        RECT 77.470000 1.125000 78.120000 1.185000 ;
        RECT 77.540000 1.055000 78.050000 1.125000 ;
        RECT 77.610000 0.000000 77.870000 0.875000 ;
        RECT 77.610000 0.875000 77.870000 0.930000 ;
        RECT 77.610000 0.930000 77.925000 0.985000 ;
        RECT 77.610000 0.985000 77.980000 1.055000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAPARTIALMETALSIDEAREA  85.19250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.230000 50.760000 76.475000 50.805000 ;
        RECT 76.230000 50.805000 76.430000 50.850000 ;
        RECT 76.230000 50.850000 76.430000 52.425000 ;
        RECT 76.230000 52.425000 76.430000 52.470000 ;
        RECT 76.230000 52.470000 76.475000 52.515000 ;
        RECT 76.280000 50.710000 76.520000 50.760000 ;
        RECT 76.300000 52.515000 76.520000 52.585000 ;
        RECT 76.350000 50.640000 76.570000 50.710000 ;
        RECT 76.370000 52.585000 76.590000 52.655000 ;
        RECT 76.420000 50.570000 76.640000 50.640000 ;
        RECT 76.440000 52.655000 76.660000 52.725000 ;
        RECT 76.490000 50.500000 76.710000 50.570000 ;
        RECT 76.510000 52.725000 76.730000 52.795000 ;
        RECT 76.560000 50.430000 76.780000 50.500000 ;
        RECT 76.580000 52.795000 76.800000 52.865000 ;
        RECT 76.630000 50.360000 76.850000 50.430000 ;
        RECT 76.650000 52.865000 76.870000 52.935000 ;
        RECT 76.700000 50.290000 76.920000 50.360000 ;
        RECT 76.720000 52.935000 76.940000 53.005000 ;
        RECT 76.770000 50.220000 76.990000 50.290000 ;
        RECT 76.790000 53.005000 77.010000 53.075000 ;
        RECT 76.825000 53.075000 77.080000 53.110000 ;
        RECT 76.840000 50.150000 77.060000 50.220000 ;
        RECT 76.870000 53.110000 77.115000 53.155000 ;
        RECT 76.900000 96.210000 77.130000 96.225000 ;
        RECT 76.910000 50.080000 77.130000 50.150000 ;
        RECT 76.915000 53.155000 77.115000 53.200000 ;
        RECT 76.915000 53.200000 77.115000 96.195000 ;
        RECT 76.915000 96.195000 77.115000 96.210000 ;
        RECT 76.980000 50.010000 77.200000 50.080000 ;
        RECT 77.050000 49.940000 77.270000 50.010000 ;
        RECT 77.120000 49.870000 77.340000 49.940000 ;
        RECT 77.190000 49.800000 77.410000 49.870000 ;
        RECT 77.260000 49.730000 77.480000 49.800000 ;
        RECT 77.330000 49.660000 77.550000 49.730000 ;
        RECT 77.400000 49.590000 77.620000 49.660000 ;
        RECT 77.470000 49.520000 77.690000 49.590000 ;
        RECT 77.540000 49.450000 77.760000 49.520000 ;
        RECT 77.610000 49.380000 77.830000 49.450000 ;
        RECT 77.680000 49.310000 77.900000 49.380000 ;
        RECT 77.750000 49.240000 77.970000 49.310000 ;
        RECT 77.820000 49.170000 78.040000 49.240000 ;
        RECT 77.890000 49.100000 78.110000 49.170000 ;
        RECT 77.960000 49.030000 78.180000 49.100000 ;
        RECT 78.030000 48.960000 78.250000 49.030000 ;
        RECT 78.100000 48.890000 78.320000 48.960000 ;
        RECT 78.170000 48.820000 78.390000 48.890000 ;
        RECT 78.240000 48.750000 78.460000 48.820000 ;
        RECT 78.310000 48.680000 78.530000 48.750000 ;
        RECT 78.380000 48.610000 78.600000 48.680000 ;
        RECT 78.450000 48.540000 78.670000 48.610000 ;
        RECT 78.520000 48.470000 78.740000 48.540000 ;
        RECT 78.590000 48.400000 78.810000 48.470000 ;
        RECT 78.615000 10.265000 78.910000 10.340000 ;
        RECT 78.615000 10.340000 78.860000 10.390000 ;
        RECT 78.615000 10.390000 78.810000 10.440000 ;
        RECT 78.615000 10.440000 78.805000 10.445000 ;
        RECT 78.615000 10.445000 78.805000 16.245000 ;
        RECT 78.615000 16.245000 78.805000 16.285000 ;
        RECT 78.615000 16.285000 78.845000 16.325000 ;
        RECT 78.620000 10.260000 78.910000 10.265000 ;
        RECT 78.660000 48.330000 78.880000 48.400000 ;
        RECT 78.665000 10.215000 78.910000 10.260000 ;
        RECT 78.685000 16.325000 78.885000 16.395000 ;
        RECT 78.705000  0.000000 78.905000  1.125000 ;
        RECT 78.705000  1.125000 78.905000  1.130000 ;
        RECT 78.705000  1.130000 78.910000  1.215000 ;
        RECT 78.710000  1.215000 78.910000  1.220000 ;
        RECT 78.710000  1.220000 78.910000 10.170000 ;
        RECT 78.710000 10.170000 78.910000 10.215000 ;
        RECT 78.730000 48.260000 78.950000 48.330000 ;
        RECT 78.755000 16.395000 78.955000 16.465000 ;
        RECT 78.800000 48.190000 79.020000 48.260000 ;
        RECT 78.825000 16.465000 79.025000 16.535000 ;
        RECT 78.870000 48.120000 79.090000 48.190000 ;
        RECT 78.895000 16.535000 79.095000 16.605000 ;
        RECT 78.940000 48.050000 79.160000 48.120000 ;
        RECT 78.965000 16.605000 79.165000 16.675000 ;
        RECT 79.010000 47.980000 79.230000 48.050000 ;
        RECT 79.035000 16.675000 79.235000 16.745000 ;
        RECT 79.080000 47.910000 79.300000 47.980000 ;
        RECT 79.105000 16.745000 79.305000 16.815000 ;
        RECT 79.150000 47.840000 79.370000 47.910000 ;
        RECT 79.175000 16.815000 79.375000 16.885000 ;
        RECT 79.220000 47.770000 79.440000 47.840000 ;
        RECT 79.240000 16.885000 79.445000 16.950000 ;
        RECT 79.270000 47.720000 79.510000 47.770000 ;
        RECT 79.280000 16.950000 79.510000 16.990000 ;
        RECT 79.320000 16.990000 79.510000 17.030000 ;
        RECT 79.320000 17.030000 79.510000 47.670000 ;
        RECT 79.320000 47.670000 79.510000 47.720000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALMETALSIDEAREA  165.2660 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715000 0.000000 79.915000 96.000000 ;
    END
  END TIE_LO_ESD
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130000 0.000000 6.390000 1.440000 ;
        RECT 6.130000 1.440000 6.390000 1.495000 ;
        RECT 6.130000 1.495000 6.445000 1.550000 ;
        RECT 6.200000 1.550000 6.500000 1.620000 ;
        RECT 6.270000 1.620000 6.570000 1.690000 ;
        RECT 6.340000 1.690000 6.640000 1.760000 ;
        RECT 6.410000 1.760000 6.710000 1.830000 ;
        RECT 6.480000 1.830000 6.780000 1.900000 ;
        RECT 6.550000 1.900000 6.850000 1.970000 ;
        RECT 6.620000 1.970000 6.920000 2.040000 ;
        RECT 6.690000 2.040000 6.990000 2.110000 ;
        RECT 6.760000 2.110000 7.060000 2.180000 ;
        RECT 6.830000 2.180000 7.130000 2.250000 ;
        RECT 6.900000 2.250000 7.200000 2.320000 ;
        RECT 6.970000 2.320000 7.270000 2.390000 ;
        RECT 7.040000 2.390000 7.340000 2.460000 ;
        RECT 7.110000 2.460000 7.410000 2.530000 ;
        RECT 7.180000 2.530000 7.480000 2.600000 ;
        RECT 7.250000 2.600000 7.550000 2.670000 ;
        RECT 7.320000 2.670000 7.620000 2.740000 ;
        RECT 7.390000 2.740000 7.690000 2.810000 ;
        RECT 7.460000 2.810000 7.760000 2.880000 ;
        RECT 7.530000 2.880000 7.830000 2.950000 ;
        RECT 7.600000 2.950000 7.900000 3.020000 ;
        RECT 7.670000 3.020000 7.970000 3.090000 ;
        RECT 7.740000 3.090000 8.040000 3.160000 ;
        RECT 7.810000 3.160000 8.110000 3.230000 ;
        RECT 7.880000 3.230000 8.180000 3.300000 ;
        RECT 7.950000 3.300000 8.250000 3.370000 ;
        RECT 8.020000 3.370000 8.320000 3.440000 ;
        RECT 8.090000 3.440000 8.390000 3.510000 ;
        RECT 8.160000 3.510000 8.460000 3.580000 ;
        RECT 8.230000 3.580000 8.530000 3.650000 ;
        RECT 8.300000 3.650000 8.600000 3.720000 ;
        RECT 8.335000 3.720000 8.670000 3.755000 ;
        RECT 8.390000 3.755000 8.705000 3.810000 ;
        RECT 8.445000 3.810000 8.705000 3.865000 ;
        RECT 8.445000 3.865000 8.705000 6.780000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 8.885000 80.000000 13.535000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 2.035000 80.000000 7.485000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 19.785000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 70.035000 80.000000 95.000000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 64.085000 80.000000 68.535000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 36.735000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 41.585000 80.000000 46.235000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 25.835000 80.000000 30.485000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 58.235000 80.000000 62.685000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 31.885000 80.000000 35.335000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.115000  95.895000 45.710000  95.955000 ;
      RECT -0.115000  95.955000  4.915000 130.220000 ;
      RECT -0.115000 131.275000  4.915000 140.050000 ;
      RECT -0.115000 140.050000  1.495000 140.150000 ;
      RECT -0.115000 145.155000  1.495000 145.210000 ;
      RECT -0.115000 145.210000  4.915000 170.090000 ;
      RECT -0.085000  93.065000  9.000000  95.255000 ;
      RECT -0.085000  95.255000 45.710000  95.895000 ;
      RECT -0.085000 130.220000  4.915000 130.225000 ;
      RECT -0.085000 130.995000  4.915000 131.275000 ;
      RECT -0.085000 170.090000  4.915000 178.645000 ;
      RECT  0.950000  18.885000  1.310000  19.055000 ;
      RECT  0.980000  21.465000  1.310000  21.635000 ;
      RECT  1.120000  22.325000  1.310000  22.495000 ;
      RECT  1.150000  19.745000  1.310000  19.915000 ;
      RECT  1.150000  20.605000  1.310000  20.775000 ;
      RECT  1.690000  45.545000  4.585000  45.715000 ;
      RECT  2.260000 145.155000  4.700000 145.210000 ;
      RECT  5.875000   5.940000  6.405000   6.465000 ;
      RECT  6.490000  88.950000  9.000000  93.065000 ;
      RECT  7.805000   5.400000 67.100000   6.230000 ;
      RECT  9.300000  32.000000  9.660000  36.750000 ;
      RECT 10.330000  32.000000 10.690000  36.750000 ;
      RECT 11.410000  32.000000 11.665000  37.260000 ;
      RECT 11.940000  31.110000 12.365000  36.765000 ;
      RECT 12.610000  32.000000 13.140000  37.260000 ;
      RECT 13.390000  32.000000 13.920000  36.750000 ;
      RECT 14.170000  32.000000 14.700000  36.750000 ;
      RECT 14.170000  36.750000 14.305000  37.260000 ;
      RECT 14.320000  26.760000 14.500000  29.470000 ;
      RECT 14.320000  29.470000 14.670000  29.570000 ;
      RECT 14.320000  29.570000 14.490000  30.110000 ;
      RECT 14.955000  32.000000 15.485000  37.260000 ;
      RECT 15.105000  26.760000 15.635000  29.690000 ;
      RECT 15.730000  32.000000 16.260000  36.750000 ;
      RECT 15.730000 179.435000 68.925000 179.450000 ;
      RECT 15.730000 179.450000 77.885000 179.980000 ;
      RECT 15.730000 179.980000 68.925000 180.205000 ;
      RECT 15.885000  26.760000 16.415000  29.470000 ;
      RECT 16.510000  32.000000 16.950000  37.260000 ;
      RECT 16.670000  26.760000 17.200000  29.690000 ;
      RECT 17.210000  32.000000 17.650000  36.750000 ;
      RECT 18.035000  26.760000 18.450000  29.470000 ;
      RECT 18.140000  32.060000 18.630000  36.750000 ;
      RECT 19.040000  26.760000 19.455000  29.470000 ;
      RECT 19.050000  32.000000 19.580000  36.750000 ;
      RECT 19.790000  26.760000 20.320000  29.470000 ;
      RECT 20.640000  32.000000 21.170000  36.750000 ;
      RECT 21.690000  26.760000 22.130000  29.470000 ;
      RECT 22.170000  32.000000 22.700000  36.755000 ;
      RECT 23.725000  32.000000 24.255000  36.755000 ;
      RECT 23.800000  26.760000 24.160000  29.470000 ;
      RECT 24.340000  25.580000 26.330000  25.905000 ;
      RECT 24.340000  25.905000 24.835000  29.690000 ;
      RECT 25.015000  26.760000 25.545000  29.470000 ;
      RECT 25.675000  32.250000 26.090000  37.000000 ;
      RECT 25.930000  59.095000 28.100000  60.125000 ;
      RECT 25.935000  57.585000 29.370000  58.865000 ;
      RECT 26.225000  19.595000 26.670000  24.375000 ;
      RECT 26.385000  32.250000 26.865000  37.330000 ;
      RECT 26.390000  26.760000 26.750000  29.690000 ;
      RECT 26.525000  67.105000 29.670000  67.815000 ;
      RECT 26.975000  19.600000 27.420000  24.365000 ;
      RECT 27.045000  32.250000 27.575000  37.000000 ;
      RECT 27.490000  63.970000 29.315000  64.550000 ;
      RECT 27.510000  26.490000 28.090000  30.360000 ;
      RECT 27.675000  68.735000 29.670000  69.445000 ;
      RECT 27.830000  32.245000 28.360000  37.330000 ;
      RECT 28.340000  59.180000 28.510000  59.710000 ;
      RECT 28.605000  32.250000 29.135000  37.005000 ;
      RECT 28.680000  18.995000 29.210000  23.750000 ;
      RECT 28.860000  95.125000 45.710000  95.255000 ;
      RECT 29.035000  56.755000 29.565000  57.285000 ;
      RECT 29.390000  18.965000 30.080000  23.745000 ;
      RECT 29.390000  32.250000 29.920000  37.330000 ;
      RECT 30.165000  32.250000 30.695000  37.000000 ;
      RECT 30.270000  18.995000 30.800000  23.745000 ;
      RECT 30.950000  32.250000 31.375000  37.330000 ;
      RECT 31.660000  32.250000 32.085000  37.005000 ;
      RECT 31.820000  18.995000 32.350000  23.745000 ;
      RECT 32.410000  32.060000 33.070000  36.750000 ;
      RECT 33.500000  31.990000 33.930000  37.080000 ;
      RECT 34.305000  31.975000 34.865000  36.750000 ;
      RECT 35.060000  31.990000 35.490000  37.080000 ;
      RECT 35.865000  31.975000 36.425000  36.750000 ;
      RECT 35.870000  26.885000 36.305000  28.235000 ;
      RECT 36.620000  31.990000 37.050000  37.080000 ;
      RECT 37.425000  31.975000 37.985000  36.750000 ;
      RECT 38.180000  31.990000 38.610000  37.080000 ;
      RECT 38.985000  31.975000 39.545000  36.750000 ;
      RECT 39.270000  26.885000 39.690000  28.235000 ;
      RECT 39.685000  95.955000 45.710000  96.105000 ;
      RECT 39.715000  31.990000 40.090000  36.750000 ;
      RECT 40.580000  32.155000 40.900000  36.710000 ;
      RECT 43.380000  24.850000 43.870000  27.560000 ;
      RECT 43.855000 180.205000 44.500000 180.370000 ;
      RECT 44.200000  33.270000 44.390000  36.510000 ;
      RECT 45.310000  36.340000 46.360000  36.970000 ;
      RECT 49.340000  32.065000 51.760000  32.445000 ;
      RECT 51.105000  32.445000 51.760000  33.690000 ;
      RECT 52.050000  24.855000 52.580000  27.565000 ;
      RECT 53.470000  24.855000 54.000000  27.565000 ;
      RECT 54.870000  24.855000 55.400000  27.565000 ;
      RECT 56.725000 180.205000 57.305000 180.370000 ;
      RECT 59.360000   2.260000 59.720000   3.430000 ;
      RECT 61.115000   5.230000 67.290000   5.345000 ;
      RECT 61.115000   5.345000 67.100000   5.400000 ;
      RECT 61.370000   5.080000 67.290000   5.230000 ;
      RECT 61.560000   4.765000 67.290000   5.080000 ;
      RECT 64.375000   0.250000 66.075000   1.000000 ;
      RECT 65.660000   6.230000 67.100000   9.570000 ;
      RECT 66.390000   9.570000 67.100000   9.575000 ;
      RECT 66.390000   9.575000 69.665000   9.745000 ;
      RECT 66.390000   9.745000 71.650000  10.185000 ;
      RECT 68.290000   1.940000 69.255000   3.960000 ;
      RECT 69.165000 128.445000 79.585000 130.115000 ;
      RECT 69.625000 179.435000 77.885000 179.450000 ;
      RECT 69.625000 179.980000 77.885000 180.205000 ;
      RECT 69.665000  10.185000 71.650000  11.425000 ;
      RECT 72.315000   1.940000 74.335000   4.420000 ;
      RECT 73.080000   8.080000 74.910000   8.830000 ;
      RECT 74.910000   5.170000 76.930000   5.800000 ;
      RECT 74.910000   5.800000 79.430000   7.820000 ;
      RECT 77.195000   3.705000 79.430000   4.420000 ;
      RECT 77.195000   4.420000 77.775000   5.170000 ;
      RECT 77.410000   3.700000 79.430000   3.705000 ;
      RECT 77.410000   7.820000 79.430000   8.080000 ;
      RECT 79.880000  19.485000 80.120000  25.015000 ;
      RECT 79.880000  30.115000 80.120000  35.725000 ;
    LAYER met1 ;
      RECT -0.115000  95.895000  1.495000 130.220000 ;
      RECT -0.115000 131.275000  1.495000 170.090000 ;
      RECT  0.000000   0.000000  5.565000   1.560000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000 62.290000   2.055000 ;
      RECT  0.000000   1.560000  5.565000   1.565000 ;
      RECT  0.000000   1.565000  5.565000   2.055000 ;
      RECT  0.000000   1.565000 35.575000   1.635000 ;
      RECT  0.000000   1.635000 35.505000   1.705000 ;
      RECT  0.000000   1.705000 35.435000   1.775000 ;
      RECT  0.000000   1.775000 35.365000   1.845000 ;
      RECT  0.000000   1.845000 35.295000   1.915000 ;
      RECT  0.000000   1.915000 35.225000   1.985000 ;
      RECT  0.000000   1.985000 35.155000   2.055000 ;
      RECT  0.000000   2.055000  5.565000   2.875000 ;
      RECT  0.000000   2.055000 80.000000 106.585000 ;
      RECT  0.000000   2.875000 11.260000   3.155000 ;
      RECT  0.000000   3.155000 67.995000   4.240000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   4.240000 76.885000   5.515000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   5.515000 80.000000  10.335000 ;
      RECT  0.000000  10.335000  1.340000  11.155000 ;
      RECT  0.000000  11.155000  0.750000  12.425000 ;
      RECT  0.000000  12.425000 80.000000  13.120000 ;
      RECT  0.000000  14.320000 76.495000  23.850000 ;
      RECT  0.000000  14.320000 80.000000  16.455000 ;
      RECT  0.000000  17.275000 78.550000  23.850000 ;
      RECT  0.000000  17.275000 78.550000  29.840000 ;
      RECT  0.000000  17.275000 79.605000  19.205000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  19.205000 79.605000  20.650000 ;
      RECT  0.000000  20.650000 78.550000  29.840000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.850000 79.605000  25.295000 ;
      RECT  0.000000  25.295000 78.845000  36.005000 ;
      RECT  0.000000  25.295000 78.845000  42.035000 ;
      RECT  0.000000  25.295000 80.000000  29.840000 ;
      RECT  0.000000  29.840000 78.845000  42.035000 ;
      RECT  0.000000  29.840000 79.605000  31.400000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.725000 78.845000  34.115000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.440000 79.605000  36.005000 ;
      RECT  0.000000  36.005000 80.000000  42.035000 ;
      RECT  0.000000  42.035000 78.635000  42.340000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.975000 78.635000  43.235000 ;
      RECT  0.000000  43.235000 80.000000  44.355000 ;
      RECT  0.000000  44.355000  1.020000  45.010000 ;
      RECT  0.000000  45.010000  0.965000  45.240000 ;
      RECT  0.000000  45.240000  0.895000  45.310000 ;
      RECT  0.000000  45.310000  0.825000  45.380000 ;
      RECT  0.000000  45.380000  0.755000  45.450000 ;
      RECT  0.000000  45.450000  0.685000  45.520000 ;
      RECT  0.000000  45.520000  0.615000  45.590000 ;
      RECT  0.000000  45.590000  0.545000  45.660000 ;
      RECT  0.000000  45.660000  0.475000  45.730000 ;
      RECT  0.000000  45.730000  0.405000  45.800000 ;
      RECT  0.000000  45.800000  0.335000  45.870000 ;
      RECT  0.000000  45.870000  0.265000  45.940000 ;
      RECT  0.000000  45.940000  0.195000  46.010000 ;
      RECT  0.000000  46.010000  0.125000  46.080000 ;
      RECT  0.000000  46.080000  0.055000  46.150000 ;
      RECT  0.000000  46.445000  0.965000  46.580000 ;
      RECT  0.000000  46.580000  1.050000  47.350000 ;
      RECT  0.000000  47.350000 80.000000  93.020000 ;
      RECT  0.000000  93.020000  1.070000  94.660000 ;
      RECT  0.000000  94.660000 11.550000  94.830000 ;
      RECT  0.000000  94.830000  1.985000  95.615000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 130.500000  4.530000 130.715000 ;
      RECT  0.000000 130.715000  1.980000 130.995000 ;
      RECT  0.000000 170.370000  1.980000 178.680000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 80.000000 179.140000 ;
      RECT  0.000000 179.140000 15.445000 180.290000 ;
      RECT  0.000000 180.290000 15.490000 200.000000 ;
      RECT  0.000000 180.290000 80.000000 198.405000 ;
      RECT  0.000000 198.405000 15.490000 200.000000 ;
      RECT  0.210000  13.400000  0.470000  14.040000 ;
      RECT  0.475000  46.125000  5.000000  46.165000 ;
      RECT  0.545000  46.055000  5.000000  46.125000 ;
      RECT  0.615000  45.985000  5.000000  46.055000 ;
      RECT  0.685000  45.915000  5.000000  45.985000 ;
      RECT  0.750000  11.155000 76.825000  12.425000 ;
      RECT  0.750000  13.120000 80.000000  16.125000 ;
      RECT  0.755000  45.845000  5.000000  45.915000 ;
      RECT  0.825000  45.775000  5.000000  45.845000 ;
      RECT  0.895000  45.705000  5.000000  45.775000 ;
      RECT  0.965000  45.635000  5.000000  45.705000 ;
      RECT  1.035000  45.565000  5.000000  45.635000 ;
      RECT  1.105000  45.495000  5.000000  45.565000 ;
      RECT  1.175000  45.425000  5.000000  45.495000 ;
      RECT  1.245000  45.290000  5.000000  45.355000 ;
      RECT  1.245000  45.355000  5.000000  45.425000 ;
      RECT  1.245000  46.165000  5.000000  46.300000 ;
      RECT  1.300000  44.635000  1.730000  45.290000 ;
      RECT  1.330000  46.300000  2.790000  47.070000 ;
      RECT  1.350000  93.300000  8.265000  94.380000 ;
      RECT  1.620000  10.615000  4.025000  10.875000 ;
      RECT  1.775000  95.615000  1.985000 106.585000 ;
      RECT  1.775000 118.955000  1.985000 130.500000 ;
      RECT  1.775000 130.995000  1.980000 140.430000 ;
      RECT  1.775000 140.430000 80.000000 144.875000 ;
      RECT  1.775000 144.875000  1.980000 170.370000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  2.010000  44.355000 80.000000  45.010000 ;
      RECT  2.260000 130.995000  4.700000 139.510000 ;
      RECT  2.260000 139.510000  4.855000 140.150000 ;
      RECT  2.260000 145.155000  4.700000 178.400000 ;
      RECT  2.265000  95.110000  8.970000  95.900000 ;
      RECT  2.265000  95.900000  4.250000 130.220000 ;
      RECT  3.070000  46.580000 80.000000  47.350000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  4.305000   8.145000 80.000000  11.150000 ;
      RECT  4.305000  11.150000 76.825000  11.155000 ;
      RECT  4.530000  96.180000 80.000000 127.980000 ;
      RECT  4.530000 125.130000 70.100000 128.135000 ;
      RECT  4.530000 128.135000 68.825000 130.425000 ;
      RECT  4.530000 130.425000 70.100000 130.500000 ;
      RECT  4.530000 130.500000 80.000000 130.715000 ;
      RECT  4.980000 130.715000 80.000000 139.230000 ;
      RECT  4.980000 144.875000 80.000000 178.680000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  5.135000 139.230000 80.000000 140.430000 ;
      RECT  5.135000 139.230000 80.000000 144.875000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  47.350000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  45.010000 80.000000  46.580000 ;
      RECT  5.565000   0.000000  6.890000   1.560000 ;
      RECT  5.565000   1.560000 22.990000   1.565000 ;
      RECT  5.845000   2.335000 10.120000   2.595000 ;
      RECT  7.170000   0.270000 10.715000   1.280000 ;
      RECT  8.545000  93.020000 11.550000  94.660000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT 10.400000   2.055000 35.085000   2.125000 ;
      RECT 10.400000   2.125000 35.015000   2.195000 ;
      RECT 10.400000   2.195000 34.945000   2.265000 ;
      RECT 10.400000   2.265000 34.880000   2.330000 ;
      RECT 10.400000   2.330000 13.640000   2.335000 ;
      RECT 10.400000   2.335000 11.260000   2.875000 ;
      RECT 10.995000   0.000000 18.955000   1.560000 ;
      RECT 11.540000   2.615000 35.170000   2.685000 ;
      RECT 11.540000   2.685000 35.100000   2.755000 ;
      RECT 11.540000   2.755000 35.070000   2.785000 ;
      RECT 11.540000   2.785000 18.385000   2.790000 ;
      RECT 11.540000   2.790000 13.990000   2.795000 ;
      RECT 11.540000   2.795000 13.985000   2.800000 ;
      RECT 11.540000   2.800000 12.220000   2.835000 ;
      RECT 11.540000   2.835000 12.185000   2.870000 ;
      RECT 11.540000   2.870000 12.180000   2.875000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 13.760000   2.610000 35.240000   2.615000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 15.725000 179.420000 77.705000 180.010000 ;
      RECT 15.770000 198.685000 56.715000 199.975000 ;
      RECT 18.505000   3.065000 19.370000   3.070000 ;
      RECT 19.235000   0.270000 21.375000   1.280000 ;
      RECT 19.490000   2.785000 28.955000   2.790000 ;
      RECT 21.655000   0.000000 22.990000   1.560000 ;
      RECT 23.270000   0.275000 26.265000   1.285000 ;
      RECT 26.545000   0.000000 33.120000   1.560000 ;
      RECT 26.545000   1.560000 34.265000   1.565000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 30.545000   2.785000 35.065000   2.790000 ;
      RECT 33.400000   0.270000 37.775000   1.280000 ;
      RECT 34.545000   1.280000 37.775000   1.285000 ;
      RECT 35.055000   2.550000 35.245000   2.610000 ;
      RECT 35.125000   2.480000 35.305000   2.550000 ;
      RECT 35.195000   2.410000 35.375000   2.480000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.265000   2.340000 35.445000   2.410000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.335000   2.270000 35.515000   2.340000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.405000   2.200000 35.585000   2.270000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.475000   2.130000 35.655000   2.200000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.515000   2.090000 43.035000   2.130000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.585000   2.020000 42.965000   2.090000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.655000   1.950000 42.895000   2.020000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 38.055000   0.000000 40.785000   1.145000 ;
      RECT 38.055000   1.145000 39.110000   1.670000 ;
      RECT 39.390000   1.425000 43.110000   1.495000 ;
      RECT 39.390000   1.495000 43.180000   1.565000 ;
      RECT 39.390000   1.565000 43.250000   1.635000 ;
      RECT 39.390000   1.635000 43.320000   1.685000 ;
      RECT 41.065000   0.270000 41.935000   1.285000 ;
      RECT 42.215000   0.000000 55.320000   1.145000 ;
      RECT 42.875000   2.130000 43.075000   2.180000 ;
      RECT 42.925000   2.180000 43.125000   2.230000 ;
      RECT 42.930000   2.230000 43.175000   2.235000 ;
      RECT 43.000000   2.235000 51.520000   2.305000 ;
      RECT 43.070000   2.305000 51.520000   2.375000 ;
      RECT 43.110000   1.685000 43.370000   1.755000 ;
      RECT 43.110000   2.375000 51.520000   2.415000 ;
      RECT 43.180000   1.755000 43.440000   1.825000 ;
      RECT 43.200000   1.825000 43.510000   1.845000 ;
      RECT 43.270000   1.145000 62.150000   1.190000 ;
      RECT 43.270000   1.845000 47.840000   1.915000 ;
      RECT 43.315000   1.190000 62.150000   1.235000 ;
      RECT 43.340000   1.915000 47.770000   1.985000 ;
      RECT 43.385000   1.235000 47.725000   1.305000 ;
      RECT 43.410000   1.985000 47.700000   2.055000 ;
      RECT 43.430000   2.055000 47.680000   2.075000 ;
      RECT 43.455000   1.305000 47.655000   1.375000 ;
      RECT 43.525000   1.375000 47.585000   1.445000 ;
      RECT 43.595000   1.445000 47.515000   1.515000 ;
      RECT 43.645000   1.515000 47.465000   1.565000 ;
      RECT 47.630000   1.795000 47.910000   1.845000 ;
      RECT 47.680000   1.745000 47.960000   1.795000 ;
      RECT 47.700000   1.725000 55.040000   1.745000 ;
      RECT 47.770000   1.655000 55.040000   1.725000 ;
      RECT 47.840000   1.585000 55.040000   1.655000 ;
      RECT 47.910000   1.515000 55.040000   1.585000 ;
      RECT 50.840000   2.195000 51.520000   2.235000 ;
      RECT 50.880000   2.155000 51.520000   2.195000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.655000 59.170000   2.695000 ;
      RECT 54.655000   1.745000 55.040000   1.760000 ;
      RECT 54.670000   1.760000 55.040000   1.775000 ;
      RECT 54.675000   1.775000 55.040000   1.780000 ;
      RECT 54.745000   1.780000 54.875000   1.850000 ;
      RECT 54.815000   1.850000 54.875000   1.920000 ;
      RECT 55.155000   2.060000 59.170000   2.655000 ;
      RECT 55.320000   0.000000 59.170000   1.145000 ;
      RECT 55.320000   1.145000 59.170000   1.235000 ;
      RECT 55.320000   1.235000 59.170000   1.920000 ;
      RECT 55.320000   1.920000 59.170000   2.060000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 198.405000 80.000000 198.420000 ;
      RECT 56.995000 198.420000 71.715000 200.000000 ;
      RECT 59.170000   0.000000 62.150000   1.145000 ;
      RECT 59.170000   1.235000 62.150000   1.920000 ;
      RECT 59.450000   2.200000 59.710000   2.850000 ;
      RECT 59.990000   1.920000 62.150000   2.195000 ;
      RECT 59.990000   2.195000 67.995000   3.130000 ;
      RECT 62.830000   0.000000 80.000000   2.055000 ;
      RECT 62.970000   0.000000 64.095000   1.190000 ;
      RECT 62.970000   1.190000 67.995000   1.960000 ;
      RECT 62.970000   1.960000 67.995000   2.195000 ;
      RECT 64.375000   0.260000 67.295000   0.910000 ;
      RECT 67.575000   0.000000 69.205000   1.190000 ;
      RECT 67.995000   1.190000 69.205000   1.960000 ;
      RECT 68.275000   2.240000 68.925000   3.960000 ;
      RECT 69.105000 128.415000 80.145000 130.145000 ;
      RECT 69.205000   0.000000 80.000000   1.190000 ;
      RECT 69.205000   1.190000 80.000000   1.960000 ;
      RECT 69.205000   1.960000 80.000000   3.365000 ;
      RECT 69.205000   3.365000 76.885000   4.240000 ;
      RECT 70.380000 128.260000 80.145000 128.415000 ;
      RECT 70.380000 130.145000 80.145000 130.220000 ;
      RECT 71.995000 198.700000 76.855000 200.000000 ;
      RECT 76.775000  16.735000 77.415000  16.995000 ;
      RECT 77.105000  11.430000 77.365000  12.145000 ;
      RECT 77.135000 198.420000 80.000000 200.000000 ;
      RECT 77.165000   3.645000 77.805000   5.235000 ;
      RECT 77.645000  11.150000 80.000000  12.425000 ;
      RECT 77.695000  16.455000 80.000000  17.275000 ;
      RECT 77.985000 179.140000 80.000000 180.290000 ;
      RECT 78.085000   3.365000 80.000000   5.515000 ;
      RECT 78.705000  42.665000 79.175000  42.695000 ;
      RECT 78.775000  42.595000 79.175000  42.665000 ;
      RECT 78.830000  21.375000 80.115000  23.125000 ;
      RECT 78.845000  42.525000 79.175000  42.595000 ;
      RECT 78.915000  42.315000 79.175000  42.455000 ;
      RECT 78.915000  42.455000 79.175000  42.525000 ;
      RECT 78.915000  42.695000 79.175000  42.955000 ;
      RECT 79.125000  32.005000 80.115000  33.835000 ;
      RECT 79.325000  21.325000 80.115000  21.375000 ;
      RECT 79.345000  23.125000 80.115000  23.195000 ;
      RECT 79.395000  21.255000 80.115000  21.325000 ;
      RECT 79.415000  23.195000 80.115000  23.265000 ;
      RECT 79.455000  42.035000 80.000000  43.235000 ;
      RECT 79.465000  21.185000 80.115000  21.255000 ;
      RECT 79.465000  31.935000 80.115000  32.005000 ;
      RECT 79.465000  33.835000 80.115000  33.905000 ;
      RECT 79.485000  23.265000 80.115000  23.335000 ;
      RECT 79.535000  21.115000 80.115000  21.185000 ;
      RECT 79.535000  31.865000 80.115000  31.935000 ;
      RECT 79.535000  33.905000 80.115000  33.975000 ;
      RECT 79.555000  23.335000 80.115000  23.405000 ;
      RECT 79.605000  17.275000 80.000000  19.205000 ;
      RECT 79.605000  21.045000 80.115000  21.115000 ;
      RECT 79.605000  31.795000 80.115000  31.865000 ;
      RECT 79.605000  33.975000 80.115000  34.045000 ;
      RECT 79.625000  23.405000 80.115000  23.475000 ;
      RECT 79.675000  20.975000 80.115000  21.045000 ;
      RECT 79.675000  31.725000 80.115000  31.795000 ;
      RECT 79.675000  34.045000 80.115000  34.115000 ;
      RECT 79.695000  23.475000 80.115000  23.545000 ;
      RECT 79.745000  20.905000 80.115000  20.975000 ;
      RECT 79.745000  31.655000 80.115000  31.725000 ;
      RECT 79.745000  34.115000 80.115000  34.185000 ;
      RECT 79.765000  23.545000 80.115000  23.615000 ;
      RECT 79.815000  20.835000 80.115000  20.905000 ;
      RECT 79.815000  31.585000 80.115000  31.655000 ;
      RECT 79.815000  34.185000 80.115000  34.255000 ;
      RECT 79.835000  23.615000 80.115000  23.685000 ;
      RECT 79.885000  19.485000 80.115000  20.765000 ;
      RECT 79.885000  20.765000 80.115000  20.835000 ;
      RECT 79.885000  23.685000 80.115000  23.735000 ;
      RECT 79.885000  23.735000 80.115000  25.015000 ;
      RECT 79.885000  30.120000 80.115000  31.515000 ;
      RECT 79.885000  31.515000 80.115000  31.585000 ;
      RECT 79.885000  34.255000 80.115000  34.325000 ;
      RECT 79.885000  34.325000 80.115000  35.725000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  3.095000   4.590000 ;
      RECT  0.000000   0.000000  3.235000   4.535000 ;
      RECT  0.000000   4.535000  3.940000   5.240000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.240000  5.260000   5.435000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.260000   8.410000 ;
      RECT  0.000000   5.490000  5.120000   8.495000 ;
      RECT  0.000000   8.410000  6.435000   9.585000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.435000  38.760000 ;
      RECT  0.000000   9.640000  6.295000  38.705000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.760000  5.835000  39.360000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.305000  5.685000  53.625000 ;
      RECT  0.000000  39.305000  5.695000  42.860000 ;
      RECT  0.000000  39.360000  5.835000  42.915000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.870000  5.685000  43.905000 ;
      RECT  0.000000  42.915000  5.825000  42.925000 ;
      RECT  0.000000  42.925000  5.825000  43.765000 ;
      RECT  0.000000  43.765000  8.055000  44.015000 ;
      RECT  0.000000  43.905000  7.915000  53.625000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.960000  7.915000  53.625000 ;
      RECT  0.000000  44.015000  8.055000  53.680000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.680000  7.835000  53.900000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.845000  7.695000  55.685000 ;
      RECT  0.000000  53.900000  7.835000  55.740000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.740000  7.175000  56.400000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.400000  7.175000  73.785000 ;
      RECT  0.000000  73.785000  7.665000  74.270000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.270000  7.665000  74.850000 ;
      RECT  0.000000  74.330000  7.525000  74.905000 ;
      RECT  0.000000  74.850000  8.070000  75.255000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.975000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.975000  7.595000  75.045000 ;
      RECT  0.000000  75.020000  7.640000  75.310000 ;
      RECT  0.000000  75.045000  7.665000  75.115000 ;
      RECT  0.000000  75.115000  7.735000  75.185000 ;
      RECT  0.000000  75.185000  7.805000  75.255000 ;
      RECT  0.000000  75.255000  7.875000  75.310000 ;
      RECT  0.000000  75.255000  8.070000  77.055000 ;
      RECT  0.000000  75.310000  7.930000  77.005000 ;
      RECT  0.000000  77.005000  7.640000  78.315000 ;
      RECT  0.000000  77.055000  7.980000  77.145000 ;
      RECT  0.000000  77.145000  7.780000  77.685000 ;
      RECT  0.000000  77.685000 76.775000  96.135000 ;
      RECT  0.000000  77.825000 76.635000  96.080000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.135000 76.545000  96.365000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.365000 80.000000 106.585000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.505000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.740000 106.585000 80.000000 118.955000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  3.745000   0.000000  5.280000   4.315000 ;
      RECT  3.745000   4.315000  5.280000   4.535000 ;
      RECT  3.885000   0.000000  5.140000   4.260000 ;
      RECT  3.955000   4.260000  5.140000   4.330000 ;
      RECT  3.960000   4.535000  5.475000   4.730000 ;
      RECT  4.025000   4.330000  5.140000   4.400000 ;
      RECT  4.095000   4.400000  5.140000   4.470000 ;
      RECT  4.165000   4.470000  5.140000   4.540000 ;
      RECT  4.215000   4.540000  5.140000   4.590000 ;
      RECT  5.285000   4.730000  5.965000   5.215000 ;
      RECT  5.770000   5.215000  6.180000   5.435000 ;
      RECT  5.770000   5.435000  6.180000   6.190000 ;
      RECT  5.770000   6.190000  6.085000   6.285000 ;
      RECT  5.770000   6.825000  8.305000   6.920000 ;
      RECT  5.770000   6.920000 13.830000   8.190000 ;
      RECT  5.770000   8.190000 13.830000   9.365000 ;
      RECT  5.790000   0.000000  5.990000   1.610000 ;
      RECT  5.790000   1.610000  8.305000   3.925000 ;
      RECT  5.790000   3.925000  8.305000   4.315000 ;
      RECT  5.790000   4.315000  8.305000   5.215000 ;
      RECT  5.845000   2.335000  6.520000   2.405000 ;
      RECT  5.845000   2.405000  6.590000   2.475000 ;
      RECT  5.845000   2.475000  6.660000   2.545000 ;
      RECT  5.845000   2.545000  6.730000   2.595000 ;
      RECT  5.885000   2.595000  6.780000   2.635000 ;
      RECT  5.910000   6.965000  8.165000   7.060000 ;
      RECT  5.910000   7.060000 13.690000   7.345000 ;
      RECT  5.910000   7.345000 13.690000   8.135000 ;
      RECT  5.925000   2.635000  6.820000   2.675000 ;
      RECT  5.930000   1.815000  6.000000   1.885000 ;
      RECT  5.930000   1.885000  6.070000   1.955000 ;
      RECT  5.930000   1.955000  6.140000   2.025000 ;
      RECT  5.930000   2.025000  6.210000   2.095000 ;
      RECT  5.930000   2.095000  6.280000   2.165000 ;
      RECT  5.930000   2.165000  6.350000   2.235000 ;
      RECT  5.930000   2.235000  6.420000   2.305000 ;
      RECT  5.930000   2.305000  6.490000   2.335000 ;
      RECT  5.930000   2.675000  6.860000   2.680000 ;
      RECT  5.930000   2.680000  6.865000   2.750000 ;
      RECT  5.930000   2.750000  6.935000   2.820000 ;
      RECT  5.930000   2.820000  7.005000   2.890000 ;
      RECT  5.930000   2.890000  7.075000   2.960000 ;
      RECT  5.930000   2.960000  7.145000   3.030000 ;
      RECT  5.930000   3.030000  7.215000   3.100000 ;
      RECT  5.930000   3.100000  7.285000   3.170000 ;
      RECT  5.930000   3.170000  7.355000   3.240000 ;
      RECT  5.930000   3.240000  7.425000   3.310000 ;
      RECT  5.930000   3.310000  7.495000   3.380000 ;
      RECT  5.930000   3.380000  7.565000   3.450000 ;
      RECT  5.930000   3.450000  7.635000   3.520000 ;
      RECT  5.930000   3.520000  7.705000   3.590000 ;
      RECT  5.930000   3.590000  7.775000   3.660000 ;
      RECT  5.930000   3.660000  7.845000   3.730000 ;
      RECT  5.930000   3.730000  7.915000   3.800000 ;
      RECT  5.930000   3.800000  7.985000   3.870000 ;
      RECT  5.930000   3.870000  8.055000   3.940000 ;
      RECT  5.930000   3.940000  8.125000   3.980000 ;
      RECT  5.930000   3.980000  8.165000   4.260000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  6.000000   4.260000  8.165000   4.330000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.070000   4.330000  8.165000   4.400000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.140000   4.400000  8.165000   4.470000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.210000   4.470000  8.165000   4.540000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.280000   4.540000  8.165000   4.610000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.345000  39.580000  9.165000  42.905000 ;
      RECT  6.345000  42.905000  9.145000  42.925000 ;
      RECT  6.350000   4.610000  8.165000   4.680000 ;
      RECT  6.365000  42.925000  8.305000  43.765000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.420000   4.680000  8.165000   4.750000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.490000   4.750000  8.165000   4.820000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.530000   0.000000 12.615000   1.380000 ;
      RECT  6.530000   1.380000 12.615000   3.695000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.560000   4.820000  8.165000   4.890000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.630000   4.890000  8.165000   4.960000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.670000   0.000000 12.475000   1.325000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.690000   5.215000  8.305000   6.825000 ;
      RECT  6.700000   4.960000  8.165000   5.030000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.770000   5.030000  8.165000   5.100000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.830000   5.100000  8.165000   5.160000 ;
      RECT  6.830000   5.160000  8.165000   6.965000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.945000   9.365000 13.830000  18.285000 ;
      RECT  6.945000  18.285000 15.245000  19.700000 ;
      RECT  6.945000  19.700000 15.245000  31.485000 ;
      RECT  6.945000  31.485000 14.830000  31.900000 ;
      RECT  6.945000  31.900000 14.830000  37.240000 ;
      RECT  6.945000  37.240000 13.095000  38.980000 ;
      RECT  6.945000  38.980000 12.495000  39.580000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.310000 13.690000  18.340000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.755000 15.105000  31.430000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.845000 14.690000  37.185000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.715000  56.630000 14.210000  57.835000 ;
      RECT  7.715000  57.835000 14.055000  57.990000 ;
      RECT  7.715000  57.990000 14.055000  58.450000 ;
      RECT  7.715000  58.450000 76.775000  73.555000 ;
      RECT  7.715000  73.555000 76.775000  74.045000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.855000  56.685000 14.070000  57.780000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.935000 13.915000  58.590000 ;
      RECT  7.855000  58.590000 76.635000  73.500000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  74.045000 76.775000  74.620000 ;
      RECT  8.205000  74.620000 76.775000  75.025000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.990000 76.635000  74.565000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.375000  54.130000 14.210000  55.970000 ;
      RECT  8.375000  55.970000 14.210000  56.630000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.515000  54.185000 14.070000  56.025000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.595000  44.245000 11.110000  47.445000 ;
      RECT  8.595000  47.445000 11.880000  48.215000 ;
      RECT  8.595000  48.215000 14.210000  48.745000 ;
      RECT  8.595000  48.745000 14.210000  53.910000 ;
      RECT  8.595000  53.910000 14.210000  54.130000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.610000  75.025000 76.775000  77.135000 ;
      RECT  8.610000  77.135000 76.775000  77.225000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000  77.225000 76.775000  77.685000 ;
      RECT  8.735000  44.300000 10.970000  45.265000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.800000 14.070000  53.965000 ;
      RECT  8.735000  48.800000 14.070000  56.025000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.970000 76.635000  77.080000 ;
      RECT  8.755000  44.280000 10.970000  44.300000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.825000  44.210000 10.970000  44.280000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.845000   3.695000 12.615000   5.410000 ;
      RECT  8.845000   5.410000 13.830000   6.625000 ;
      RECT  8.845000   6.625000 13.830000   6.920000 ;
      RECT  8.895000  44.140000 10.970000  44.210000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.965000  44.070000 10.970000  44.140000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.680000 13.690000   7.060000 ;
      RECT  9.035000  44.000000 10.970000  44.070000 ;
      RECT  9.060000  43.775000 11.110000  44.245000 ;
      RECT  9.105000  43.930000 10.970000  44.000000 ;
      RECT  9.175000  43.860000 10.970000  43.930000 ;
      RECT  9.245000  43.790000 10.970000  43.860000 ;
      RECT  9.315000  43.720000 10.970000  43.790000 ;
      RECT  9.375000  43.660000 10.970000  43.720000 ;
      RECT  9.445000  43.590000 11.030000  43.660000 ;
      RECT  9.515000  43.520000 11.100000  43.590000 ;
      RECT  9.585000  43.450000 11.170000  43.520000 ;
      RECT  9.655000  43.380000 11.240000  43.450000 ;
      RECT  9.725000  43.310000 11.310000  43.380000 ;
      RECT  9.795000  43.240000 11.380000  43.310000 ;
      RECT  9.865000  43.170000 11.450000  43.240000 ;
      RECT  9.935000  43.100000 11.520000  43.170000 ;
      RECT 10.005000  43.030000 11.590000  43.100000 ;
      RECT 10.075000  42.960000 11.660000  43.030000 ;
      RECT 10.145000  42.890000 11.730000  42.960000 ;
      RECT 10.215000  42.820000 11.800000  42.890000 ;
      RECT 10.285000  42.750000 11.870000  42.820000 ;
      RECT 10.355000  42.680000 11.940000  42.750000 ;
      RECT 10.425000  42.610000 12.010000  42.680000 ;
      RECT 10.495000  42.540000 12.080000  42.610000 ;
      RECT 10.565000  42.470000 12.150000  42.540000 ;
      RECT 10.635000  42.400000 12.220000  42.470000 ;
      RECT 10.705000  42.330000 12.290000  42.400000 ;
      RECT 10.775000  42.260000 12.360000  42.330000 ;
      RECT 10.845000  42.190000 12.430000  42.260000 ;
      RECT 10.915000  42.120000 12.500000  42.190000 ;
      RECT 10.985000  42.050000 12.570000  42.120000 ;
      RECT 11.055000  41.980000 12.640000  42.050000 ;
      RECT 11.125000  41.910000 12.710000  41.980000 ;
      RECT 11.195000  41.840000 12.780000  41.910000 ;
      RECT 11.265000  41.770000 12.850000  41.840000 ;
      RECT 11.335000  41.700000 12.920000  41.770000 ;
      RECT 11.405000  41.630000 12.990000  41.700000 ;
      RECT 11.475000  41.560000 13.060000  41.630000 ;
      RECT 11.545000  41.490000 13.130000  41.560000 ;
      RECT 11.615000  41.420000 13.200000  41.490000 ;
      RECT 11.650000  44.005000 29.985000  47.215000 ;
      RECT 11.650000  47.215000 29.985000  47.675000 ;
      RECT 11.685000  41.350000 13.270000  41.420000 ;
      RECT 11.740000  41.295000 13.340000  41.350000 ;
      RECT 11.790000  44.060000 29.845000  47.160000 ;
      RECT 11.810000  41.225000 13.340000  41.295000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.880000  41.155000 13.340000  41.225000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.950000  41.085000 13.340000  41.155000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.020000  41.015000 13.340000  41.085000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.090000  40.945000 13.340000  41.015000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.160000  40.875000 13.340000  40.945000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.230000  40.805000 13.340000  40.875000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.300000  40.735000 13.340000  40.805000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.370000  40.665000 13.340000  40.735000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.440000  40.595000 13.340000  40.665000 ;
      RECT 12.465000  40.370000 13.480000  41.405000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.510000  40.525000 13.340000  40.595000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.580000  40.455000 13.340000  40.525000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.650000  40.385000 13.340000  40.455000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.720000  40.315000 13.340000  40.385000 ;
      RECT 12.745000  40.290000 13.340000  40.315000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.815000  40.220000 13.365000  40.290000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.885000  40.150000 13.435000  40.220000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.955000  40.080000 13.505000  40.150000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 13.025000  40.010000 13.575000  40.080000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.095000  39.940000 13.645000  40.010000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.155000   0.000000 16.170000   2.380000 ;
      RECT 13.155000   2.380000 16.955000   3.160000 ;
      RECT 13.155000   3.160000 16.955000   5.180000 ;
      RECT 13.155000   5.180000 16.955000   6.395000 ;
      RECT 13.165000  39.870000 13.715000  39.940000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.235000  39.800000 13.785000  39.870000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.220000 16.815000   5.125000 ;
      RECT 13.305000  39.730000 13.855000  39.800000 ;
      RECT 13.320000  39.520000 13.480000  40.370000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.375000  39.660000 13.925000  39.730000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.445000  39.590000 13.995000  39.660000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.515000  39.520000 14.065000  39.590000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.585000  39.450000 14.135000  39.520000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.655000  39.380000 14.205000  39.450000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.690000  39.345000 15.195000  39.380000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.760000  39.275000 15.230000  39.345000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.830000  39.205000 15.300000  39.275000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.900000  39.135000 15.370000  39.205000 ;
      RECT 13.910000  47.675000 29.985000  48.515000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.970000  39.065000 15.440000  39.135000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 14.020000  40.600000 29.985000  41.635000 ;
      RECT 14.020000  41.635000 29.985000  44.005000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.040000  38.995000 15.510000  39.065000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.110000  38.925000 15.580000  38.995000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.160000  40.655000 29.845000  41.690000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.180000  38.855000 15.650000  38.925000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.250000  38.785000 15.720000  38.855000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.320000  38.715000 15.790000  38.785000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.370000   6.395000 16.955000   6.615000 ;
      RECT 14.370000   6.615000 16.470000   7.100000 ;
      RECT 14.370000   7.100000 16.470000  11.600000 ;
      RECT 14.370000  11.600000 16.565000  11.695000 ;
      RECT 14.370000  11.695000 16.565000  12.320000 ;
      RECT 14.370000  12.320000 16.470000  12.415000 ;
      RECT 14.370000  12.415000 16.470000  18.055000 ;
      RECT 14.370000  18.055000 16.470000  19.470000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.390000  38.645000 15.860000  38.715000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.460000  38.575000 15.930000  38.645000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.560000 16.745000   6.630000 ;
      RECT 14.510000   6.630000 16.675000   6.700000 ;
      RECT 14.510000   6.700000 16.605000   6.770000 ;
      RECT 14.510000   6.770000 16.535000   6.840000 ;
      RECT 14.510000   6.840000 16.465000   6.910000 ;
      RECT 14.510000   6.910000 16.395000   6.980000 ;
      RECT 14.510000   6.980000 16.330000   7.045000 ;
      RECT 14.510000   7.045000 16.330000  11.655000 ;
      RECT 14.510000  11.655000 16.330000  11.705000 ;
      RECT 14.510000  11.705000 16.380000  11.750000 ;
      RECT 14.510000  11.750000 16.425000  12.265000 ;
      RECT 14.510000  12.265000 16.380000  12.310000 ;
      RECT 14.510000  12.310000 16.335000  12.355000 ;
      RECT 14.510000  12.355000 16.330000  12.360000 ;
      RECT 14.510000  12.360000 16.330000  18.000000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.530000  38.505000 16.000000  38.575000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.560000  40.060000 29.985000  40.600000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000  18.000000 16.330000  18.070000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.600000  38.435000 16.070000  38.505000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000  18.070000 16.330000  18.140000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.670000  38.365000 16.140000  38.435000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000  18.140000 16.330000  18.210000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.740000  38.295000 16.210000  38.365000 ;
      RECT 14.750000  48.515000 29.985000  51.370000 ;
      RECT 14.750000  51.370000 29.565000  51.790000 ;
      RECT 14.750000  51.790000 24.535000  53.195000 ;
      RECT 14.750000  53.195000 24.535000  56.895000 ;
      RECT 14.750000  56.895000 24.210000  57.220000 ;
      RECT 14.750000  57.220000 22.940000  57.765000 ;
      RECT 14.750000  57.765000 22.940000  57.780000 ;
      RECT 14.765000  57.780000 76.775000  57.990000 ;
      RECT 14.790000  18.210000 16.330000  18.280000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.810000  38.225000 16.280000  38.295000 ;
      RECT 14.860000  18.280000 16.330000  18.350000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.880000  38.155000 16.350000  38.225000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.460000 29.845000  51.315000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.650000 24.395000  56.840000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.140000 24.395000  56.840000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.080000 22.800000  57.710000 ;
      RECT 14.930000  18.350000 16.330000  18.420000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.950000  38.085000 16.420000  38.155000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.975000  57.990000 76.775000  58.450000 ;
      RECT 15.000000  18.420000 16.330000  18.490000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.020000  38.015000 16.490000  38.085000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.070000  18.490000 16.330000  18.560000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.090000  37.945000 16.560000  38.015000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.935000 76.635000  58.590000 ;
      RECT 15.140000  18.560000 16.330000  18.630000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.160000  37.875000 16.630000  37.945000 ;
      RECT 15.210000  18.630000 16.330000  18.700000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.230000  37.805000 16.700000  37.875000 ;
      RECT 15.280000  18.700000 16.330000  18.770000 ;
      RECT 15.300000  37.735000 16.770000  37.805000 ;
      RECT 15.350000  18.770000 16.330000  18.840000 ;
      RECT 15.370000  32.130000 16.225000  34.380000 ;
      RECT 15.370000  34.380000 17.435000  35.590000 ;
      RECT 15.370000  35.590000 17.435000  37.335000 ;
      RECT 15.370000  37.335000 17.305000  37.470000 ;
      RECT 15.370000  37.665000 16.840000  37.735000 ;
      RECT 15.420000  18.840000 16.330000  18.910000 ;
      RECT 15.440000  37.595000 16.910000  37.665000 ;
      RECT 15.490000  18.910000 16.330000  18.980000 ;
      RECT 15.510000  32.185000 16.085000  34.435000 ;
      RECT 15.510000  34.435000 16.085000  34.505000 ;
      RECT 15.510000  34.505000 16.155000  34.575000 ;
      RECT 15.510000  34.575000 16.225000  34.645000 ;
      RECT 15.510000  34.645000 16.295000  34.715000 ;
      RECT 15.510000  34.715000 16.365000  34.785000 ;
      RECT 15.510000  34.785000 16.435000  34.855000 ;
      RECT 15.510000  34.855000 16.505000  34.925000 ;
      RECT 15.510000  34.925000 16.575000  34.995000 ;
      RECT 15.510000  34.995000 16.645000  35.065000 ;
      RECT 15.510000  35.065000 16.715000  35.135000 ;
      RECT 15.510000  35.135000 16.785000  35.205000 ;
      RECT 15.510000  35.205000 16.855000  35.275000 ;
      RECT 15.510000  35.275000 16.925000  35.345000 ;
      RECT 15.510000  35.345000 16.995000  35.415000 ;
      RECT 15.510000  35.415000 17.065000  35.485000 ;
      RECT 15.510000  35.485000 17.135000  35.555000 ;
      RECT 15.510000  35.555000 17.205000  35.625000 ;
      RECT 15.510000  35.625000 17.275000  35.645000 ;
      RECT 15.510000  35.645000 17.295000  37.280000 ;
      RECT 15.510000  37.280000 17.225000  37.350000 ;
      RECT 15.510000  37.350000 17.155000  37.420000 ;
      RECT 15.510000  37.420000 17.085000  37.490000 ;
      RECT 15.510000  37.490000 17.050000  37.525000 ;
      RECT 15.510000  37.525000 16.980000  37.595000 ;
      RECT 15.560000  18.980000 16.330000  19.050000 ;
      RECT 15.575000  32.120000 16.085000  32.185000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.630000  19.050000 16.330000  19.120000 ;
      RECT 15.645000  32.050000 16.085000  32.120000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.700000  19.120000 16.330000  19.190000 ;
      RECT 15.715000  31.980000 16.085000  32.050000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.770000  19.190000 16.330000  19.260000 ;
      RECT 15.785000  19.470000 16.470000  31.255000 ;
      RECT 15.785000  31.255000 16.225000  31.500000 ;
      RECT 15.785000  31.500000 16.225000  31.715000 ;
      RECT 15.785000  31.715000 16.225000  32.130000 ;
      RECT 15.785000  31.910000 16.085000  31.980000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.840000  19.260000 16.330000  19.330000 ;
      RECT 15.855000  31.840000 16.085000  31.910000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.910000  19.330000 16.330000  19.400000 ;
      RECT 15.925000  19.400000 16.330000  19.415000 ;
      RECT 15.925000  19.415000 16.330000  31.200000 ;
      RECT 15.925000  31.200000 16.260000  31.270000 ;
      RECT 15.925000  31.270000 16.190000  31.340000 ;
      RECT 15.925000  31.340000 16.120000  31.410000 ;
      RECT 15.925000  31.410000 16.085000  31.445000 ;
      RECT 15.925000  31.445000 16.085000  31.770000 ;
      RECT 15.925000  31.770000 16.085000  31.840000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.445000  39.095000 29.985000  40.060000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.710000   0.000000 22.215000   2.150000 ;
      RECT 16.710000   2.150000 22.215000   2.935000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.765000  31.730000 23.335000  34.150000 ;
      RECT 16.765000  34.150000 23.335000  35.360000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.850000   0.000000 22.075000   2.095000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.905000  31.785000 23.195000  34.095000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.985000  38.555000 22.955000  39.095000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 17.010000   7.330000 22.625000  14.545000 ;
      RECT 17.010000  14.545000 23.515000  15.435000 ;
      RECT 17.010000  15.435000 23.515000  24.940000 ;
      RECT 17.010000  24.940000 23.335000  25.120000 ;
      RECT 17.010000  25.120000 23.335000  31.485000 ;
      RECT 17.010000  31.485000 23.335000  31.730000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.150000   7.385000 22.485000  14.600000 ;
      RECT 17.150000   7.385000 22.485000  15.490000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.490000 23.375000  24.885000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.065000 23.195000  31.540000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.180000  38.355000 23.135000  38.555000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.445000   6.895000 22.625000   7.330000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.495000   2.935000 22.215000   6.480000 ;
      RECT 17.495000   6.480000 22.575000   6.845000 ;
      RECT 17.495000   6.845000 22.625000   6.895000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.880000 22.075000   6.540000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.975000  35.360000 23.335000  37.565000 ;
      RECT 17.975000  37.565000 23.335000  38.355000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.115000  31.540000 23.195000  37.620000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.305000 23.195000  37.620000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 22.755000   0.000000 26.460000   1.835000 ;
      RECT 22.755000   1.835000 28.350000   4.130000 ;
      RECT 22.755000   4.130000 29.070000   4.850000 ;
      RECT 22.755000   4.850000 29.070000   6.255000 ;
      RECT 22.755000   6.255000 29.070000   6.665000 ;
      RECT 22.895000   0.000000 26.320000   1.975000 ;
      RECT 22.895000   0.000000 26.320000   4.185000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   4.185000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.905000 28.930000   6.200000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.165000   6.665000 29.070000   6.920000 ;
      RECT 23.165000   6.920000 31.550000  14.315000 ;
      RECT 23.165000  14.315000 31.550000  15.205000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.610000 28.930000   7.060000 ;
      RECT 23.305000   7.060000 31.410000  14.260000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.875000  25.345000 29.985000  36.515000 ;
      RECT 23.875000  36.515000 30.250000  36.780000 ;
      RECT 23.875000  36.780000 30.250000  37.685000 ;
      RECT 23.875000  37.685000 29.985000  37.950000 ;
      RECT 23.875000  37.950000 29.985000  39.095000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.015000  25.405000 29.845000  37.630000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.835000 30.110000  37.245000 ;
      RECT 24.015000  37.245000 30.110000  37.630000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.895000 29.845000  39.235000 ;
      RECT 24.055000  15.205000 31.550000  16.005000 ;
      RECT 24.055000  16.005000 29.985000  17.570000 ;
      RECT 24.055000  17.570000 29.985000  25.165000 ;
      RECT 24.055000  25.165000 29.985000  25.345000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.150000 31.410000  15.950000 ;
      RECT 24.195000  15.950000 29.845000  25.225000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.515000 29.845000  25.225000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.095000  53.425000 76.775000  57.125000 ;
      RECT 25.095000  57.125000 76.775000  57.780000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.235000  53.480000 76.635000  57.180000 ;
      RECT 25.235000  53.480000 76.635000  57.920000 ;
      RECT 25.235000  53.480000 76.635000  73.500000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.260000  53.260000 76.775000  53.425000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.945000  52.575000 76.775000  53.260000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.165000  52.350000 76.090000  52.575000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 27.000000   0.000000 28.350000   1.835000 ;
      RECT 27.140000   0.000000 28.210000   1.975000 ;
      RECT 28.890000   0.000000 30.610000   2.320000 ;
      RECT 28.890000   2.320000 31.165000   2.880000 ;
      RECT 28.890000   2.880000 31.165000   3.900000 ;
      RECT 28.890000   3.900000 31.165000   4.505000 ;
      RECT 29.030000   0.000000 30.470000   2.380000 ;
      RECT 29.030000   2.380000 30.470000   2.450000 ;
      RECT 29.030000   2.450000 30.540000   2.520000 ;
      RECT 29.030000   2.520000 30.610000   2.590000 ;
      RECT 29.030000   2.590000 30.680000   2.660000 ;
      RECT 29.030000   2.660000 30.750000   2.730000 ;
      RECT 29.030000   2.730000 30.820000   2.800000 ;
      RECT 29.030000   2.800000 30.890000   2.870000 ;
      RECT 29.030000   2.870000 30.960000   2.935000 ;
      RECT 29.030000   2.935000 31.025000   3.845000 ;
      RECT 29.100000   3.845000 31.025000   3.915000 ;
      RECT 29.170000   3.915000 31.025000   3.985000 ;
      RECT 29.240000   3.985000 31.025000   4.055000 ;
      RECT 29.310000   4.055000 31.025000   4.125000 ;
      RECT 29.380000   4.125000 31.025000   4.195000 ;
      RECT 29.450000   4.195000 31.025000   4.265000 ;
      RECT 29.490000   4.505000 31.285000   4.620000 ;
      RECT 29.520000   4.265000 31.025000   4.335000 ;
      RECT 29.590000   4.335000 31.025000   4.405000 ;
      RECT 29.610000   4.620000 31.550000   4.890000 ;
      RECT 29.610000   4.890000 31.550000   6.920000 ;
      RECT 29.660000   4.405000 31.025000   4.475000 ;
      RECT 29.730000   4.475000 31.025000   4.545000 ;
      RECT 29.745000   4.545000 31.025000   4.560000 ;
      RECT 29.750000   4.560000 31.025000   4.565000 ;
      RECT 29.750000   4.565000 31.025000   4.635000 ;
      RECT 29.750000   4.635000 31.100000   4.705000 ;
      RECT 29.750000   4.705000 31.170000   4.775000 ;
      RECT 29.750000   4.775000 31.240000   4.845000 ;
      RECT 29.750000   4.845000 31.310000   4.915000 ;
      RECT 29.750000   4.915000 31.380000   4.945000 ;
      RECT 29.750000   4.945000 31.410000   7.060000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.525000  17.795000 79.180000  36.285000 ;
      RECT 30.525000  36.285000 79.180000  36.550000 ;
      RECT 30.525000  38.180000 79.180000  47.610000 ;
      RECT 30.525000  47.610000 76.090000  50.700000 ;
      RECT 30.525000  50.700000 76.090000  51.620000 ;
      RECT 30.525000  51.620000 76.090000  52.350000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.665000  17.855000 79.175000  36.230000 ;
      RECT 30.665000  38.235000 79.175000  42.955000 ;
      RECT 30.665000  42.955000 75.950000  52.490000 ;
      RECT 30.665000  42.955000 79.040000  47.555000 ;
      RECT 30.665000  47.555000 75.950000  52.490000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.645000 75.950000  51.675000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.790000  36.550000 79.180000  37.915000 ;
      RECT 30.790000  37.915000 79.180000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.930000  17.855000 79.175000  42.955000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.150000   0.000000 31.675000   2.095000 ;
      RECT 31.150000   2.095000 31.675000   2.620000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.235000  17.090000 79.180000  17.795000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.290000   0.000000 31.535000   2.040000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.360000   2.040000 31.535000   2.110000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.430000   2.110000 31.535000   2.180000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.500000   2.180000 31.535000   2.250000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.705000   4.105000 45.105000   4.275000 ;
      RECT 31.705000   4.275000 45.105000   4.660000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.940000   4.245000 44.965000   4.315000 ;
      RECT 31.940000  16.380000 79.180000  17.090000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 32.010000   4.315000 44.965000   4.385000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.080000   4.385000 44.965000   4.455000 ;
      RECT 32.090000   4.660000 45.105000   5.145000 ;
      RECT 32.090000   5.145000 45.715000   5.760000 ;
      RECT 32.090000   5.760000 45.715000   6.920000 ;
      RECT 32.090000   6.920000 78.570000  10.110000 ;
      RECT 32.090000  10.110000 78.475000  10.205000 ;
      RECT 32.090000  10.205000 78.475000  16.235000 ;
      RECT 32.090000  16.235000 78.475000  16.380000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.150000   4.455000 44.965000   4.525000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.215000   0.000000 35.320000   1.840000 ;
      RECT 32.215000   1.840000 34.995000   2.165000 ;
      RECT 32.215000   2.165000 34.995000   4.025000 ;
      RECT 32.215000   4.025000 45.105000   4.105000 ;
      RECT 32.220000   4.525000 44.965000   4.595000 ;
      RECT 32.230000   4.245000 44.965000   4.605000 ;
      RECT 32.230000   4.595000 44.965000   4.605000 ;
      RECT 32.230000   4.605000 44.965000   5.205000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.815000 45.575000   7.060000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.430000   8.230000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.365000 78.565000   9.910000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.045000 78.430000  10.055000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.065000 78.420000  16.290000 ;
      RECT 32.230000  10.065000 78.420000  17.855000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.355000   0.000000 35.180000   1.785000 ;
      RECT 32.355000   1.785000 35.110000   1.855000 ;
      RECT 32.355000   1.855000 35.040000   1.925000 ;
      RECT 32.355000   1.925000 34.970000   1.995000 ;
      RECT 32.355000   1.995000 34.900000   2.065000 ;
      RECT 32.355000   2.065000 34.855000   2.110000 ;
      RECT 32.355000   2.110000 34.855000   4.165000 ;
      RECT 32.355000   4.165000 44.965000   4.245000 ;
      RECT 35.535000   2.390000 38.250000   3.855000 ;
      RECT 35.535000   3.855000 45.105000   4.025000 ;
      RECT 35.675000   2.450000 38.110000   3.995000 ;
      RECT 35.675000   3.995000 44.965000   4.165000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.720000   2.405000 38.110000   2.450000 ;
      RECT 35.790000   2.335000 38.110000   2.405000 ;
      RECT 35.860000   0.000000 38.250000   2.070000 ;
      RECT 35.860000   2.070000 38.250000   2.390000 ;
      RECT 35.860000   2.265000 38.110000   2.335000 ;
      RECT 35.930000   2.195000 38.110000   2.265000 ;
      RECT 36.000000   0.000000 38.110000   2.125000 ;
      RECT 36.000000   2.125000 38.110000   2.195000 ;
      RECT 38.790000   0.000000 45.105000   3.855000 ;
      RECT 38.930000   0.000000 44.965000   3.995000 ;
      RECT 38.930000   0.000000 44.965000   4.605000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 45.645000   0.000000 49.715000   0.220000 ;
      RECT 45.645000   0.220000 49.450000   0.485000 ;
      RECT 45.645000   0.485000 49.450000   0.965000 ;
      RECT 45.645000   0.965000 66.400000   1.135000 ;
      RECT 45.645000   1.135000 66.400000   1.615000 ;
      RECT 45.645000   1.615000 68.135000   4.100000 ;
      RECT 45.645000   4.100000 77.010000   4.920000 ;
      RECT 45.645000   4.920000 77.010000   5.375000 ;
      RECT 45.785000   0.000000 49.310000   0.165000 ;
      RECT 45.785000   0.165000 49.310000   0.430000 ;
      RECT 45.785000   0.165000 49.505000   0.235000 ;
      RECT 45.785000   0.235000 49.435000   0.305000 ;
      RECT 45.785000   0.305000 49.365000   0.375000 ;
      RECT 45.785000   0.375000 49.310000   0.430000 ;
      RECT 45.785000   0.430000 49.310000   1.105000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.240000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   4.240000 76.870000   4.865000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.100000   5.375000 78.570000   5.530000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.255000   5.530000 78.570000   6.920000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.475000 76.870000   5.515000 ;
      RECT 46.395000   5.515000 78.430000   7.060000 ;
      RECT 49.310000   0.000000 49.575000   0.165000 ;
      RECT 50.255000   0.000000 66.695000   0.240000 ;
      RECT 50.255000   0.240000 66.695000   0.485000 ;
      RECT 50.395000   0.000000 50.640000   0.185000 ;
      RECT 50.465000   0.185000 66.555000   0.255000 ;
      RECT 50.500000   0.485000 66.695000   0.840000 ;
      RECT 50.500000   0.840000 66.570000   0.965000 ;
      RECT 50.535000   0.255000 66.555000   0.325000 ;
      RECT 50.605000   0.325000 66.555000   0.395000 ;
      RECT 50.640000   0.000000 66.260000   4.865000 ;
      RECT 50.640000   0.395000 66.555000   0.430000 ;
      RECT 50.640000   0.785000 66.485000   0.855000 ;
      RECT 50.640000   0.855000 66.415000   0.925000 ;
      RECT 50.640000   0.925000 66.345000   0.995000 ;
      RECT 50.640000   0.995000 66.275000   1.065000 ;
      RECT 50.640000   1.065000 66.260000   1.080000 ;
      RECT 66.260000   0.000000 66.555000   0.185000 ;
      RECT 66.260000   0.430000 66.555000   0.785000 ;
      RECT 67.235000   0.000000 68.135000   0.870000 ;
      RECT 67.235000   0.870000 68.135000   1.135000 ;
      RECT 67.375000   0.000000 67.995000   0.815000 ;
      RECT 67.445000   0.815000 67.995000   0.885000 ;
      RECT 67.500000   1.135000 68.135000   1.615000 ;
      RECT 67.515000   0.885000 67.995000   0.955000 ;
      RECT 67.585000   0.955000 67.995000   1.025000 ;
      RECT 67.640000   1.025000 67.995000   1.080000 ;
      RECT 67.640000   1.080000 67.995000   1.755000 ;
      RECT 69.065000   0.000000 76.140000   2.110000 ;
      RECT 69.065000   2.110000 77.010000   2.985000 ;
      RECT 69.065000   2.985000 77.010000   4.100000 ;
      RECT 69.205000   0.000000 76.000000   3.005000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.040000 76.870000   4.240000 ;
      RECT 76.570000  50.910000 79.435000  52.365000 ;
      RECT 76.570000  52.365000 79.435000  53.050000 ;
      RECT 76.710000  50.965000 79.435000  52.310000 ;
      RECT 76.775000  50.900000 79.435000  50.965000 ;
      RECT 76.780000  52.310000 79.435000  52.380000 ;
      RECT 76.845000  50.830000 79.435000  50.900000 ;
      RECT 76.850000  52.380000 79.435000  52.450000 ;
      RECT 76.915000  50.760000 79.435000  50.830000 ;
      RECT 76.920000  52.450000 79.435000  52.520000 ;
      RECT 76.985000  50.690000 79.435000  50.760000 ;
      RECT 76.990000  52.520000 79.435000  52.590000 ;
      RECT 77.055000  50.620000 79.435000  50.690000 ;
      RECT 77.060000   0.000000 77.470000   0.925000 ;
      RECT 77.060000   0.925000 77.350000   1.045000 ;
      RECT 77.060000   1.045000 77.250000   1.565000 ;
      RECT 77.060000   1.565000 77.250000   1.605000 ;
      RECT 77.060000  52.590000 79.435000  52.660000 ;
      RECT 77.100000   1.605000 78.570000   2.535000 ;
      RECT 77.125000  50.550000 79.435000  50.620000 ;
      RECT 77.130000  52.660000 79.435000  52.730000 ;
      RECT 77.195000  50.480000 79.435000  50.550000 ;
      RECT 77.200000  52.730000 79.435000  52.800000 ;
      RECT 77.255000  53.050000 79.435000  96.135000 ;
      RECT 77.255000  96.135000 79.435000  96.280000 ;
      RECT 77.265000  50.410000 79.435000  50.480000 ;
      RECT 77.270000  52.800000 79.435000  52.870000 ;
      RECT 77.335000  50.340000 79.435000  50.410000 ;
      RECT 77.340000  52.870000 79.435000  52.940000 ;
      RECT 77.395000  52.940000 79.435000  52.995000 ;
      RECT 77.395000  52.995000 79.435000  96.080000 ;
      RECT 77.395000  96.280000 80.000000  96.365000 ;
      RECT 77.405000  50.270000 79.435000  50.340000 ;
      RECT 77.465000  96.080000 79.435000  96.150000 ;
      RECT 77.475000  50.200000 79.435000  50.270000 ;
      RECT 77.505000   1.745000 78.430000   1.815000 ;
      RECT 77.535000  96.150000 79.435000  96.220000 ;
      RECT 77.545000  50.130000 79.435000  50.200000 ;
      RECT 77.575000   1.815000 78.430000   1.885000 ;
      RECT 77.595000  96.220000 79.435000  96.280000 ;
      RECT 77.615000  50.060000 79.435000  50.130000 ;
      RECT 77.645000   1.885000 78.430000   1.955000 ;
      RECT 77.665000  96.280000 80.000000  96.350000 ;
      RECT 77.685000  49.990000 79.435000  50.060000 ;
      RECT 77.715000   1.955000 78.430000   2.025000 ;
      RECT 77.735000  96.350000 80.000000  96.420000 ;
      RECT 77.755000  49.920000 79.435000  49.990000 ;
      RECT 77.785000   2.025000 78.430000   2.095000 ;
      RECT 77.805000  96.420000 80.000000  96.490000 ;
      RECT 77.820000  96.490000 80.000000  96.505000 ;
      RECT 77.825000  49.850000 79.435000  49.920000 ;
      RECT 77.855000   2.095000 78.430000   2.165000 ;
      RECT 77.895000  49.780000 79.435000  49.850000 ;
      RECT 77.925000   2.165000 78.430000   2.235000 ;
      RECT 77.965000  49.710000 79.435000  49.780000 ;
      RECT 77.995000   2.235000 78.430000   2.305000 ;
      RECT 78.010000   0.000000 78.565000   0.815000 ;
      RECT 78.010000   0.815000 78.565000   1.045000 ;
      RECT 78.030000   2.535000 78.570000   5.375000 ;
      RECT 78.035000  49.640000 79.435000  49.710000 ;
      RECT 78.065000   2.305000 78.430000   2.375000 ;
      RECT 78.105000  49.570000 79.435000  49.640000 ;
      RECT 78.135000   2.375000 78.430000   2.445000 ;
      RECT 78.150000   0.000000 78.425000   0.760000 ;
      RECT 78.170000   2.445000 78.430000   2.480000 ;
      RECT 78.170000   2.480000 78.430000   5.515000 ;
      RECT 78.175000  49.500000 79.435000  49.570000 ;
      RECT 78.220000   0.760000 78.425000   0.830000 ;
      RECT 78.245000  49.430000 79.435000  49.500000 ;
      RECT 78.290000   0.830000 78.425000   0.900000 ;
      RECT 78.295000   0.900000 78.425000   0.905000 ;
      RECT 78.315000  49.360000 79.435000  49.430000 ;
      RECT 78.350000   1.045000 78.565000   1.275000 ;
      RECT 78.350000   1.275000 78.570000   1.280000 ;
      RECT 78.350000   1.280000 78.570000   1.605000 ;
      RECT 78.385000  49.290000 79.435000  49.360000 ;
      RECT 78.455000  49.220000 79.435000  49.290000 ;
      RECT 78.525000  49.150000 79.435000  49.220000 ;
      RECT 78.595000  49.080000 79.435000  49.150000 ;
      RECT 78.665000  49.010000 79.435000  49.080000 ;
      RECT 78.735000  48.940000 79.435000  49.010000 ;
      RECT 78.805000  48.870000 79.435000  48.940000 ;
      RECT 78.875000  48.800000 79.435000  48.870000 ;
      RECT 78.945000  10.505000 79.435000  16.185000 ;
      RECT 78.945000  16.185000 79.435000  16.675000 ;
      RECT 78.945000  48.730000 79.435000  48.800000 ;
      RECT 79.015000  48.660000 79.435000  48.730000 ;
      RECT 79.045000   0.000000 79.435000   1.065000 ;
      RECT 79.045000   1.065000 79.435000   1.070000 ;
      RECT 79.050000   1.070000 79.435000  10.400000 ;
      RECT 79.050000  10.400000 79.435000  10.505000 ;
      RECT 79.085000  10.560000 79.435000  16.130000 ;
      RECT 79.085000  48.590000 79.435000  48.660000 ;
      RECT 79.135000  10.510000 79.435000  10.560000 ;
      RECT 79.155000  16.130000 79.435000  16.200000 ;
      RECT 79.155000  48.520000 79.435000  48.590000 ;
      RECT 79.185000   0.000000 79.435000   1.010000 ;
      RECT 79.190000   1.010000 79.435000   1.015000 ;
      RECT 79.190000   1.015000 79.435000  10.455000 ;
      RECT 79.190000  10.455000 79.435000  10.510000 ;
      RECT 79.225000  16.200000 79.435000  16.270000 ;
      RECT 79.225000  48.450000 79.435000  48.520000 ;
      RECT 79.295000  16.270000 79.435000  16.340000 ;
      RECT 79.295000  48.380000 79.435000  48.450000 ;
      RECT 79.365000  16.340000 79.435000  16.410000 ;
      RECT 79.365000  48.310000 79.435000  48.380000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.100000 106.585000 ;
      RECT  0.000000 118.955000  0.100000 178.610000 ;
      RECT  0.000000 178.610000  2.960000 181.470000 ;
      RECT  0.000000 178.800000  0.150000 178.950000 ;
      RECT  0.000000 178.950000  0.300000 179.100000 ;
      RECT  0.000000 179.100000  0.450000 179.250000 ;
      RECT  0.000000 179.250000  0.600000 179.400000 ;
      RECT  0.000000 179.400000  0.750000 179.550000 ;
      RECT  0.000000 179.550000  0.900000 179.700000 ;
      RECT  0.000000 179.700000  1.050000 179.850000 ;
      RECT  0.000000 179.850000  1.200000 180.000000 ;
      RECT  0.000000 180.000000  1.350000 180.150000 ;
      RECT  0.000000 180.150000  1.500000 180.300000 ;
      RECT  0.000000 180.300000  1.650000 180.450000 ;
      RECT  0.000000 180.450000  1.800000 180.600000 ;
      RECT  0.000000 180.600000  1.950000 180.750000 ;
      RECT  0.000000 180.750000  2.100000 180.900000 ;
      RECT  0.000000 180.900000  2.250000 181.050000 ;
      RECT  0.000000 181.050000  2.400000 181.200000 ;
      RECT  0.000000 181.200000  2.550000 181.350000 ;
      RECT  0.000000 181.350000  2.700000 181.500000 ;
      RECT  0.000000 181.470000 80.000000 200.000000 ;
      RECT  0.000000 181.500000  2.850000 181.570000 ;
      RECT  0.000000 181.570000  7.970000 184.570000 ;
      RECT  0.000000 184.570000  7.965000 184.575000 ;
      RECT  0.000000 184.575000  3.005000 196.995000 ;
      RECT  0.000000 196.995000 80.000000 200.000000 ;
      RECT  1.320000   0.000000 45.565000  36.930000 ;
      RECT  1.320000  36.930000 46.275000  37.640000 ;
      RECT  1.320000  37.640000 60.310000  47.660000 ;
      RECT  1.320000  47.660000 61.410000  74.310000 ;
      RECT  1.320000  74.310000 62.735000  75.635000 ;
      RECT  1.320000  75.635000 68.390000  76.345000 ;
      RECT  1.320000  76.345000 68.390000 102.210000 ;
      RECT  1.320000 102.210000 78.280000 106.585000 ;
      RECT  1.320000 118.955000 78.280000 176.780000 ;
      RECT  1.320000 176.780000 80.000000 178.110000 ;
      RECT  1.320000 178.110000 80.000000 180.140000 ;
      RECT  1.415000   0.945000 45.465000   1.675000 ;
      RECT  1.420000   0.000000 45.465000   0.945000 ;
      RECT  1.420000   1.675000 45.465000   3.950000 ;
      RECT  1.420000   3.950000  4.425000  36.970000 ;
      RECT  1.420000  36.970000 45.465000  37.120000 ;
      RECT  1.420000  37.120000 45.615000  37.270000 ;
      RECT  1.420000  37.270000 45.765000  37.420000 ;
      RECT  1.420000  37.420000 45.915000  37.570000 ;
      RECT  1.420000  37.570000 46.065000  37.720000 ;
      RECT  1.420000  37.720000 46.215000  37.740000 ;
      RECT  1.420000  37.740000  4.425000  74.350000 ;
      RECT  1.420000  74.350000 61.310000  74.500000 ;
      RECT  1.420000  74.500000 61.460000  74.650000 ;
      RECT  1.420000  74.650000 61.610000  74.800000 ;
      RECT  1.420000  74.800000 61.760000  74.950000 ;
      RECT  1.420000  74.950000 61.910000  75.100000 ;
      RECT  1.420000  75.100000 62.060000  75.250000 ;
      RECT  1.420000  75.250000 62.210000  75.400000 ;
      RECT  1.420000  75.400000 62.360000  75.550000 ;
      RECT  1.420000  75.550000 62.510000  75.700000 ;
      RECT  1.420000  75.700000 62.660000  75.735000 ;
      RECT  1.420000  75.735000 67.640000  75.885000 ;
      RECT  1.420000  75.885000 67.790000  76.035000 ;
      RECT  1.420000  76.035000 67.940000  76.185000 ;
      RECT  1.420000  76.185000 68.090000  76.335000 ;
      RECT  1.420000  76.335000 68.240000  76.385000 ;
      RECT  1.420000  76.385000 68.290000 106.585000 ;
      RECT  1.420000 118.955000  4.460000 121.960000 ;
      RECT  1.420000 121.960000  4.425000 173.875000 ;
      RECT  1.420000 173.875000  4.475000 176.880000 ;
      RECT  1.420000 176.880000  4.475000 176.960000 ;
      RECT  1.420000 176.960000  4.555000 177.040000 ;
      RECT  1.420000 177.040000  7.970000 178.070000 ;
      RECT  1.440000 178.070000 80.000000 178.090000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 178.090000 80.000000 178.110000 ;
      RECT  1.460000 178.110000  7.970000 178.145000 ;
      RECT  1.645000 178.145000 80.000000 178.295000 ;
      RECT  1.795000 178.295000 80.000000 178.445000 ;
      RECT  1.945000 178.445000 80.000000 178.595000 ;
      RECT  2.000000 106.585000 78.280000 118.955000 ;
      RECT  2.095000 178.595000 80.000000 178.745000 ;
      RECT  2.245000 178.745000 80.000000 178.895000 ;
      RECT  2.395000 178.895000 80.000000 179.045000 ;
      RECT  2.545000 179.045000 80.000000 179.195000 ;
      RECT  2.695000 179.195000 80.000000 179.345000 ;
      RECT  2.845000 179.345000 80.000000 179.495000 ;
      RECT  2.995000 179.495000 80.000000 179.645000 ;
      RECT  3.000000 184.570000 77.000000 197.000000 ;
      RECT  3.145000 179.645000 80.000000 179.795000 ;
      RECT  3.295000 179.795000 80.000000 179.945000 ;
      RECT  3.390000 179.945000 80.000000 180.040000 ;
      RECT  4.420000   3.000000 42.465000  38.215000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.740000 57.210000  50.760000 ;
      RECT  4.420000  50.760000 58.310000  75.595000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.735000 65.285000 103.585000 ;
      RECT  4.420000 121.955000 75.175000 176.825000 ;
      RECT  4.460000 103.585000 65.285000 105.310000 ;
      RECT  4.460000 105.310000 75.175000 121.955000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.865000 180.140000 80.000000 181.470000 ;
      RECT  4.965000 178.070000  7.970000 178.110000 ;
      RECT  4.965000 178.145000  7.970000 181.570000 ;
      RECT  7.965000 177.040000 75.175000 179.880000 ;
      RECT  7.965000 179.880000 77.000000 184.570000 ;
      RECT 42.460000   3.950000 45.465000  36.970000 ;
      RECT 42.465000  37.740000 52.000000  40.745000 ;
      RECT 46.495000   0.000000 62.520000   5.430000 ;
      RECT 46.495000   5.430000 61.960000   5.990000 ;
      RECT 46.495000   5.990000 59.300000   7.300000 ;
      RECT 46.495000   7.300000 59.300000  11.060000 ;
      RECT 46.495000  11.060000 61.170000  12.930000 ;
      RECT 46.495000  12.930000 61.170000  18.080000 ;
      RECT 46.495000  18.080000 60.310000  18.940000 ;
      RECT 46.495000  18.940000 60.310000  35.570000 ;
      RECT 46.495000  35.570000 47.660000  36.315000 ;
      RECT 46.495000  36.315000 47.880000  36.535000 ;
      RECT 46.495000  36.535000 47.880000  36.540000 ;
      RECT 46.495000  36.540000 47.880000  36.610000 ;
      RECT 46.565000  36.610000 47.780000  36.710000 ;
      RECT 46.595000   0.000000 62.420000   3.005000 ;
      RECT 46.595000   3.005000 49.600000   5.390000 ;
      RECT 46.595000   5.390000 62.270000   5.540000 ;
      RECT 46.595000   5.540000 62.120000   5.690000 ;
      RECT 46.595000   5.690000 61.970000   5.840000 ;
      RECT 46.595000   5.840000 61.920000   5.890000 ;
      RECT 46.595000   5.890000 60.420000   6.040000 ;
      RECT 46.595000   6.040000 60.270000   6.190000 ;
      RECT 46.595000   6.190000 60.120000   6.340000 ;
      RECT 46.595000   6.340000 59.970000   6.490000 ;
      RECT 46.595000   6.490000 59.820000   6.640000 ;
      RECT 46.595000   6.640000 59.670000   6.790000 ;
      RECT 46.595000   6.790000 59.520000   6.940000 ;
      RECT 46.595000   6.940000 59.370000   7.090000 ;
      RECT 46.595000   7.090000 59.220000   7.240000 ;
      RECT 46.595000   7.240000 59.200000   7.260000 ;
      RECT 46.595000   7.260000 59.200000  35.470000 ;
      RECT 46.595000  11.100000 59.200000  11.250000 ;
      RECT 46.595000  11.250000 59.350000  11.400000 ;
      RECT 46.595000  11.400000 59.500000  11.550000 ;
      RECT 46.595000  11.550000 59.650000  11.700000 ;
      RECT 46.595000  11.700000 59.800000  11.850000 ;
      RECT 46.595000  11.850000 59.950000  12.000000 ;
      RECT 46.595000  12.000000 60.100000  12.150000 ;
      RECT 46.595000  12.150000 60.250000  12.300000 ;
      RECT 46.595000  12.300000 60.400000  12.450000 ;
      RECT 46.595000  12.450000 60.550000  12.600000 ;
      RECT 46.595000  12.600000 60.700000  12.750000 ;
      RECT 46.595000  12.750000 60.850000  12.900000 ;
      RECT 46.595000  12.900000 61.000000  12.970000 ;
      RECT 46.595000  18.040000 60.920000  18.190000 ;
      RECT 46.595000  18.190000 60.770000  18.340000 ;
      RECT 46.595000  18.340000 60.620000  18.490000 ;
      RECT 46.595000  18.490000 60.470000  18.640000 ;
      RECT 46.595000  18.640000 60.320000  18.790000 ;
      RECT 46.595000  18.790000 60.210000  18.900000 ;
      RECT 46.595000  35.470000 47.560000  36.355000 ;
      RECT 46.595000  36.355000 47.560000  36.425000 ;
      RECT 46.595000  36.425000 47.630000  36.495000 ;
      RECT 46.595000  36.495000 47.700000  36.500000 ;
      RECT 46.650000  36.500000 47.705000  36.555000 ;
      RECT 46.705000  36.555000 47.760000  36.610000 ;
      RECT 48.310000  37.640000 60.210000  37.740000 ;
      RECT 48.460000  37.490000 60.210000  37.640000 ;
      RECT 48.610000  37.340000 60.210000  37.490000 ;
      RECT 48.760000  37.190000 60.210000  37.340000 ;
      RECT 48.810000  36.545000 60.310000  37.000000 ;
      RECT 48.810000  37.000000 60.310000  37.640000 ;
      RECT 48.910000  36.585000 52.145000  37.040000 ;
      RECT 48.910000  37.040000 60.210000  37.190000 ;
      RECT 49.025000  36.470000 60.210000  36.585000 ;
      RECT 49.040000  35.570000 60.310000  36.315000 ;
      RECT 49.040000  36.315000 60.310000  36.545000 ;
      RECT 49.140000  35.470000 52.145000  36.585000 ;
      RECT 49.140000  36.355000 60.210000  36.470000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.015000 56.200000  12.345000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.215000 58.070000  16.795000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.655000 57.210000  32.470000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.910000  37.830000 57.210000  38.285000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.140000  32.470000 57.210000  37.600000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 56.825000   3.005000 62.420000   5.390000 ;
      RECT 57.205000  18.900000 60.210000  37.040000 ;
      RECT 57.205000  37.740000 60.210000  47.760000 ;
      RECT 57.210000  47.760000 61.310000  50.765000 ;
      RECT 58.065000  12.970000 61.070000  18.040000 ;
      RECT 58.305000  50.765000 61.310000  74.350000 ;
      RECT 60.685000   7.875000 62.520000   7.930000 ;
      RECT 60.685000   7.930000 62.520000  10.485000 ;
      RECT 60.685000  10.485000 62.520000  12.320000 ;
      RECT 60.785000   7.915000 62.365000   7.945000 ;
      RECT 60.785000   7.945000 62.395000   7.970000 ;
      RECT 60.785000   7.970000 62.420000  10.445000 ;
      RECT 60.930000   7.770000 62.220000   7.915000 ;
      RECT 60.935000  10.445000 62.420000  10.595000 ;
      RECT 61.080000   7.620000 62.070000   7.770000 ;
      RECT 61.085000  10.595000 62.420000  10.745000 ;
      RECT 61.190000   7.370000 62.465000   7.875000 ;
      RECT 61.230000   7.470000 61.920000   7.620000 ;
      RECT 61.235000  10.745000 62.420000  10.895000 ;
      RECT 61.385000  10.895000 62.420000  11.045000 ;
      RECT 61.535000  11.045000 62.420000  11.195000 ;
      RECT 61.685000  11.195000 62.420000  11.345000 ;
      RECT 61.695000  19.515000 62.325000  34.720000 ;
      RECT 61.795000  19.555000 62.225000  34.680000 ;
      RECT 61.795000  34.680000 62.075000  34.830000 ;
      RECT 61.795000  34.830000 61.925000  34.980000 ;
      RECT 61.835000  11.345000 62.420000  11.495000 ;
      RECT 61.925000  19.425000 62.225000  19.555000 ;
      RECT 61.985000  11.495000 62.420000  11.645000 ;
      RECT 62.075000  19.275000 62.225000  19.425000 ;
      RECT 62.135000  11.645000 62.420000  11.795000 ;
      RECT 62.285000  11.795000 62.420000  11.945000 ;
      RECT 63.080000  36.325000 78.280000  72.880000 ;
      RECT 63.080000  72.880000 78.280000  73.965000 ;
      RECT 63.180000  36.365000 67.095000  39.370000 ;
      RECT 63.180000  39.370000 66.185000  69.835000 ;
      RECT 63.180000  69.835000 71.940000  72.840000 ;
      RECT 63.195000  36.350000 78.180000  36.365000 ;
      RECT 63.330000  72.840000 78.180000  72.990000 ;
      RECT 63.345000  36.200000 78.180000  36.350000 ;
      RECT 63.480000  72.990000 78.180000  73.140000 ;
      RECT 63.495000  36.050000 78.180000  36.200000 ;
      RECT 63.630000  73.140000 78.180000  73.290000 ;
      RECT 63.645000  35.900000 78.180000  36.050000 ;
      RECT 63.780000  73.290000 78.180000  73.440000 ;
      RECT 63.795000  35.750000 78.180000  35.900000 ;
      RECT 63.930000  73.440000 78.180000  73.590000 ;
      RECT 63.945000  35.600000 78.180000  35.750000 ;
      RECT 63.995000  18.390000 78.280000  35.410000 ;
      RECT 63.995000  35.410000 78.280000  36.325000 ;
      RECT 64.080000  73.590000 78.180000  73.740000 ;
      RECT 64.095000  18.430000 67.290000  21.435000 ;
      RECT 64.095000  21.435000 67.100000  35.450000 ;
      RECT 64.095000  35.450000 78.180000  35.600000 ;
      RECT 64.190000   0.000000 78.280000  18.195000 ;
      RECT 64.190000  18.195000 78.280000  18.390000 ;
      RECT 64.190000  18.335000 78.180000  18.430000 ;
      RECT 64.205000  73.740000 78.180000  73.865000 ;
      RECT 64.290000   0.000000 78.180000   7.455000 ;
      RECT 64.290000   2.690000 78.180000   2.735000 ;
      RECT 64.290000   2.735000 78.225000   2.780000 ;
      RECT 64.290000   2.780000 78.270000   2.785000 ;
      RECT 64.290000   2.785000 78.180000  18.235000 ;
      RECT 64.290000  18.235000 78.180000  18.335000 ;
      RECT 66.180000  37.610000 75.175000  70.865000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 67.095000  19.675000 75.175000  36.695000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.290000   3.000000 75.175000   3.935000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.030000 75.270000   4.455000 ;
      RECT 67.290000   4.455000 75.175000  19.480000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 68.680000  73.965000 78.280000  75.345000 ;
      RECT 68.870000  73.865000 78.180000  74.015000 ;
      RECT 69.020000  74.015000 78.180000  74.165000 ;
      RECT 69.170000  74.165000 78.180000  74.315000 ;
      RECT 69.320000  74.315000 78.180000  74.465000 ;
      RECT 69.470000  74.465000 78.180000  74.615000 ;
      RECT 69.620000  74.615000 78.180000  74.765000 ;
      RECT 69.770000  74.765000 78.180000  74.915000 ;
      RECT 69.920000  74.915000 78.180000  75.065000 ;
      RECT 70.060000  75.345000 78.280000 102.210000 ;
      RECT 70.070000  75.065000 78.180000  75.215000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.160000  73.865000 78.180000 118.955000 ;
      RECT 70.160000  75.215000 78.180000  75.305000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.060000 75.175000 105.310000 ;
      RECT 75.175000  18.430000 78.180000  35.450000 ;
      RECT 75.175000  36.365000 78.180000  72.840000 ;
      RECT 75.175000 118.955000 78.180000 176.880000 ;
      RECT 75.175000 176.880000 80.000000 179.885000 ;
      RECT 75.270000   2.785000 78.275000   7.455000 ;
      RECT 76.995000 179.885000 80.000000 196.995000 ;
      RECT 78.180000   1.160000 78.190000   1.490000 ;
      RECT 79.870000   0.000000 80.000000 176.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000 80.000000   1.635000 ;
      RECT  0.000000   7.885000  4.675000   8.485000 ;
      RECT  0.000000   7.885000 80.000000   8.485000 ;
      RECT  0.000000  13.935000  4.675000  14.535000 ;
      RECT  0.000000  13.935000 80.000000  14.535000 ;
      RECT  0.000000  18.785000  4.675000  19.385000 ;
      RECT  0.000000  18.785000 80.000000  19.385000 ;
      RECT  0.000000  24.835000  4.675000  25.435000 ;
      RECT  0.000000  24.835000 80.000000  25.435000 ;
      RECT  0.000000  30.885000  4.675000  31.485000 ;
      RECT  0.000000  30.885000 80.000000  31.485000 ;
      RECT  0.000000  35.735000  4.675000  36.335000 ;
      RECT  0.000000  35.735000 80.000000  36.335000 ;
      RECT  0.000000  40.585000  4.675000  41.185000 ;
      RECT  0.000000  40.585000 80.000000  41.185000 ;
      RECT  0.000000  46.635000  4.675000  47.335000 ;
      RECT  0.000000  46.635000 80.000000  47.435000 ;
      RECT  0.000000  57.035000 80.000000  57.835000 ;
      RECT  0.000000  57.135000  4.675000  57.835000 ;
      RECT  0.000000  63.085000  4.675000  63.685000 ;
      RECT  0.000000  63.085000 80.000000  63.685000 ;
      RECT  0.000000  68.935000  4.675000  69.635000 ;
      RECT  0.000000  68.935000 80.000000  69.635000 ;
      RECT  0.000000  95.400000  3.005000 104.215000 ;
      RECT  0.000000  95.400000 80.000000 104.315000 ;
      RECT  0.000000 104.215000  9.485000 104.365000 ;
      RECT  0.000000 104.315000  7.705000 106.285000 ;
      RECT  0.000000 104.365000  9.335000 104.515000 ;
      RECT  0.000000 104.515000  9.185000 104.665000 ;
      RECT  0.000000 104.665000  9.035000 104.815000 ;
      RECT  0.000000 104.815000  8.885000 104.965000 ;
      RECT  0.000000 104.965000  8.735000 105.115000 ;
      RECT  0.000000 105.115000  8.585000 105.265000 ;
      RECT  0.000000 105.265000  8.435000 105.415000 ;
      RECT  0.000000 105.415000  8.285000 105.565000 ;
      RECT  0.000000 105.565000  8.135000 105.715000 ;
      RECT  0.000000 105.715000  7.985000 105.865000 ;
      RECT  0.000000 105.865000  7.835000 106.015000 ;
      RECT  0.000000 106.015000  7.685000 106.165000 ;
      RECT  0.000000 106.165000  7.665000 106.185000 ;
      RECT  0.000000 106.185000  1.600000 106.585000 ;
      RECT  0.000000 106.285000  1.700000 106.585000 ;
      RECT  0.000000 118.955000  1.600000 119.355000 ;
      RECT  0.000000 118.955000  1.700000 119.255000 ;
      RECT  0.000000 119.255000  9.685000 121.550000 ;
      RECT  0.000000 119.355000  7.350000 119.505000 ;
      RECT  0.000000 119.505000  7.500000 119.655000 ;
      RECT  0.000000 119.655000  7.650000 119.805000 ;
      RECT  0.000000 119.805000  7.800000 119.955000 ;
      RECT  0.000000 119.955000  7.950000 120.105000 ;
      RECT  0.000000 120.105000  8.100000 120.255000 ;
      RECT  0.000000 120.255000  8.250000 120.405000 ;
      RECT  0.000000 120.405000  8.400000 120.555000 ;
      RECT  0.000000 120.555000  8.550000 120.705000 ;
      RECT  0.000000 120.705000  8.700000 120.855000 ;
      RECT  0.000000 120.855000  8.850000 121.005000 ;
      RECT  0.000000 121.005000  9.000000 121.155000 ;
      RECT  0.000000 121.155000  9.150000 121.305000 ;
      RECT  0.000000 121.305000  9.300000 121.455000 ;
      RECT  0.000000 121.455000  9.450000 121.605000 ;
      RECT  0.000000 121.550000 80.000000 175.385000 ;
      RECT  0.000000 121.605000  9.600000 121.650000 ;
      RECT  0.000000 121.650000 15.900000 124.655000 ;
      RECT  0.000000 124.655000  3.005000 172.380000 ;
      RECT  0.000000 172.380000  4.670000 175.385000 ;
      RECT  1.365000  14.535000  4.675000  18.785000 ;
      RECT  1.365000  14.535000 78.635000  18.785000 ;
      RECT  1.455000  70.310000  4.675000  94.885000 ;
      RECT  1.570000  47.435000 78.430000  57.035000 ;
      RECT  1.670000   1.635000 78.330000   4.640000 ;
      RECT  1.670000   1.635000 78.330000   7.885000 ;
      RECT  1.670000   4.640000  4.675000   7.885000 ;
      RECT  1.670000   8.485000  4.675000  13.935000 ;
      RECT  1.670000   8.485000 78.330000  13.935000 ;
      RECT  1.670000  19.385000  4.675000  24.835000 ;
      RECT  1.670000  19.385000 78.330000  24.835000 ;
      RECT  1.670000  25.435000  4.675000  30.885000 ;
      RECT  1.670000  25.435000 78.330000  30.885000 ;
      RECT  1.670000  31.485000  4.675000  35.735000 ;
      RECT  1.670000  31.485000 78.330000  35.735000 ;
      RECT  1.670000  36.335000  4.675000  40.585000 ;
      RECT  1.670000  36.335000 78.330000  40.585000 ;
      RECT  1.670000  41.185000  4.675000  46.635000 ;
      RECT  1.670000  41.185000 78.330000  46.635000 ;
      RECT  1.670000  47.335000  4.675000  57.135000 ;
      RECT  1.670000  57.835000  4.675000  63.085000 ;
      RECT  1.670000  57.835000 78.330000  63.085000 ;
      RECT  1.670000  63.685000  4.675000  68.935000 ;
      RECT  1.670000  63.685000 78.330000  68.935000 ;
      RECT  1.670000  69.635000  4.675000  70.310000 ;
      RECT  1.670000  69.635000 78.330000  95.400000 ;
      RECT  1.670000  94.885000 78.330000 104.215000 ;
      RECT  1.670000 175.385000  4.675000 196.995000 ;
      RECT  1.670000 175.385000 78.330000 200.000000 ;
      RECT  1.670000 196.995000 78.330000 200.000000 ;
      RECT  3.000000  98.400000 77.000000 101.210000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.650000 77.000000 172.385000 ;
      RECT  4.455000  73.310000 75.330000  91.880000 ;
      RECT  4.670000   3.000000 75.330000  73.310000 ;
      RECT  4.670000  91.880000 75.330000  98.400000 ;
      RECT  4.670000 172.385000 75.330000 197.000000 ;
      RECT  9.880000 121.400000 12.460000 121.650000 ;
      RECT 12.800000 104.315000 80.000000 121.550000 ;
      RECT 12.900000  95.400000 80.000000 121.650000 ;
      RECT 15.900000 101.210000 77.000000 124.650000 ;
      RECT 75.325000   4.640000 78.330000   7.885000 ;
      RECT 75.325000   7.885000 80.000000   8.485000 ;
      RECT 75.325000   8.485000 78.330000  13.935000 ;
      RECT 75.325000  13.935000 80.000000  14.535000 ;
      RECT 75.325000  14.535000 78.635000  18.785000 ;
      RECT 75.325000  18.785000 80.000000  19.385000 ;
      RECT 75.325000  19.385000 78.330000  24.835000 ;
      RECT 75.325000  24.835000 80.000000  25.435000 ;
      RECT 75.325000  25.435000 78.330000  30.885000 ;
      RECT 75.325000  30.885000 80.000000  31.485000 ;
      RECT 75.325000  31.485000 78.330000  35.735000 ;
      RECT 75.325000  35.735000 80.000000  36.335000 ;
      RECT 75.325000  36.335000 78.330000  40.585000 ;
      RECT 75.325000  40.585000 80.000000  41.185000 ;
      RECT 75.325000  41.185000 78.330000  46.635000 ;
      RECT 75.325000  46.635000 80.000000  47.335000 ;
      RECT 75.325000  47.335000 78.330000  57.135000 ;
      RECT 75.325000  57.135000 80.000000  57.835000 ;
      RECT 75.325000  57.835000 78.330000  63.085000 ;
      RECT 75.325000  63.085000 80.000000  63.685000 ;
      RECT 75.325000  63.685000 78.330000  68.935000 ;
      RECT 75.325000  68.935000 80.000000  69.635000 ;
      RECT 75.325000  69.635000 78.330000  94.885000 ;
      RECT 75.325000 175.385000 78.330000 196.995000 ;
      RECT 75.330000 172.380000 80.000000 175.385000 ;
      RECT 76.995000 121.650000 80.000000 172.380000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 124.670000 ;
      RECT  0.000000 124.670000 31.315000 147.815000 ;
      RECT  0.000000 147.815000 80.000000 200.000000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT 54.455000 124.670000 80.000000 147.815000 ;
  END
END sky130_fd_io__top_gpiov2
END LIBRARY