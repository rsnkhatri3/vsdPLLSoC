`default_nettype none
`timescale 1 ns / 1 ps

module simple_por(
    inout vdd3v3,
    inout vdd1v8,
    inout vss,
    output porb_h,
    output porb_l,
    output por_l
);










endmodule
`default_nettype wire
