magic
tech sky130A
magscale 1 2
timestamp 1606744421
<< metal2 >>
rect 99 0 4879 148
rect 5179 0 5579 107
rect 10078 0 14858 148
<< metal3 >>
rect 99 0 4879 391
rect 5179 0 7379 545
rect 7578 0 9778 2266
rect 10078 0 14858 18037
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 7329 27865 7594 29187
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__hvc_clampv2  sky130_fd_io__hvc_clampv2_0
timestamp 1606744421
transform 1 0 0 0 1 0
box 0 0 15000 40000
<< labels >>
flabel metal2 5179 0 5579 107 2 FreeSans 1000 90 0 0 OGC_HVC
port 4 nsew default bidirectional
flabel metal5 7329 27865 7594 29187 0 FreeSans 2000 0 0 0 P_PAD
port 17 nsew default bidirectional
rlabel metal4 s 14746 10625 15000 11221 1 AMUXBUS_A
port 8 nsew default bidirectional
rlabel metal4 s 14746 9673 15000 10269 1 AMUXBUS_B
port 7 nsew default bidirectional
rlabel metal3 s 7578 0 9778 2266 1 DRN_HVC
port 2 nsew default bidirectional
rlabel metal3 s 10078 0 14858 18037 1 P_CORE
port 1 nsew default bidirectional
rlabel metal3 s 5179 0 7379 545 1 SRC_BDY_HVC
port 3 nsew default bidirectional
rlabel metal5 s 14746 1797 15000 2687 1 VCCD
port 14 nsew default bidirectional
rlabel metal5 s 14746 427 15000 1477 1 VCCHIB
port 15 nsew default bidirectional
rlabel metal5 s 14807 3007 15000 3657 1 VDDA
port 13 nsew default bidirectional
rlabel metal5 s 14746 14007 15000 18997 1 VDDIO
port 10 nsew default bidirectional
rlabel metal5 s 14746 12837 15000 13687 1 VDDIO_Q
port 9 nsew default bidirectional
rlabel metal5 s 14746 9547 15000 11347 1 VSSA
port 5 nsew default bidirectional
rlabel metal5 s 14746 8337 15000 9227 1 VSSD
port 6 nsew default bidirectional
rlabel metal5 s 14746 5187 15000 6077 1 VSSIO
port 12 nsew default bidirectional
rlabel metal5 s 14746 11667 15000 12517 1 VSSIO_Q
port 16 nsew default bidirectional
rlabel metal5 s 14746 6397 15000 7047 1 VSWITCH
port 11 nsew default bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 15000 40000
string GDS_FILE /home/roshan/Desktop/pdks/sky130A/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 9954396
string GDS_START 9944920
<< end >>
