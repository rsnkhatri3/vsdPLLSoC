`include "sky130_fd_io__top_ground_hvc_wpad.v"
`include "sky130_fd_io__top_ground_lvc_wpad.v"
//`include "sky130_fd_io__top_power_hvc_wpadv2.v"
`include "sky130_fd_io__top_power_lvc_wpad.v"
`include "sky130_fd_io__top_gpiov2.v"
`include "sky130_ef_io__vddio_hvc_pad.v"
`include "sky130_ef_io__vdda_hvc_pad.v"
`include "sky130_ef_io__corner_pad.v"


module chip_io (input GPIO_0,
                input GPIO_1,
	        input GPIO_2,
	        input GPIO_3, 
		output B_0_pll,
	        output B_1_pll, 
		output B_2_pll, 
		output B_3_pll, 
		input REF_CLK, 
		output REF_CLK_pll, 
		output CLK, 
		input CLK_pll, 
		input VCO_IN, 
		output VCO_IN_pll, 
		input EN_CP, 
		output EN_CP_pll, 
		input EN_VCO, 
		output EN_VCO_pll, 
		output B_CP, 
		input B_CP_pll, 
		output B_VCO, 
		input B_VCO_pll, 
		input VDDA2, 
		input VSSA, 
		input VDDD2,
		input VSSD,
		input VDDR,
		input GNDR,
		input VDDO,
		input GNDO,
		input PORB);






wire GPIO_0;
wire GPIO_1;
wire GPIO_2;
wire GPIO_3;
wire TIE_HI_ESD;
wire TIE_LO_ESD;
wire B_1_pll;
wire B_2_pll;
wire B_3_pll;
wire B_0_pll;

wire REF_CLK;
wire REF_CLK_pll;

wire CLK;
wire CLK_pll;

wire VCO_IN;
wire VCO_IN_pll;

wire EN_CP;
wire EN_CP_pll;

wire EN_VCO;
wire EN_VCO_pll;

wire B_CP;
wire B_CP_pll;

wire B_VCO;
wire B_VCO_pll;


wire   VDDA;
wire   VSSA;
wire   VSSD;
wire   VDDD;

wire   VDDR;
wire   GNDR;
wire   VDDO;
wire   GNDO;

wire   VDDIO;
wire   VSSIO;

wire   VDDA1;
wire   VSSA1;

wire   VCCD1;
wire   VSSD1;

//assign VDDIO = VDDR_pll;
assign VSSIO = GNDR_pll;

assign VDDA1 = VDDO_pll;
assign VSSA1 = GNDO_pll;

assign VCCD1 = VDDD_pll;
assign VSSD1 = VSSD_pll;



wire   VDDA_pll;
wire   VSSA_pll;
wire   VSSD_pll;
wire   VDDD_pll;

wire   VDDR_pll;
wire   GNDR_pll;
wire   VDDO_pll;
wire   GNDO_pll;

wire   PORB;






























sky130_fd_io__top_gpiov2 GPIO_0_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(GPIO_0), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(B_0_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );



sky130_fd_io__top_gpiov2 GPIO_1_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(GPIO_1), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(B_1_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );


sky130_fd_io__top_gpiov2 GPIO_2_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(GPIO_2), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(B_2_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),  
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );



sky130_fd_io__top_gpiov2 GPIO_3_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                         
                                  .PAD(GPIO_3), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(B_3_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );


sky130_fd_io__top_gpiov2 ENb_VCO_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(EN_VCO), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(EN_VCO_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                 
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );



sky130_fd_io__top_gpiov2 ENb_CP_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(EN_CP), 
                                  
                                  .DM({VSSD1,VSSD1,VCCD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(EN_CP_pll), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VCCD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(VSSD1), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );


sky130_fd_io__top_gpiov2 B_VCO_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(B_VCO), 
                                  
                                  .DM({VCCD1,VCCD1,VSSD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VSSD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(B_VCO_pll), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );


sky130_fd_io__top_gpiov2 B_CP_PAD (.IN_H(),
                                  .PAD_A_NOESD_H(),
                                  .PAD_A_ESD_0_H(),
                                  .PAD_A_ESD_1_H(),
                                  
                                  .PAD(B_CP), 
                                  
                                  .DM({VCCD1,VCCD1,VSSD1}), 
                                  .HLD_H_N(VDDIO), 
                                 
                                  .IN(), 
                                  
                                  .INP_DIS(VSSD1), 
                                  .IB_MODE_SEL(VSSD1), 
                                  .ENABLE_H(PORB),      //DOUBT
                                  .ENABLE_VDDA_H(VSSA1),   
                                  .ENABLE_INP_H(TIE_LO_ESD),   
                                  .OE_N(VSSD1),
                                  .TIE_HI_ESD(TIE_HI_ESD), 
                                  .TIE_LO_ESD(TIE_LO_ESD), 
                                  .SLOW(VSSD1), 
                                  .VTRIP_SEL(VSSD1), 
                                  .HLD_OVR(VSSD1), 
                                  .ANALOG_EN(VSSD1), 
                                  .ANALOG_SEL(VSSD1), 
                                  .ENABLE_VDDIO(VCCD1),         
                                  .ENABLE_VSWITCH_H(VSSA1),     
                                  .ANALOG_POL(VSSD1), 
                                  .OUT(B_CP_pll), 
                                  .AMUXBUS_A(), 
                                  .AMUXBUS_B()
                                  
                                 // .VSSA(VSSA1), 
                                 // .VDDA(VDDA1), 
                                 // .VSWITCH(VDDIO), 
                                 // .VDDIO_Q(), 
                                 // .VCCHIB(VCCD1), 
                                 // .VDDIO(VDDIO), 
                                 // .VCCD(VCCD1), 
                                 // .VSSIO(VSSIO),
                                 // .VSSD(VSSD1), 
                                 // .VSSIO_Q()
                                );                                


sky130_fd_io__top_power_lvc_wpad VCO_IN_PAD ( .P_PAD(VCO_IN), 
                                   .AMUXBUS_A(), 
                                   .AMUXBUS_B()
                                  // .P_CORE(VCO_IN_pll), 
                                  // .BDY2_B2B(VSSA1), 
                                  // .DRN_LVC1(VDDA1), 
                                  // .DRN_LVC2(), 
                                  // .OGC_LVC(), 
                                  // .SRC_BDY_LVC1(VSSA1), 
                                  // .SRC_BDY_LVC2(), 
                                   
                                  // .VSSA(VSSA1), 
                                  // .VDDA(VDDA1), 
                                  // .VSWITCH(VDDIO), 
                                  // .VDDIO_Q(), 
                                  // .VCCHIB(VCCD1), 
                                  // .VDDIO(VDDIO), 
                                  // .VCCD(VCCD1), 
                                  // .VSSIO(VSSIO), 
                                  // .VSSD(VSSD1), 
                                  // .VSSIO_Q()
                                        );




sky130_fd_io__top_power_lvc_wpad REF_CLK_PAD ( .P_PAD(REF_CLK), 
                                   .AMUXBUS_A(), 
                                   .AMUXBUS_B()
                                  // .P_CORE(REF_CLK_pll), 
                                  // .BDY2_B2B(VSSA1), 
                                  // .DRN_LVC1(VDDA1), 
                                  // .DRN_LVC2(), 
                                  // .OGC_LVC(), 
                                  // .SRC_BDY_LVC1(VSSA1), 
                                  // .SRC_BDY_LVC2(), 
                                   
                                   //.VSSA(VSSA1), 
                                  // .VDDA(VDDA1), 
                                  // .VSWITCH(VDDIO), 
                                  // .VDDIO_Q(), 
                                  // .VCCHIB(VCCD1), 
                                  // .VDDIO(VDDIO), 
                                  // .VCCD(VCCD1), 
                                  // .VSSIO(VSSIO), 
                                  // .VSSD(VSSD1), 
                                  // .VSSIO_Q()
                                        );


sky130_fd_io__top_power_lvc_wpad CLK_PAD ( .P_PAD(CLK), 
                                   .AMUXBUS_A(), 
                                   .AMUXBUS_B()
                                  // .P_CORE(CLK_pll), 
                                  // .BDY2_B2B(VSSA1), 
                                  // .DRN_LVC1(VDDA1), 
                                  // .DRN_LVC2(), 
                                  // .OGC_LVC(), 
                                  // .SRC_BDY_LVC1(VSSA1), 
                                  // .SRC_BDY_LVC2(), 
                                   
                                  // .VSSA(VSSA1), 
                                  // .VDDA(VDDA1), 
                                  // .VSWITCH(VDDIO), 
                                  // .VDDIO_Q(), 
                                  // .VCCHIB(VCCD1), 
                                  // .VDDIO(VDDIO), 
                                  // .VCCD(VCCD1), 
                                  // .VSSIO(VSSIO), 
                                  // .VSSD(VSSD1), 
                                  // .VSSIO_Q()
                                        );                                        



sky130_fd_io__top_power_lvc_wpad VDDA_PAD ( .P_PAD(VDDA), 
                                   .AMUXBUS_A(), 
                                   .AMUXBUS_B()
                                  // .P_CORE(VDDA_pll), 
                                  // .BDY2_B2B(VSSA1), 
                                  // .DRN_LVC1(VDDA1), 
                                  // .DRN_LVC2(), 
                                  // .OGC_LVC(), 
                                  // .SRC_BDY_LVC1(VSSA1), 
                                  // .SRC_BDY_LVC2(), 
                                   
                                   //.VSSA(VSSA1), 
                                  // .VDDA(VDDA1), 
                                  // .VSWITCH(VDDIO), 
                                  // .VDDIO_Q(), 
                                  // .VCCHIB(VCCD1), 
                                  // .VDDIO(VDDIO), 
                                  // .VCCD(VCCD1), 
                                  // .VSSIO(VSSIO), 
                                  // .VSSD(VSSD1), 
                                  // .VSSIO_Q()
                                        );      


sky130_fd_io__top_ground_lvc_wpad VSSA_PAD ( .G_PAD(VSSA), 
                                    .AMUXBUS_A(), 
                                    .AMUXBUS_B()
                                   // .G_CORE(VSSA_pll), 
                                   // .BDY2_B2B(VSSA1), 
                                   // .DRN_LVC1(VDDA1), 
                                   // .DRN_LVC2(), 
                                   // .OGC_LVC(), 
                                   // .SRC_BDY_LVC1(VSSA1), 
                                   // .SRC_BDY_LVC2(), 
                                    
                                   // .VSSA(VSSA1), 
                                   // .VDDA(VDDA1), 
                                   // .VSWITCH(VDDIO), 
                                   // .VDDIO_Q(), 
                                   // .VCCHIB(VCCD1), 
                                   // .VDDIO(VDDIO), 
                                   // .VCCD(VCCD1), 
                                   // .VSSIO(VSSIO), 
                                   // .VSSD(VSSD1), 
                                   // .VSSIO_Q()
                                         );



sky130_fd_io__top_ground_lvc_wpad VSSD_PAD ( .G_PAD(VSSD), 
                                    .AMUXBUS_A(), 
                                    .AMUXBUS_B()
                                   // .G_CORE(VSSD_pll), 
                                   // .BDY2_B2B(VSSA1), 
                                   // .DRN_LVC1(VDDA1), 
                                   // .DRN_LVC2(), 
                                   // .OGC_LVC(), 
                                   // .SRC_BDY_LVC1(VSSA1), 
                                   // .SRC_BDY_LVC2(), 
                                    
                                   // .VSSA(VSSA1), 
                                   // .VDDA(VDDA1), 
                                   // .VSWITCH(VDDIO), 
                                   // .VDDIO_Q(), 
                                   // .VCCHIB(VCCD1), 
                                   // .VDDIO(VDDIO), 
                                   // .VCCD(VCCD1), 
                                   // .VSSIO(VSSIO), 
                                   // .VSSD(VSSD1), 
                                   // .VSSIO_Q()
                                         );



sky130_fd_io__top_power_lvc_wpad VDDD_PAD ( .P_PAD(VDDD), 
                                   .AMUXBUS_A(), 
                                   .AMUXBUS_B()
                                  // .P_CORE(VDDD_pll), 
                                  // .BDY2_B2B(VSSA1), 
                                  // .DRN_LVC1(VDDA1), 
                                  // .DRN_LVC2(), 
                                  // .OGC_LVC(), 
                                 //  .SRC_BDY_LVC1(VSSA1), 
                                  // .SRC_BDY_LVC2(), 
                                   
                                  // .VSSA(VSSA1), 
                                  // .VDDA(VDDA1), 
                                 //  .VSWITCH(VDDIO), 
                                  // .VDDIO_Q(), 
                                  // .VCCHIB(VCCD1), 
                                  // .VDDIO(VDDIO), 
                                  // .VCCD(VCCD1), 
                                  // .VSSIO(VSSIO), 
                                  // .VSSD(VSSD1), 
                                  // .VSSIO_Q()
                                        );      






sky130_ef_io__vddio_hvc_pad  VDDR_PAD (.AMUXBUS_A(), 
                                      .AMUXBUS_B(), 
                                      .DRN_HVC(VDDA),
	                              .SRC_BDY_HVC(VSSA1),
	                              .VSSA(VSSA1), 
	                              .VDDA(VDDA1), 
	                              .VSWITCH(VDDIO), 
	                              .VDDIO_Q(), 
	                              .VCCHIB(VCCD1), 
	                              .VDDIO(VDDR), 
	                              .VCCD(VCCD1),
	                              .VSSIO(VSSIO), 
	                              .VSSD(VSSD1), 
	                              .VSSIO_Q()
                                       );



sky130_fd_io__top_ground_hvc_wpad GNDR_PAD ( .G_PAD(GNDR),
                                    .AMUXBUS_A(), 
                                    .AMUXBUS_B()
                                   // .G_CORE(GNDR_pll), 
                                   // .DRN_HVC(VDDA1), 
                                   // .OGC_HVC(), 
                                   // .SRC_BDY_HVC(VSSA1),
                                   // .VSSA(VSSA1), 
                                   // .VDDA(VDDA1), 
                                   // .VSWITCH(VDDIO), 
                                   // .VDDIO_Q(), 
                                  //  .VCCHIB(VCCD1), 
                                   // .VDDIO(VDDIO), 
                                    //.VCCD(VCCD1), 
                                    //.VSSIO(VSSIO), 
                                   // .VSSD(VSSD1), 
                                   // .VSSIO_Q()
                                         );



sky130_ef_io__vdda_hvc_pad  VDDO_PAD (.AMUXBUS_A(), 
                                      .AMUXBUS_B(), 
                                      .DRN_HVC(VDDA),
	                              .SRC_BDY_HVC(VSSA1),
	                              .VSSA(VSSA1), 
	                              .VDDA(VDDO), 
	                              .VSWITCH(VDDIO), 
	                              .VDDIO_Q(), 
	                              .VCCHIB(VCCD1), 
	                              .VDDIO(VDDIO), 
	                              .VCCD(VCCD1),
	                              .VSSIO(VSSIO), 
	                              .VSSD(VSSD1), 
	                              .VSSIO_Q()
                                       );
  



sky130_fd_io__top_ground_hvc_wpad GNDO_PAD ( .G_PAD(GNDO),
                                    .AMUXBUS_A(), 
                                    .AMUXBUS_B()
                                   // .G_CORE(GNDO_pll), 
                                   // .DRN_HVC(VDDA1), 
                                   // .OGC_HVC(), 
                                   // .SRC_BDY_HVC(VSSA1),
                                   // .VSSA(VSSA1), 
                                   // .VDDA(VDDA1), 
                                   // .VSWITCH(VDDIO), 
                                   // .VDDIO_Q(), 
                                   // .VCCHIB(VCCD1), 
                                   // .VDDIO(VDDIO), 
                                   // .VCCD(VCCD1), 
                                   // .VSSIO(VSSIO), 
                                   // .VSSD(VSSD1), 
                                   // .VSSIO_Q()
                                         );
 
 
sky130_ef_io__corner_pad corner_1 (.AMUXBUS_A(), 
                                   .AMUXBUS_B(), 
	                           .VSSA(VSSA1), 
	                           .VDDA(VDDA1), 
	                           .VSWITCH(VDDIO), 
	                           .VDDIO_Q(), 
	                           .VCCHIB(VCCD1), 
	                           .VDDIO(VDDIO), 
	                           .VCCD(VCCD1),
	                           .VSSIO(VSSIO), 
	                           .VSSD(VSSD1), 
	                           .VSSIO_Q()
                                       );
  
  
  
sky130_ef_io__corner_pad corner_2 (.AMUXBUS_A(), 
                                   .AMUXBUS_B(), 
	                           .VSSA(VSSA1), 
	                           .VDDA(VDDA1), 
	                           .VSWITCH(VDDIO), 
	                           .VDDIO_Q(), 
	                           .VCCHIB(VCCD1), 
	                           .VDDIO(VDDIO), 
	                           .VCCD(VCCD1),
	                           .VSSIO(VSSIO), 
	                           .VSSD(VSSD1), 
	                           .VSSIO_Q()
                                       );
 
 
sky130_ef_io__corner_pad corner_3 (.AMUXBUS_A(), 
                                   .AMUXBUS_B(), 
	                           .VSSA(VSSA1), 
	                           .VDDA(VDDA1), 
	                           .VSWITCH(VDDIO), 
	                           .VDDIO_Q(), 
	                           .VCCHIB(VCCD1), 
	                           .VDDIO(VDDIO), 
	                           .VCCD(VCCD1),
	                           .VSSIO(VSSIO), 
	                           .VSSD(VSSD1), 
	                           .VSSIO_Q()
                                       );
 
 
 
sky130_ef_io__corner_pad corner_4 (.AMUXBUS_A(), 
                                   .AMUXBUS_B(), 
	                           .VSSA(VSSA1), 
	                           .VDDA(VDDA1), 
	                           .VSWITCH(VDDIO), 
	                           .VDDIO_Q(), 
	                           .VCCHIB(VCCD1), 
	                           .VDDIO(VDDIO), 
	                           .VCCD(VCCD1),
	                           .VSSIO(VSSIO), 
	                           .VSSD(VSSD1), 
	                           .VSSIO_Q()
                                       );
 
 

 
 
 
                                     
endmodule                                         
                                         




